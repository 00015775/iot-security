PK
     Ps�[N�Y�R�  R�     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_0":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_0":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1":["pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_5"],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_1":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_2":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_2":["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_27"],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_3":["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9"],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_3":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_4":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_4":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_5":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_5":["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1"],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_6":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_6":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_7":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_7":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_8":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_8":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9":["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_3"],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9":["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_4","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_1"],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_10":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_10":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_11":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_11":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_12":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_12":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_13":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_13":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_14":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_14":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_15":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_15":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_16":[],"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_16":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_0":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_1":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_2":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_3":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_4":["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9"],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5":["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9"],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_6":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_7":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_8":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_9":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_10":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_11":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_12":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_13":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_14":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_15":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_16":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_17":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_18":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_19":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_20":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_21":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_22":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_23":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_24":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_25":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_26":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_27":["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_2"],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_28":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_29":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_30":[],"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_31":[],"pin-type-component_0df04e1e-7267-4d16-94d0-338b96ff5fbd_0":[],"pin-type-component_0df04e1e-7267-4d16-94d0-338b96ff5fbd_1":[],"pin-type-component_0b7f63ea-a2de-4b3f-a624-8eac33fdc1f7_0":[],"pin-type-component_0b7f63ea-a2de-4b3f-a624-8eac33fdc1f7_1":[],"pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0":["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1"],"pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_1":["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9"],"pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_0":[],"pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_1":[],"pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_2":[]},"pin_to_color":{"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_0":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_0":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1":"#005F39","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_1":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_2":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_2":"#ff2600","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_3":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_3":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_4":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_4":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_5":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_5":"#005F39","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_6":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_6":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_7":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_7":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_8":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_8":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9":"#b51a00","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_10":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_10":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_11":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_11":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_12":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_12":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_13":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_13":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_14":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_14":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_15":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_15":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_16":"#000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_16":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_0":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_1":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_2":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_3":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_4":"#b51a00","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_6":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_7":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_8":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_9":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_10":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_11":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_12":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_13":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_14":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_15":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_16":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_17":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_18":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_19":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_20":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_21":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_22":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_23":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_24":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_25":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_26":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_27":"#ff2600","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_28":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_29":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_30":"#000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_31":"#000000","pin-type-component_0df04e1e-7267-4d16-94d0-338b96ff5fbd_0":"#000000","pin-type-component_0df04e1e-7267-4d16-94d0-338b96ff5fbd_1":"#000000","pin-type-component_0b7f63ea-a2de-4b3f-a624-8eac33fdc1f7_0":"#000000","pin-type-component_0b7f63ea-a2de-4b3f-a624-8eac33fdc1f7_1":"#000000","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0":"#005F39","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_1":"#b51a00","pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_0":"#000000","pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_1":"#000000","pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_2":"#000000"},"pin_to_state":{"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_0":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_0":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_1":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_2":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_2":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_3":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_3":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_4":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_4":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_5":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_5":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_6":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_6":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_7":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_7":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_8":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_8":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_10":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_10":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_11":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_11":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_12":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_12":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_13":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_13":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_14":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_14":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_15":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_15":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_16":"neutral","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_16":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_0":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_1":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_2":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_3":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_4":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_6":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_7":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_8":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_9":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_10":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_11":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_12":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_13":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_14":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_15":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_16":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_17":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_18":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_19":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_20":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_21":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_22":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_23":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_24":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_25":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_26":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_27":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_28":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_29":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_30":"neutral","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_31":"neutral","pin-type-component_0df04e1e-7267-4d16-94d0-338b96ff5fbd_0":"neutral","pin-type-component_0df04e1e-7267-4d16-94d0-338b96ff5fbd_1":"neutral","pin-type-component_0b7f63ea-a2de-4b3f-a624-8eac33fdc1f7_0":"neutral","pin-type-component_0b7f63ea-a2de-4b3f-a624-8eac33fdc1f7_1":"neutral","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0":"neutral","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_1":"neutral","pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_0":"neutral","pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_1":"neutral","pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_2":"neutral"},"next_color_idx":6,"wires_placed_in_order":[["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_27","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_2"],["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9"],["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9"],["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_3"],["pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1"],["pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1"],["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_4","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9"],["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_1"],["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_5"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_27","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_2"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9"]]],[[["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5"]],[]],[[],[["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9"]]],[[],[["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_3"]]],[[],[["pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1"]]],[[["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0"]],[]],[[],[["pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1"]]],[[],[["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_4","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9"]]],[[],[["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_1"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_5"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_0":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_0":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1":"0000000000000002","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_1":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_2":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_2":"0000000000000000","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_3":"0000000000000001","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_3":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_4":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_4":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_5":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_5":"0000000000000002","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_6":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_6":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_7":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_7":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_8":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_8":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9":"0000000000000001","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9":"0000000000000003","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_10":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_10":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_11":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_11":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_12":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_12":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_13":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_13":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_14":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_14":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_15":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_15":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_16":"_","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_16":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_0":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_1":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_2":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_3":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_4":"0000000000000003","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5":"0000000000000001","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_6":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_7":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_8":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_9":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_10":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_11":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_12":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_13":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_14":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_15":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_16":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_17":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_18":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_19":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_20":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_21":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_22":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_23":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_24":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_25":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_26":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_27":"0000000000000000","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_28":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_29":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_30":"_","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_31":"_","pin-type-component_0df04e1e-7267-4d16-94d0-338b96ff5fbd_0":"_","pin-type-component_0df04e1e-7267-4d16-94d0-338b96ff5fbd_1":"_","pin-type-component_0b7f63ea-a2de-4b3f-a624-8eac33fdc1f7_0":"_","pin-type-component_0b7f63ea-a2de-4b3f-a624-8eac33fdc1f7_1":"_","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0":"0000000000000002","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_1":"0000000000000003","pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_0":"_","pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_1":"_","pin-type-component_2677a2d4-47ab-4974-aa4d-91ba8a64f2f9_2":"_"},"component_id_to_pins":{"d3d841d9-84c0-4783-b9b7-3d9d99c59f90":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"0df04e1e-7267-4d16-94d0-338b96ff5fbd":["0","1"],"0b7f63ea-a2de-4b3f-a624-8eac33fdc1f7":["0","1"],"741beb8c-3e81-420b-83f9-9c980f603734":["0","1"],"f8f07702-f832-4a42-87ea-64a72d994d50":[],"2677a2d4-47ab-4974-aa4d-91ba8a64f2f9":["0","1","2"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_27","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_2"],"0000000000000001":["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_3"],"0000000000000002":["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0","pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_5"],"0000000000000003":["pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9","pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_4","pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_1"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3"},"all_breadboard_info_list":["ce2376b2-6fad-4481-865e-d6c07eea78ee_17_2_False_880_340_up"],"breadboard_info_list":["ce2376b2-6fad-4481-865e-d6c07eea78ee_17_2_False_880_340_up"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[1341.25,462.50000000000045],"typeId":"23db5403-7550-740c-a02b-8b3755757442","componentVersion":1,"instanceId":"d3d841d9-84c0-4783-b9b7-3d9d99c59f90","orientation":"up","circleData":[[1322.5,605],[1337.5,605],[1352.5,605],[1367.5,605],[1382.5,605],[1397.5,605],[1412.5,605],[1427.5,605],[1457.5,605],[1472.5,605],[1487.5,605],[1502.5,605],[1517.5,605],[1532.5,605],[1268.5,320.00000000000034],[1283.5,320.00000000000034],[1298.5,320.00000000000034],[1313.5,320.00000000000034],[1328.5,320.00000000000034],[1343.5,320.00000000000034],[1358.5,320.00000000000034],[1373.5,320.00000000000034],[1388.5,320.00000000000034],[1403.5,320.00000000000034],[1427.5,320.00000000000034],[1442.5,320.00000000000034],[1457.5,320.00000000000034],[1472.5,320.00000000000034],[1487.5,320.00000000000034],[1502.5,320.00000000000034],[1517.5,320.00000000000034],[1532.5,320.00000000000034]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"cabb5eed-764a-4254-9f14-10ad922ef5bd\",\"explorerHtmlId\":\"8eae3b46-36e2-4d26-b3c3-313aef96005d\",\"nameHtmlId\":\"001bd08b-6a2f-4d1c-87ee-b69ac60f8f77\",\"nameInputHtmlId\":\"79e009c9-8ef6-4d7a-9248-bd8c4dec713f\",\"explorerChildHtmlId\":\"9a492043-39bc-441d-b8d0-74f4d5bc1d36\",\"explorerCarrotOpenHtmlId\":\"ed0de702-c154-4e16-b6bb-2ca2223f8cf8\",\"explorerCarrotClosedHtmlId\":\"043fb8f4-cd20-4f93-887a-d93db74574fc\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"ba1888ef-4bfd-469e-938d-64128c39725c\",\"explorerHtmlId\":\"994697c6-87c0-418f-bb4b-ac8cc3885c49\",\"nameHtmlId\":\"fe32aff7-d5ef-48bf-87d0-dc7c2e994f21\",\"nameInputHtmlId\":\"61a2a8af-8996-45b0-9773-dc97c223277c\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"c0e20c32-e700-4943-aebe-7af05ed74423\",\"explorerHtmlId\":\"9fa41b06-0b9d-4272-bcae-cf69dc41b9a0\",\"nameHtmlId\":\"3be67a60-6434-4df5-b573-a388a1db6b41\",\"nameInputHtmlId\":\"e1e53cd0-b227-419a-97b5-3958bc0daece\",\"code\":\"\"},0,","codeLabelPosition":[1341.25,305.0000000000004],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[947.4374995000001,458.2385495],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"0df04e1e-7267-4d16-94d0-338b96ff5fbd","orientation":"left","circleData":[[947.5,485],[947.5,429.2958484999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"1000","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[925,380],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"0b7f63ea-a2de-4b3f-a624-8eac33fdc1f7","orientation":"up","circleData":[[902.5,380],[947.5,380]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[876.7518610000003,124.60839349999992],"typeId":"3ce813a8-322b-4f90-a9f5-e0d3b4eaeefb","componentVersion":1,"instanceId":"741beb8c-3e81-420b-83f9-9c980f603734","orientation":"left","circleData":[[947.5,215],[936.6004419999999,215.06061799999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Simple Fan (2-wire with NPN Transistor): \n  Required Components:\n   - 1x NPN Transistor (2N2222, BC547, or similar)\n   - 1x 1kΩ Resistor\n   - 1x Diode 1N4007 (for protection)\n\nArduino Pin 4 → 1kΩ Resistor → Transistor Base (middle pin)\nTransistor Emitter (left/right pin) → Arduino GND\nTransistor Collector (left/right pin) → Fan GND (-)\nFan VCC (+) → Arduino 5V\nDiode (1N4007): Cathode to Arduino 5V, Anode to Fan GND","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1251.5520649625084,139.29935981486483],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"f8f07702-f832-4a42-87ea-64a72d994d50","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[804.1677175,380.30182700000023],"typeId":"10d13646-c889-4b39-93c7-eebbfe2262dd","componentVersion":1,"instanceId":"2677a2d4-47ab-4974-aa4d-91ba8a64f2f9","orientation":"left","circleData":[[842.5,395],[842.5,380],[842.5,365]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"21.58897","left":"758.94182","width":"813.55818","height":"608.41103","x":"758.94182","y":"21.58897"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_2\",\"endPinId\":\"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_27\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_2_4\",\"rawEndPinId\":\"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_27\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1007.5000000000_380.0000000000\\\",\\\"1022.5000000000_380.0000000000\\\",\\\"1022.5000000000_290.0000000000\\\",\\\"1472.5000000000_290.0000000000\\\",\\\"1472.5000000000_320.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9\",\"endPinId\":\"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9_0\",\"rawEndPinId\":\"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_485.0000000000\\\",\\\"835.0000000000_485.0000000000\\\",\\\"835.0000000000_650.0000000000\\\",\\\"1397.5000000000_650.0000000000\\\",\\\"1397.5000000000_605.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_3\",\"endPinId\":\"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_3_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_9_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.5000000000_395.0000000000\\\",\\\"902.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1\",\"endPinId\":\"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_5\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_5_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.5000000000_365.0000000000\\\",\\\"910.0000000000_365.0000000000\\\",\\\"910.0000000000_320.0000000000\\\",\\\"970.0000000000_320.0000000000\\\",\\\"970.0000000000_417.5000000000\\\",\\\"947.5000000000_417.5000000000\\\",\\\"947.5000000000_425.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1\",\"endPinId\":\"pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ce2376b2-6fad-4481-865e-d6c07eea78ee_0_1_2\",\"rawEndPinId\":\"pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"872.5000000000_365.0000000000\\\",\\\"880.0000000000_365.0000000000\\\",\\\"880.0000000000_297.5000000000\\\",\\\"947.5000000000_297.5000000000\\\",\\\"947.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#b51a00\",\"startPinId\":\"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9\",\"endPinId\":\"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_4\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9_4\",\"rawEndPinId\":\"pin-type-component_d3d841d9-84c0-4783-b9b7-3d9d99c59f90_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1007.5000000000_485.0000000000\\\",\\\"1007.5000000000_477.5000000000\\\",\\\"1037.5000000000_477.5000000000\\\",\\\"1037.5000000000_635.0000000000\\\",\\\"1382.5000000000_635.0000000000\\\",\\\"1382.5000000000_605.0000000000\\\"]}\"}","{\"color\":\"#b51a00\",\"startPinId\":\"pin-type-breadboard_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9\",\"endPinId\":\"pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ce2376b2-6fad-4481-865e-d6c07eea78ee_1_9_2\",\"rawEndPinId\":\"pin-type-component_741beb8c-3e81-420b-83f9-9c980f603734_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"977.5000000000_485.0000000000\\\",\\\"970.0000000000_485.0000000000\\\",\\\"970.0000000000_672.5000000000\\\",\\\"782.5000000000_672.5000000000\\\",\\\"782.5000000000_252.5000000000\\\",\\\"936.6004420000_252.5000000000\\\",\\\"936.6004420000_215.0606180000\\\"]}\"}"],"projectDescription":""}PK
     Ps�[               jsons/PK
     Ps�[�赚#  �#     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino UNO","category":["Microcontroller"],"userDefined":false,"id":"23db5403-7550-740c-a02b-8b3755757442","subtypeDescription":"","subtypePic":"0b351edc-7875-4477-b820-546ce15be531.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Fan","category":["User Defined"],"userDefined":true,"id":"3ce813a8-322b-4f90-a9f5-e0d3b4eaeefb","subtypeDescription":"","subtypePic":"9ce856c6-be81-4769-87b3-53be9928d02a.png","iconPic":"627fe4d2-0152-4b97-938d-4b9176d7a483.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"12.40259","numDisplayRows":"10.33548","pins":[{"uniquePinIdString":"0","positionMil":"17.51879,45.11974","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"17.11467,117.78346","isAnchorPin":false,"label":"5V"}],"pinType":"wired"},"properties":[],"componentVersion":1,"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":" A3144 Magnetic Hall Effect Sensor","category":["User Defined"],"id":"10d13646-c889-4b39-93c7-eebbfe2262dd","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6a97e33c-aa93-4e7b-a2bd-349ce97096b8.png","iconPic":"e65d6d59-bd1f-4659-a32c-fe6c1b0070ef.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"2.74401","numDisplayRows":"6.03012","pins":[{"uniquePinIdString":"0","positionMil":"39.21268,45.95745","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"139.21268,45.95745","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"239.21268,45.95745","isAnchorPin":false,"label":"OUT"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     Ps�[               images/PK
     Ps�[P��/ǽ  ǽ  /   images/0b351edc-7875-4477-b820-546ce15be531.png�PNG

   IHDR  u  v   ��:   sBIT|d�    IDATx���}tSwz/��$۲0���Mblc0fB��3���@��0�b�!d�qN�bν'�tAgڣ�rf��i��Ճ���M�8�Ms�z��� N�`L�~��-�/��ClE�e[/{k���Y+kY��O��g?���S��ҡ�D�P�C���{HDDDDD�;����_��{�R�=�p����V)v9""""��Ή�:�t(I�R�)xZ�Q��5�cR�GBנP�@��x�1�cR��+o6I���t�|�&�I ����W��ǙM~��<>/(�^h�J""""
O����=�p���`T��F��:ix./M�8�IV�0<<,�0������ ~�}�M�Kb�J�/^:���Q��)��ӣ ]��+���!�L-[�,(q��~cP�Qx��+u>HT�*�GT�K�N�F#�0�����BN�T���@{��c�NQ9*���!�S�=�p�n�DDDDD��abg�{�aR祄W��="""""�G('v�~I�v|b��
[�M�6ן)�B�;JX�&"""�^�N�dRDO�f੅�`�b���y��A�����DF=T*~��"�bb�������_��g}� �L|v;>��f�@�|y`��6��~�PN�JU�Pث�B�GIDDD^B1��^Jx�PI�g9������~�1��y��\oo/���@�Z����80w��Y���G'Q�f
���c��	��0����'�C
���䎈��h�P�:�aLv��0�Ə��8��/�ҡ:m�Ҡ ^��٨���w��cqyX˸�˸�Ըb����q7��
B�b�J��X���Z���qu\e����MRʕP��{`<�}���R�a��A�<�,]�q��G��s"�������m>=?*v�~I��v\���H�����_�W�J�@�g�DDDDA
]1���1!����(F~�r;"""���N���);`W�*���	F~�r���`�#"""

�r�f��0e�tk�f����봯��f �S&&�ݮC�RA�R1.�2.�W,6����O�P ֋�y�q7��I��f��b�`xx `�Za��  � ��������"��<x��:�����e�?�S `||f�FGGKllRSS��!�2.�2��q�b��1:j���H��R*��?���\�e\�<n8`RG����`�Zq���ޅ��?�6�������9Z-���/��#�uB�)�o�<`�P�B�|ǟ_W*�P��D h��q�?>�v�Wg�˸�˸���B��J�9s�tA*\����xu1ʸ�˸��L���������z��c;Vcn������ݻ���|���>�����ݻHNLD�R	����	L���X`������͎/&&�y��]�����BZf&������(�k�Z���?}(��"<����8f}��6��1���F�oV�[���pa�P(`���q�q%�+�@.H]/D�q7�qCYd���fý{���ڊ�`�Ղ�y�H���%&c�}p���� ��#QJE,���0������F���`Q����b����ܩ����)lF��� 7&����q�q7Xq������˸��	���&A[k+�:��א9/��x���`��8J qJ%�J$ƨ`�����������'�=�RRR�z���.�Z��ƕ6c�MPR8.�ZZZ�~�ʕ�D�0c\�e\ƕ�J����;ר�fɒ<Q.D�q72ӟ�|U��Ʉ/._��cu��j��Q����qc
̍�A�J��]��f5z�菡/-EFF�#�"v4�=W#�x�I�ꛦ@�`
�����&�)�e\�e\�X,V�_���~�q7��"��d��_��G���I0wv`��W�1
t11xT���}�O���B{{��1"�ݎ�oa0�K4������:��d�o��a�ڄ�9��&��$�� �T���x�_���＃��nIbE"��� �&�D����(�0��r###�M}=p���`W�A(M�*H���D�u4��?��ݻ��$""""�DLꢘ�f���1|�7��SWWP�����k���gQ6��t��W��!Q4aR��Z[��#;I�� 't�X�ɱ1�{���ٳA������(0��R###�ZW�m"�;�2�r:j��qq���Z���m� !�r�a2�MY"��������(����B�sc����e��F��vxW~�kV눈���|��.
Y,�7��|�C==r�c�����~�vÜV(V��ЫE&uQ���Z�#���N��,N�D�݆�S��J�
�J���@DDD�b�@4��ݥؖ�,�Y��5O�C��`���54`�ܹ�Z���
�����s����{H�'��9?>T��A'Ʊ��ӽ~nll�!�q�qe������u			�˸�BqC�� �L����z����_H�X,�tu ���m0�X��!t~�%��^QJn
@7��C�^�N� @�MY!�q��Ұx�b�~gxxV��7H�q�qŌ+�����;V���Ì˸�+s�P��Q���/��T���/�P<�Q*�Q����,�PB��.N"%��@������D�/!!j��q�q7hqŒ��������{j�:�J�2.�7T1��2��혫���phn���cm]��~'�PB�B�����=��WU(��K/��^�1.�2.����Q����˸�x�P��Qftp�PȾ��LT
��^ht�Uj��h����^:��P(���u�J����.�			���^Mkf\�e\��5�X
E��!)�f*)�2.�70��2C�3�'�J���.���(xZεu��!�*]LLFGG���+�x�v;�2.�2�$qŢT*#���q�\1��211*����ƬT
�G��P���P��/^n
fܹ�*W /r�͆��Q��ĸ�˸���v�,�g\�e���5uDaJ�b&�F�t()X1���P�Jc�����E�ؘ�(�*Y��B��J���nΏ�ؔ�6G!""""q1�#
sBb7�Ǉ$��oʙ����(ېh��j4rcF���,��B�@A�Mِ��������])�x�P�æ(~�����w2�����:�<�������a1.�2.�J�A�<|�rیω���q7��"^9{)��C%1P�	��K��?��Ǽn����+z�իG��~��|y��	Q�-���	Ld/Ď��I����%9n����Ʉ�f~��@���ʡ
�BiP EQD3���,�+uQF����/>Gl|<F����G�v;�͐{aK���1P�Ѿ��'v،C�Û/x���ĩT�
����Qx`Re2�z|u�#h�ڐL���vL���Z�B=�O+�|Z�w쯼��ݎ(lm6�\����

{�(Q(P L�%"""����.�:�ڝ^<��>�R?O��&��		S�#Y����;�?P�v;,6;�=���P�i�Oʩݑ�8N��Z�>��  �ͷq����#"""�hƤ.����M��ۛ^=�؎՘+�ǳ`u�?�-�B�Z7f�#5�		r�h���4��� �Ä �m\���.�2��,��`�Z�����Iu46m�5�������CDD���A�{�i�3����*�P܌���۠��?�{(DS�4jԾ��-��.@��2��I5�v�PV���t�ㅙ�0���/+�'""���J]R'$ ��߃��fHU�6�s�h�j��B4E�~1����� ��q ���#;E���AY�竺=ې�Q��ݏQw���gBbW�gJ�����$�()�%i�����ꛤQ���#�����U4��`	�����I]�Z�y3>�������H�6F�6<U�W�y����6��Q�� P�w�3�[�� �a�ԕ�03�oECKǔ�7u����h����X��3Wd%��$�U��P���V�0[��kB��IΧ$�Ez$͉��B3�zM0�;Ө��ك�O���G�؁�Y}�rпk9�:6?�f4�t�� �9% Z:`�o�}��1���P����(�#'U��7�a8�i�n(5T� �T������R�π�]����Iա��է/OIn�vJ���Caf:*��(�L��A��I]�R'$������e$��b�����2a��j�!q�rV�$�؍ӈ��t�Q�|��4�q��}�^??ntK��J[`�1��[U;a�o��TI�03M�=��.�"�@W�F� �]��8V,q\��t�$/��b�����9�Iա�j�󮼐 U�_���-h�Daf:��lsܬ��.I�FyAJ�fKrq�� ��B3J�`ܽ	m�&�w�|��+�B�!$��bT�_����]��$�%yYh�ډE;O�d���1�p�ؚ<��_��B�]Q���B���)�����s~�m�&g���HҨQ��.˿CR�(ңzG)�zMh���o���AR%�rbR����p��e��Q��`�b�� ,6�J��/�"�����'��^�Ռ��x�I|��Ը��� ��+nt�>���:���˜�i��P�w����[��:��iҜx���L�<�ԫ��:	��s�*]����b�P߈���h�쁡����0�����fA����8Ū�+U�IS���ls\ؾ��(q�V���0l~ʭr"er'�o%�G0`�¸{�:{�>��ӗ/m~J��M8\+w�k~�><-J�$�U�W�����g����U��r$�6!�5�7:���F��)��5l~����`��*�^�S��*�����2�Z���|�#�%��(�����?�	]����ڂ�ؙ'&`��P��͎�+����^%vb��&�3�s����Gб�ȹ��5����h=�t�^��4���gO�	�J��=DI^�ǋ�����VSg���\����k�����f���:{P��%JL)�XP��Ǩh�pT�&�-h��ASg���sRu��v�y��1����vK��-I�vN��:��B3�o�qU�v�#BE�����b)��r;?��\q|��r{�����Ϸ���oEݞm0��$i����9��k
ڍ:�����^�O��o-��(�NH��?z	��7�@F��:����Yl6Xl6<��z}PbF#�+�l��TqgJ�H��wocw�_���6�fck*��=f��4���#p�J'֜T�E}��V���rR�n���z��
����sKĎ+�f/4;�r����V �zMn�[CKrR�S�����dm[E��9�q��b^��A��M0���V-��b��n������3��{1�}0[Q��ǎX{�IV}5�7b`Ă��U(������0[��TeMҨk7E�Ć&u�y�����������I_��yX���{�R��g���J��%vR����I��	�_b�K?F~َ��|���:bO���iHr�<����6���]mA��RwoBCK�V��X��<����C��R��e�����ݛд�nu�;J��ԕ�WjBr��Q�di�#����B3��ls�w���>V�_�;'ޙX�y�?0b�m�p�w0[a�Ќ�T�֯���j�5���0��PV�ܣS*7�a(+F�ي�3W��h)/�s~O�|�B\C� n�;oX	�_��I����Q	��N&�$�I�:*ۓ�/���(_����Hä� 8���j���~�0��+I�q��	&�
<��V�$$ub%���+�kb���5���Q/A�`�xu�t�l5ቶiH�;J���O�i��tęr���	�/��W����3WP^���-�><-�U��T �)�U�v$)��-q0�7��܀�*��.W-�u|�;���*li"�6�7����/4;�f��%VBYx��VT}x�ys	�d7w��\AҜx�t�����K�r�|��g�8���,�ñ�I���ZQ��<�B(܌��j'>����r \$�z�$�3��wl�j̍~�mƥ�%l-7��h���=Q�����0n�#&�Q���	�����{�3u%�=v�44#��[̔�(�FG���#K��ێ�1K��v/X���&i�h{mϔ��+�d��<%u{�9�	�֯Dݵ[nI�q�&$͉w�o�".�m���ׄ�w?F���:���H�`�-�3���>(���C��{��J�4'^�q�$'U7�1�	[P��3j��A����_�
	^�>/�r/l{!��TF,S���3.0��Y�~%��e=�� |�#4u��|6���,�+u�F���5�{��܌k�|Z�s���N�d�f�æV���ǲ?�C�Nn�>���1Y�&<�J��S\MW�4�����d`�"ZBmӐ�F0u{�9���0��n�6g�W9)Z�,�FI^�dӢB�1n����dO8Z:B�
�{������ӽ.�_�lǏ��P����*ؘԑGz=2~�:���q���	�qq�%%�n�atx��a�'<_H��혰�a�c:[|<����d�ȅ�{�T�gm�-���<�8����g�8�)��t��>ga�]�$_DDN����/����S��e�����`�b��4�S������9|s�"�{�C��F������v�Y,Ǹ��ݎ���1O��%6bޢEr�I�R����bb�������_��g}�߿/P+��C51Ԙ�΃�l���-�Y���ʊ�����$R�]7[�Nh�`Jw8��G�4$O�w0M6\�1���(Zp�exj�#���{cc�]|����LR������ہ�۝�u7O�뜺hQH�7�]˳�����s������ΰL�����q�g��{}&��[�M�x	ӳ�O��ݙ�����~��;�q=6�u]�S^���M������R�]7ݴ�$�ڹg��Y�S��q�X��|%U����g��d��w#�N�F~Fηv-f��'��z)��ԑ�ع2��$�Ŝ9j|��9ѹ�g��3l6qo8���0G��Wmw<�������fO��!n�(/ȃa�S���"6��tp�:�.@s�}��|+�!/?#�+� ���j/ݐ<f��'��z)���E����P�Th���x��=��B9?]U����F��U��u�~q��2�&���q��Ձ��w]!6/_��Wc߱��� q]ﾇ���b�'p���o�-y�q��E<��2<�jYT�'�ߋ�[ס��)��kr3 &�U�}]�3�P�w;��q3>��ɋ8x�d㐋R����j��s�O����R�".���_$�E%yYh���l�!eB8����$��q���|k'v�s��B�B��lE͹&�w� ���ηv:�h8O\���Z�G�6����gp���{�9g�'o:aL���:"�($T�=ڂ��J���|�ś�w�I|k���E�yM�7?#mJU�sּQ+I���ϭZ6��-���Lꈈ�����FU�WN��^�y�h�ϸ�$u{� ���,Gv�Źp�s�^
��q-�I4}/jvn��XVr�dSm���2}�պH��ʤ��H&����=�$�;0b	�F�MXrRuAm�ϸ���������}?**�b�êJ���-�[�,jΓh�^�۸��y���Bo�-z����A��8�uݴ�9��m�7��7T0�#�r�� !�}Ͼ�ix0<����q A��i2{�Ed\Wf�Ǥj��DW��+�����\�578��uT#��L���;�F��V-CG�P�.z��<����i��dRMì9ׄ-�\�.��A�h�V� &uDQ����T*��
T*�����װXş��so��I��TJ�`�"\��+H1�]����T	N �����T�����ͷe	y���,xU�h;O���z�v9���0+?8���2��ȩ��F�I]��Y>���Gg��y�wa�\uF]������סP��P�����4�Q��~�l�	���i��$g>z�� ��>���mbv�j�������Nː+n�JҨQ��9�:�TA�F��Mn�ih�@��Ge!�3��q��ͬ���nv�:�:(��z�D��n��d��|\����4�H�v)`RDm�Ch���;��G֜�ٟH>��l�|g@�a����<����<���;���6H Q    IDAT,$͉��}2I����-�v�LҨQ�g�c��ӗ�~f�oD[� rR�Ά*rOդ�s�l6/_��Ϡ��e5�=$����{hl������k{���W�'�v�8y���?�_ock��鏮-��w���Ps�	�cZ��#�:""��`ܽɹI���R��}Թ��� ��O!'U'�vEz����	����J�f�di6�:����N���e�;�1��j>B�>����?(y�h;O�����|4�~t���h����D��:""S��0[QQ�w$y~����(ң��G��K�f��f��0n���t���)z��F�EU$�on�4�h;O���F���PŤ��H���>}�Y6��۳%yY�>sE�΅I���n�lE��+n���"I�F�F͆)�N�bתe0����|#���������o��cDD<L�\\\�^4	�%8���&$Jm.SO�d�03]�ꜧ1L69��9&t��N�:[|?���X�F�,����jl""
&u!*F��J5}�>�(�ʐH�
EP^/Q��>}Y��j*���>�$/K�M�#���N$��ߢ��-ؼ|1��fmz����i��1Q�aR���P��������oJg6��9o|�	��A$�6��@ݵ[�*]��������T�_��<T�����&׺�a��ŲĖ�)ɇI]����\�+}��K]}���F��0�o�Z�aE��^�O_���%yY0^hv&�9)ZG�ˇ���y3�=���  K��L��A�(�tDD�I]���i�_���AsHT���j�JT�_9�c��FѧdV�����AT�a(+v�Y[�	��Fne �5���JN��An� ��\���D�]�����:"� 0[=�U�����-��ڂ�T�s���^��Id��f%��?�ڿ���IQDbRGD$���#^=/'U��i;ö����k�4F��i�(�]�����O��HCVr"���s]E�.���řIQ*/�C��%�f%\���3�  �]�"�u/l�MD��03Ezf�;g�q�zM����K��E��<wo���-0�7�M�2�ބ��[R}��w�֯DE�9��o�s�ٱF��n���S��L&��i{m��}�\5u�x]� 
G����d.'U��^���p�]�Q��w�àe{�9���^���Y{�#��uO@�Q56E'9���"=�w�:f��N9~I^e�(/ȋ��I&u��̕)�f�ø{��lC�ύS�����^�=�۳9)ZN|���P��U;QR}d�4.o�9��۟�^ۃ�^SD~�&�Z���qpL�du.���V�;�	n}�6���֮�%u}����)YbQ��+��(�;�a�a+���,��ن��+#�bǤ.J4u����T�(u|��8�K�P����O�]l
���v::�M��}�$/�Q�+�C�F�'͉w��Ä.��^���K7�.6E9��$�������M�=H�p�Pä.��8Od��<M�l��Aҟ����#�"I5��ls�l9}u�n9+ܳMY&""
Ur%Wf+�Vf��xS4I�v4 ���L�HN� ���p��Q�++FN�M�=0^hs�DQ������>IDDaN���x�U�W"'E����M�f^����K�ύ4L�DyA*����������﹖��VT��1eŨ(� �w����-�>}��<��M��.f딵tD�"��FE��y��Q
CY1�Qؓ+�2�7b`����Փ��-0��4"�8`R��֯D���S��D��QJSg��>�$�U����Q;�U�Q���)���g��0^hFaf:J�]e�VʊQw���QX�3��>s�g� 'U��usĂ�Ξo�"i���1��@��/sRu0�ބ$�zʖ�0[�1�><�ܾ�zG);V�������H�Ҡ�H���+��ك�w?���DD6�M����t�������$��?���+80��p���?,Gݞm+iު۳����LV���l��w?"ѳ�O��ݙυ{��ۯ�7w7Hꮶ��j��
^^����t&uDDv�K�b]3&i�0��03U��x̊"��Y$΂aR烵smXk��ܤ���VǨ#�N[�ɱ��mU�n�;۰{��!̝fBRRt��Q᫶;~�����f�˸20[�w:���7��]1f�U��B�_V�m�%$|Ez4�t����y��I��~�j��Z�q�Q�R���������!��KN��U�(EN����MҨ���P��Q��N����*F���>���	���䬘U���hܷ��ݛ`��r$q�W:�Y�E"&u^���~�slԺD�q����Ά&��#���%�F���Z���	8���T��圮�%��2s�����7w{�S(����|#w�L��4�;�W�zM(�(Z:D�j��yA�T�(��Qw�I���''P�~<ܲ�[�N	d��: """
?rW�\��������C��l&uDDDDDDޒ�b�:�L�V�(u&���� �oq���*fR��Q���h��A�ύ0^hƀي�w?v.Aj�ډ�"�dc�+uDQ���Hиw|�^���C�0.�$�3a C}�ǥ?���)��;J1`�F�>u��E��{C�J9���:(X�	s������&G�l�lE��Gg�� L��ԭ�X�#�R�{�`��ݮ��9K-D�o;��H���df+�O_�r�iܽ	%K��4+/�CE�%yY��ꮶ����.Ԯ�_�~�[�jO\�XW�(����(�c��U;a�oDCK�v:��=����F4u��j�JT���������nݼ���
�I����ԡ;'U���?���᪢H��<Y����b&��+��BҜx��MҨ��Q�/�0�#�R�rL�;U���h���PyA��BN�n�}d�d�P��h��m��9m#����^���i��䡩�Ǒ$�T�0�����6>O���7��{
�M�=HҨQ򰃢�di6�V��e�%u���h�5����L��MN��W,���q�¾�Ez��&��\���i�#T�f��૜T��>��(���sw��E��K��/����dUw�����H�r%(�LwV�\-�B���U���0-�P��hn�R��P��&A4��9�:�䡡�f���"�����)�7&'����4կ� o��#�g����-��܎���&7s�sv=��1�����%i��
�l���&W�;J���s��p͞��>���
�4�H�ހ�:""""��]mA�槜2O*��h�왶�2y/Z	chh�pTU&W�Z��2�q�a���,�v&�B�Vw�e��?�ꐓ�CÉOݎ��ҁ�<f�;�ϭ>s�y��wor����Kv��{�C (�<�j[�p�\�[ ϯz��O��b��Z'���t�i�m�&��ن�=�7$�OnL�"Шz4#�݇e"&V���sS��>�jb,�q������3c��$/u�nI:�
&L��vE�Y��Φ�H��؅����4n��U�
3��p��m�eCKJ�]�Uw��m
f��%�W�������2%U�|1��q8x�"���]O.��Gq��.��e�}��g�CG�Z��x>Ea�\[ߠ�1�.�L���+&uD��e�x��$���ĳ�p;� ��w^�,���EX���Ci�j\""�ʹ�+�C�^O����zf�_�ufBu��f;�֯DyA^@S���{la_�~%�֯t{��j�]�Ȧ�geM�
UɆ�gϵ7YCK��rVq��®���Qs�	 P{�j/����L�]W���;�]���'��|�Y�Z�b�W	��B�䛁W���	���(b}���˪N���A��;/��  ���������5.���K|��t�,y��r6Ez���9s�ʖ7rRuHҨ=&��L��Օ�e�-E����}����n��L7ƺ�-0l~
���0[��2��j��
�d�[;q�uj���}'�㍀`��}m��<�s��E2&uDL�krB����`$vL�HJ9)Zgh�!L1�JI^rRu�H�Mi,�4'~��,ꮶ�03I��4N�6�9���칾�%���.���S �����E8���:��ΔXI��1�#")��9�|�0M�x�ٱmA�S!gC[�	�~����f��$5m������kKա���?{��s����j�w�pt��$����*iN���n�ȑ�y����1a��H�����r !!a,!!!V��^zD?2fW���#���?|D�1�;����7��N�fK褊�Mb%EbǄ���TQ�G���0^h������C}#��7�:3�9m1'U��Ι��~_LO׈E��:��K@M;����w���vT��������E�>e�	d���������P(Rl6[�7�x�b���h4���[
 q
;  �_(�a�4h4J ��Ð���x��i�YG:Ψz�\V����N���n闟�������ݛ���g�J��B�W	S��+h�t44��9���2eSs_�����U.��l��p�d��:]zJRZ:`(+�j�_ݵ[���t
3�e�|���G�
�X[z�+�O���6��^�����INN����Wm�
7�Lꈈ�䒤Q��/+P��Ѩ���E��N�JK�3���,��r%"""��!l�0ymI��������������I:Ez��):peE��{
�f&tQ��:"""""�0�JQ��N�";Y+�0�����z�=�"l�s&uDDQ,?#�{�C'�P�������>�j>���.f��#J�|�0Fu:�l�)���f��A�j_������>cn]��#���hX�#�pm��A[�i����T�sASg�c�Ym�+��(/�s�Z����f��n���z0`����e��'i�0��mJ[w��������&��z�8+uDDU���c߱�rCTLꈢ��x5�t���/��S���0��03�~�|�𸡾�ou>nܽ	�ݛP�QO�e�o��
��Iա��� ��=� 8:�5u� 'U��M��a9J��` ��F�������Z��#"���5uD�rRu��Q���� ��\AҜxT�_��k�����U0^h���U��1�2�Q�~�W퓫�\AyA��P��i��03U�FSg ���C}#��l��A��7���A��ADDD~bRGe�֯D�F��ӗ=�|��I5�4j�z^�Zx��>�o�5�03��騻ڂ$����:�4'ާcE#&uDQ�$/f+Z:<�|�l������-(��Bݞmh��P�,'U���Y��03 �������LꈢLҜx�X|���<����F)��b���&)3%h���z�I��xEz������IDDD��Ѭ�VG�w?vLߜ��Y�~�Ǧ(��bʊ����T�3�ބ�Tݔ�~DDDD��:�(30b	h�����Q^��槜�T\;UΖ�yb(+FyA�����?"""�h'߮�D$��k���Q��77YyA�s����+1�7?r�ss;��/4;��4;�qwoB����x�c�}��hfLꈢL���0[QU����'o.4T)/���|��I��v��S�����?@��l�TaBGDDD�#N�$�2f+�><���{�6��SeŨZ�-Ω�M�=�>sŹ����9Ͳj�JT���EN�ι�x��G9咢Nv���Zd�$�m �67�c�\�e2[q��>���k_A�F���4�g̃N����A|��=9��u��:�(Tw�%�&GW���xSg��'��h�5�� m��q>����H��RYQ�G�F�8��8\�Y���~�(�g��L�ks3�� ����_��`ڟ5�v�\k'�o�z�=��*�F�|���f"+9q��)���i�2��8w��[�"�=��������BZF���'��t�,š�Өa��#��_]����4Ծ�Yɉhl�¾cgq��ޔ�w��d�bד˰c������w���[��6>o�k¾cg �6���uO  j/}�|�u���~��'/N;v�F��[��U���?�'/8��؂����®w��z�=d�hQ��)�O�Z�)X��~#b�J��V�|���������O�?��R�@���_��ɏ��DRQ��Ԕ(��3r !!�k�N�P���~�t7�r�(�}�5j�,r{lB��X�bUP)��o�u|jK+���bhb|O[>~���H��u�(��Κ��k�2���V�w�ηvJCj��\�-�\l^�X��w������5Ed�L���[׹%X�V-Á��ܞ����q����P�q�����p�'/�%э�](�����E�s���7p��E\��
�c<y��oLy|�����}�+�q{|��  ��������_!?c�Ǳ��c���n�����7��s��9��"��o���-n�TG���δ�����
���a��_���]n1�q�o~�L<;�����Y�7G��e���/)f��X�#""�'����p{,sI.�sf��x-!6�w����o&�P�%�ZŐ�6>ϭZ6�z�t5*�b�'$KxYɉxqm!^\[����8|x���ӨQ�s��=��������Q:n�L>W�s`Mn��&;y�X�1m�|k��Ǘdz��c ���X� ��؅�ɳ�G�5��Sn���k���@JB<�-��X,w^*�O��ޫ(Ê�#��>&uDD��AF|U� ������^��B��~��I�t��q��8��i���9�$�8f�d�}�<~v�o,
�ؕ0��d�����p������xs딤�d��d�N���*�k�s���8�ډA˨������?5q9���qJ�[���}�㞎8�E��V�c��}oʴda<��p�鷍�]n�����Z&�6�}J��쭎)cl�?�-��)�g'k����޹�N�tR")��lْ�P(*�@\\�)>>>I����}� �-�r�HU�W�_��?�el���}�G�M�&���%A�Pa|�
�Ō����A��>� �`��c�{�F�W���f�~�v<S����Á:F�?xl!��q�����_�!p$��/�������O��{�!��dMn&�� u�
:���B�~��wܞ�x���"I�ƪ��`�2��?:�������7���Y�����͆�w7���|k6<��F���.�?E��.}������څ�N�gh���X�$�[����;�L����:ׄ�'/:�ҝ�:}׻ﻍ���˨�|�ۿ�8�K���;�S����|�|kηv��>��-:�����_��?���������9�������}/t=C#h�@Y�b(
��@�q���.����Y�P(�34�m_�F�5�*�����q��&H)Z���t�����?����#.��Q��:�dU�W�PV��fﮞH�\gw{,1)���n�����I�Z@��a^�b�'L��;_��2�r�G��	SߤZ&���F�S�5w��HC���g̓%�7��%����۸zʚ2!i���63!�6g����MY;(�ף��5uDDRF'�KY�R��Xb����p��-$ν���ˠP�_��K~F��n�m��/6/_��?y�GN����D$�.��Wv��MGX��ӨQ{�\��ų���n��4�pg2[�$k�SovonŮ'���U� ޻�?+7'""�R�e#!1s��	 �զaђ����t\�R1���8�Ņ~b#�]O.ùW���N����{e�ٹa�'� ;E���
��N �G'u^�Cv���݀��Dh�����B���x�e��[皘 ������>���.��5���m�s���L�$
+uDD䗌��ߊo:�����FO����ڧ���V-s�W�dS����n�͋k����uʪ��[��(��ȹ���}�κ}>�nj��]�ۏPhb�����6���`6[1<t�c#r'(�=��3���O^�8],P�k�^EY�&t�����r��v�R��HCv��c2y<D����<u����'��X�#"��d-�.���u�:t����=$�H��]���e�}��kr8��J񼷗?��q�߻e�?�uk��!�{d2[q�ս5���,L�B�-�    IDAT�Q#?c�3�DM���P_�]Ҫ�������{���P޿|��9�2��^���������?CaSw6�!10�#""�`||f`�L`��M����3f(�\[(j�r���o��ý������5��آ_�2�d�J��N�.�׻��K7P����_�b�G��y�ٹ��9�f�k�2�=՞[�Ǜo#��oI��Wy�*�����\���Jvq�ܺ��s"0�#""�%$$  t:Gu�61�ί?C�|xL�l���mA����8 B���A�^���.}�S�⪣�_���/߀6>{�=�]��T�4��iԨ��.�vR�G��|{������qp�:Iײy�0�g��N�$���4����I�F������jo¼�Q�5)��a���m `��)F�)ڀ�E����ɋ�iWb����ɋ8x�"^\[��W�=�0�Į�bK�	����[��ֹ&<�j�o\�wr���B�k�,�:�b���'l*��1k'u�l���}�7<������{���%v\cG�bRGDDS(Uq��O��wU1j<�Y�{�����;�Q١��nj������lE͹&<yQ�QM�hm����k�:�?�]��nS}e2[q��E�6�Ry��c*��uO���B��X��=�6(�i�صj��sq�������w�\��qn]���f߱����t�cp$%�T,'�^{��hS�3�ܶ��vL3Y�����
g�B\�o��A�(j/}���8���#�pp�:d%'���7�wg?þ���{�*|��%""�hS�C��sal\<2�W  ���a}��v&�h�e��B��������~O!�Ǡe������V�<�����6>5;7x�$Ц(�ͭ�<r
��Q���+��y���[|�lj��pp�:���ܺ���.���oL����in窘�b���~}&�^1�x�mQ*�:�:��	�����	{���O^D͹&����7�:߇5��h|e��gϯzܯs���4 "� ��b�͏<�W����q�����ohԌ���qv��C��6%���KG�Qc�������K7������йjl�7j���Ϙ�ڊ-3>'��1B��yc}P:W��]���;~U�6/��)�a$l�1�����E�L*���+�� �۸�����"d�:��zq�I����J��0��Q���z��;��>�l������ߙ�L��G��;�T�o\�״�}��e*�l-��R�+~vv=�{� t��4�mד��n��7�]��hvٚ@.��Q���{}�?�u�(��k��Jr�E��W����bo��Ϙ�׺T]|�$�������3WP}�J���f��ɉ��I]��N��E?֥U9%z��@������ZC�1�c���~��z�=��(�!�;��.���f%'bד�^����'8���?G���x�m�+�bp������o8��:�2;E�5�����=V��Y�z�\�۱�����:""�Iv�q���ҍ�K�B����Pvx׻�!?#�{��U�ńN0h�.�q�Wn�ij���E~'ukr3�������T��P�,����uX�F�,�����޴9��m�;vv�ϡ�o�}�f&kr3Q�s��ݞ�˺T���nKͯ�&wLf+�:�aMnfT�8��#""�d�'|z���N�� �7>x�_	�p�*l�i	����>�إ4+9ѯ�ukr3q���۸�6��?���z�x5Á>c��]Z�Ө�ݢd�����^�[;��Z�S���߇�(�[;q��E�X�����v�|�_�ŵuaH��F9�2�#""r���e>%.Bӏp���S~��g�õ���k/:���[ס�r�����1<����)����^qͤi{��8����f�9���Em[�y�~����_7=Lf+�j>�ؽ����)Z�)���8���[o�|��H�����c���ɋ�u��G�SA[�c2[E�н�p{	O����q:�&蛗/�����]+�pv��gn����I���ǣ�S�����y�K��S�6Q	Or$vLꈈ��i�3n<<Y{�`Ht��Še�GNy����f��e�C>_���?g ��������>�o�t�pt��k��E��!f�)����yڭ'&��c���V-�Zw��ޔ��q:��<���1�#""zhMn�O��bP���%�2���ِض�N^����VwMf+�s��yc=�7�c���'١�Se���uAٻ�S�x������K7<V�}�Z[V��������N�&�n��`&vLꈈ�Z����}�!���'>���)�P�ꍎ�!���r3`ד���k{���#ܺ.��� BE�}����D��)��L�;e-ݠeT�
��)� ����{��&�O^Ĺ[�x~�㨯��J&I#X��:""��|�8��<�����s&�}����{>�/��8���4j�=鲒��F}s+NL�����P�N��n��7��^!��p3#+9ѧ�)e�\غιf�����7�!q#�cRGDD��/�߻�#	�}�>�qJ���n�''>�������OIK�6¨<2�<�n�1x�as\�u�&�����Og����2��Rh�:����DDD�|�=���A�׋��n�&����Lh����۞�^���֮���7�M~F��]=Ϸvz=�-;y�J���Nt��mV}��-"��lŁ��.�/���XG�醍��Wx�xs�xޜO7�K��{��a���*�>6�:"""������rm��E���7����h����ـ*%�u��V��͹W���g����+Q8���uR�671��]���﯆.^�s7��V5皰E��b�*������ۢ�5�tS��H��4��S����8�p��/o�k
�6$$=�;N�$""��)Oӹ�g�N���ߓ�/��r���ـ�]J���{l).�u5�u����Vv6�c��+)�����K٠��/�}+��@V�܈M��)�e(�I1�I|����w���x�N�ӹ����M#�2}.�W>�}W���u�����"B{���je0�����J]�ߚ���sq��]���lG�{Q�&2$�;&uDDD>2Y"sO����~U0"uj�/�G�ur�ٻ������y�X����5�b�]�I��k=}�&o�0��[�9G'i�����:"""r�Te����Q��Gܧac�P6�&�/�y)����1�#"""')׶E�Ó��5�vEl��W׻��I�X{�I�EJ���N�׏"���:"""��s��\�ʛ���ͭX�s#�����BY�GAY�8p�":�ݛ��1��S%y�[����]��8��m4�v���7�T2)���qK"""�g���������� �"l��c�_��&7��/��0�{����u�ZG�д��}o�Y''�J~F��s�Ө�����-&3���<r
�+�q>&��uR���[�0Y��o���F�] �0�#""�o��z��Г��V����Zq��zr�߿_�s���������4j|�ڞ���_�z�����WQ��󾍫a2[�*a����N���66/_�|,н���F�씩7|i��Өq�'/8�4��������E	;N�$""�o�n"m��6>5�6�M�Qc������ƛ�F�^_��y�`&;yj��E����|�V9�vs н��F)v�.X�a��/۠T�-t떩Ϙ�]����B�ǟ��Lꈈ� �6���H�Ey(�ٹA��ʵ�(�db�2��ٟ���^T�<%��C�r+'�ي}�>q{,н�<M���ٻ���;��H���e!"8�Xp�d0�f�T�2"����=A�dfrj5�����`������cMrƐ��(g-r	V0Nl.��E�`ld���ڒ��R_��;�����[?���r�~��<�H����<�'Q�wK�_P!ъ6��  �"�bf�y�g������+�,��mј�#X+y������ӽ:`Ц��X�t��e,�^D���'��x��We4��Eya���F�;9c���P�/��h�� �+����;k�~�"��Ƶz���*��灻�g*<r��:?ҭ	��P�7��;^xY�O�;��������|v��dT��<sf<{�S,����7|�p�$;�����=�Ԗh��Ǵ��c������"v�:  �8�L3O5�)+�k��BvݺV�xP^F�v�yh������*~�a=s�����zC>�Gό*���3򔌑:i*ܼ��3�źw�ۧυ����|5��=q����w�=֕�ЁǶ�ÿo�-�Wh��"
v�:  ����}�����0Wm���Ѝ��<pg�ih�Z��f�7��ĝ_��o�ᕤ'f��3 X�蝹f+/#ݐѺ���z��>l����9k=Z�{ׅWO���
��.p"M}mF3���c�C�?��zC����p�`G� ���'��ւ���I^F�<�=��N��h��%���myံ��i�?[^8`�3�����Ϳ�k̺�x��4'�>�A�g�q�'"�jj��oה��4�y��9}oe͠ue+�Nen�<�(�����k�`G� `�h@�����*��{]o���L�ڞ0&�u:���sa�9=m�C�Dx{�F�9����!��}�v����F�֕��3�6�,�軤����/��3��̙��W<#b���ٜ�	=3�0N$fO5�kK�|��P �4m�����i�� /}垘*]:��ㅗc�s]�
Â]����Q.	�f����HK���~L���-}�7�nH���_?6�㼌th�mT6���j�H��_?�����;��>o\S�[W�b�F��=�ˣQk���hb��hԡ�C�`G� `��_?���n]kȺ�D��;j�+��x��ԉ�K��r0����6W��z^�륦k�<=�n��~����������״��A��������"��W��{oW�_�3���N��hǈ�3gf��ٵ�`��޸Vo?�+������S���#�{�o��b!�5Uj��%=���k���*������I��
��l۷o��X,�jPzz�HFFFA�������1����n 9�ׯGn�|T?`�}ӵ:;�S�a1xx�Z5��ӵO���P�ק�O�j�>'���}�����7]�W?�X�/��$JMY�~��;��f�꺽o��_��l���u�Z=��u��Ks�tq����>�=��>�{n�TinV��nS}M������ڕ�.-TEQ��33��ժ���#�~^�޻I����-U�s>�=C���r0��ݖ����{'㪜�=�ԵEya���F�/�^V��3�uin�vݺV�k��۔�f׈�#�קue+t뵫����ڻs���s׆�{��ׯ/���G�W[�����>���<U�j׭kuནQ��a��H��?��:���Gkt�z �L<��Q����c�o�lІ�Fx�+��<B���:0k�ቾKz�翉�o�?���~�E~k�Jb��tOD5N~��g�[�f��Q��Wն�Ks���e������z=��=�]�.������R}MUܣ�������k�J�|T:��U��ը�jK��Q�o�>�/,WF�~	 @8�=��}ݳ(�h��H�+�9�;�z��Ԟ�V�+[���_ZU�btRl�fk��̜j�oP#좩�:�ξ~տ�ꢙh�4Li��x����%�k��:�I
{~���|X��a�%�<�_�Չ�~}m���Hm��REa��>����5e%:��v�}ӵ1]����O��;�j2����nԺ���gS�Go\���ᾘ]g_����1�~����L��ghT�>���rm��ڶQEyq<�קW;>�ۧ{U��PuiaT���������z��.�^��FO�:uqHwT�Ϩ����麇����;��y�1W���?����~,��-U����Θ2��{'����bj�/˾}��V�T5 ;;�l~~~l�u�<��N�R� &�̽���*SS�JjY�x�+MM����bL�,9#.����[I������g�rS�{�9�	�j��%m�6���;�~���Ж�r�++�-�W���y���:���^C�_EQ�*
��N�]ZS8�SQ��'�U}M՜"1�t����̙��-U�:��v�e�����W���[,��0B�<B�x��a;Z�=��_?jHI��l�Z�}_�'�}�b	,�M�g�ߊV��SϿ~,��Έ>z��o��C|$����3>v�'T���'�YXغ�Z��dF(
��x�xlFp�պ���|?�B)  \Ů��z��]��>������h��I�t�C�����z����W�-���
sD��(O��G��{�^:ܡ��ް�N��V��{o���^~�d�]8��> S�e�1��oI��� A��a�c����k�D�%�u�����1��U����J�7_רS�S
������v��ۧ�E=ʹ�0�J���1������^��{5��,d׭kC���	}󧇴��
U�{ȩg~�֢�����+[��L�N�]ҁ��3F�������P�%�P\�#�tך?�������望�R�����ŢQϤʬ�����������d��D�����=8��!��]�᪢0O��)?ӡue%q�6�f���L��<pgB�v:������#ij{�[V�PEa��T�6$��R�>V�uh'�.i�C��X����5}���=���?���z��	�0�/$��;!��`���4����nB��Z���2?}l�IW_��5.�<�H�J�sT�]���옟c�Xd�X�i��б��9���co{2�軤��^5<�m�*��pF�����vEy�(��at"%3�IS�58�rv�x�u"u*��f/��H����v�?��g��7�r��ict��H֬r���d�Ŀ����gҫ4�'�j�ߍ����?�G��0��A��x=��H�O�����jo|(�s;�]T]�+j}�A�U�QS�5���
2jo|HY�k~E]����}���˞�#) �,�H�W�#�u~�1�R%Q�.�^��v��FB���W�����bڠ|1y���)A��SL��(O��{�*
��o��>�k�����:�w)l��p�G5��U�r�������{����g���{���W,�=c���@@���# O�P��b�U@u��'�-�: 0������oPS�fu����S=3^o����,�W�Oތ9Ѕ��9tV�.�QFf��)�)�[|ۦՋI0�xl�)<���pGB�q�ݓ:��o�>2r;�X=���{Be���[j���Pn�Z��¼�7�Gb�^���7���?c�����ڦIϰ���~`O�UzF�����R�q���X���5�c��O���O�z�Ԝ��7�q��?���"�=[�O;�W���u�����KW���-�/<��EO�-ȵ�,�@�EJȲ3B �Hǹ�*���f~��Ӱ�35J�s���7�����k�[7��z��O���h�!m�Xm��3%I%�*��9tV}���▘��L\Y�d:�wI[^80���b��ׯݯ���}��}4{m�b�!���t�����Ӫ��im�*׉�KZW�bN@���\{tL�n]Z���]j�y����e�k�w�~߫�փ���K��&<����I��ǆ���#�4��{2d:����g���뫵c}�Z�ר�'o��~��j�'�%C ���,����j������%5�>���b�6�u `2-G;UW�F;�W�y�65��MՖ���~��F����yNN���^5�xኛ�;ߩ�K��h�u�<ˬ���w�Q���3��YО׏�dDg��Ѯ�U_S�=ܹ�G�9%5o_�������ۣ=ܩ�����-e+B����:�}�o����GN�jW��9Ӳ��{�Zo�
�W����5��jxxX��.�ᰫxE���	oC0�u���h�%�[7�q�F5l���x�`�t�����n'�k9 ������l��F_x�EO�mͳ[�,ғF�S"��)�\æ�?���͡���fW|�Z]�=���ߑ=-]EJw��n��bY>�)����ۧ{��;ݨ�����K��gm�����s�}G�����j=b������E0:���A�^~�d���=��yL��~x�ywG���،-&��	�{n�F\�P��ٕ�?|����Ј�3c����B�XW�B������p�{|�����*=q% �t�#������d�    IDATu�Z=���q{��/��F����v�QU>���!g�k>?ӡ�wԆ��{��A�=����O]��������Lӛ�Vk�Ƶ:r�wƿ/����S�?]o���3U�����\Ymv�9/�\��UPP���jY,���,;�W��zMh}�l͇ޟ�~�?�Pæ��3[��T�Ԛ����>�:��.�)c�V_|j�)5�|co�U��w�&��	�<jz�jy�>�>����o����%��b���Z��z䛼�1���̑�jU 0w���D�%��{U�n]�g�ݔ���>:������,#.���~L�wLMI��Ji�s�'��[�jM��W��Kou��;qy�tO��G�{B�5��XÕ����w�N��N�vb������{u�T��U�umQ��T�Y����_dL/��j�F\�}t&��	�軤k��gs�jm��SI�s���ܢue+f��RU�-/P���Ϩ$���\�ۯ�wԆ�o����ޫV+?ӡ]���V� �1����{�O�5��j{�Ka�W޲z�v��S-�`�
K箅��[������wy�Z���Ӧ���z���{~�8I�����ڱ�zN�kj;��G��23���w��uz�᫟��~�5�[{��~k{��.��� ��h=~*���k`DMmG�ކ��J]�N�I��^�vISB�=�_O����7̎��=���;�[�s�v�?���t���=�_{^?��~��?~C����]Љ�Kz����tʗ��`��/�����go71=��>o�u|��V�	��k�TQ�7��#��ծ0[\l�Z�-aF�wm\��53�`�e���0O�gmi����ue+tǬ���j]ي9[`��^�k>�aij�qKUy(�Mn�鰇�|^v������E8�7�5���]�=�Iψ�3.j�K�50r�"&�~"Ia��I
��;�ھ�B��������}��k������� ��*��UwcE����	M��e������}���'C0�m��ӄN�
�GZ�T���k�+o�|�e��#w��)Q/�Ow���=�I���1m����m�茜�ۇ��u8�����>����u|�J��3��{/���+����<a��=�Ԉ;�}f�]��.�uI���z��M�}��՞׏���j����[uy삡�-�t� ӡ��]�Ѱˣ����V�B`����eFH#�G2]���>�ᗿ!�{0� L��������Tæ�P��. ��Z��e~}�{R�%��ͻ&imX��>}nj-�+o���JwTMM�="���Q�軤{/��ӽ�v4.Z�~���#�u��aG�"�tO�����a�%�u�IZ��T������-/���u�	��[%L}���g��qy�ďߘq<�����;Bk�z�FC�ئ�������{d��C#d�}����ȭ��}8r�W�=���33�����I�軤�_?�-U塯���P��S��r�x�==��7B#fӧ�N�{�k�v�릿�g~�������N=�ũ_���/���J��^�k1���U$�?���)+w��3c�w*��ڎ��z��nP��݆O�����y�.Co��~�5�/�k�B �PS�fՖ������t��M5j�����%�~�?��m��Hekn��s�9��V��V�#[nט|^��F�~���p%�}��� ו���Iq��3�O��m�EX*�jN�]҉�K3ʾ�*�_���<:����S��{�vzi[�i�{�\hs�`_x���:τ=���^U��8�����K�;TQ�7�ks�+o��׏�9^��U�+[!I3B���9>��h��������R�=�{n��\)|�'�.����{|�s��~�O����zo�{ZJ�N��is���3���SZUPF����;��L���݄}���B�4��)���O��f셧Z�a��^S�����:B �L�7�]#�@��YW�&T9,�i9Z]�Qc�^��=!ɮ@�+�-���IҤU�u�O�ե�C������42�*#.Oد���wΝ����FL�;>�ߍh�'��.��ْ����K��>�Ν�@��(�`�q��ר��t��\Fp�ѷ���z�ڱ�Z�[7�ն�<���@��ŧ�O�m�X�����5u `"�������4�o�w=B2X,6��W���MZ��Z�y9r��]y�*i�my  fc��U~�t�����+��5֫��Sr|����l�E���;��`�Y	�׆G��x�Oޜ*f���@@?OŴ��F_x�%��)�: 0����?�@��Ȝ�d���Q��g�TKs�++�L9y�dO�Qzf�` H���1]g�ٵb�M��s]�kt�3y'���M\��i�[Ԗ����9�k�[7���!U�ݣ.�a�'��ymyiT�	�o��}�D{�/�$�nm��F6[pyp��|�E�b��]�:#�$t/�ͦ�K��
 �Q^����^���Y�Z]�^�44����S�P_��}v��gj}�����WN_'���������F��9uk�f�Z�-i~kTSu ��4��w���C�G�bY4��e�Q8s���>Y'G��d���2r�W^�_���r����'$���� �����ʟ��V����r��S�K���l�Z��R��oC��?Sæ�9A���)�~�ID�.gk��k����y�uF$���/6���>Ց��G�)�B� 蛿����v  ���Pqh��O�d���ҭ�Ϻ�d�ov�+���ۡ��٣���W��Ψ�y-��Nijf��A��'P���J���e���N�   ��o�98��')i�Y����T�a�@@B  @d�wnU�j9ک��|Ֆ�������8w1��A��P�  ,k�?yS��^h�W�7�*�P��Ў�Ւ����k��Eiܻ��_F;zH�  �Gp�dI���"�R� �l�:  "P����?}]���uu}���T燞o�nij�)x?D�����H]æ����Xܲ�Muf���uQ���f  ��L_s5}J��a�G]#j�߬���<�n �A�  ��~�g��f�~�G���
���T7�T�O��q�F�%*�Q�d�X�=$� p�奪-/���~Iu�kTY�0�`�z KK�*),���t�4  �*��r��O���Eu�����R5l�YpS\�K��g|<}ۂ��fǹ�Qm���P����������!� �G��5顏�'s4�cW��snN K9ʊ�A�F=�*��:q��y$��%Ip=]p���������M5j޹M�z��vD�;��F�Z��RÏ~1�܆M5��;�]T��筴���y�R�^k9�*�_W�F��?8����FT����q�5l�	�D�<j~�9�g���HS!)�`��H�9�ػc쟟jMu[$��6D}M� 0��֤���B[s��W�y��*�,����Ue��(-;��X,Y,}�y4t�du��e���r;�WOU�tyB��Z?�DM��U����d:���}3�Nנ3���6��-/Uˣ��dD����T�,�t��~��n����v��ᦢ6n�0��'o2�`Q���E�����: �~߄��㲧�H
�/�2����5��f��$I�w�*v���T���h���Kp���G���G���Q������7�	{�VY����|��TS��<�,�W��m��^z��p;=��<jj;���ҩ X�F�;��� ��X,z����JϋOu���O�m�(����R  ���:����х�?�u��ώԨě�uA뇟�x-P")���v$t~pM^A�C��6J�褩i�;~�3u$Zjp��� ����BO�ӧ[����f�ێs��?M�l��ϓ�  &��%�xro��bm��RB �X{�C����io|hΈMp�g�f�M��n��?}=��*�M���;rUZ�N�׮Sz����a���N��|m��=�(S��S��s��pU�n�}��|o���.OJ�,�{��
gӿނ���h���a��8F ���b�]9�ػ#U�ϳ[�b��u ��Ֆ��Yw�~�G͇ޟ�*����\���q�b�HF�r
oP~�-�)�VNA���t��*\q��ӭ��i���,���٦����p#n�Ey��F����:%��g��CA�#�j���f�����*kKַ�&}���o��a����z���"Q��~���`�kܺaF�hj;Z�4�XGA�#4:��r��׬Յ�:{����UPT�tG��v�,KB��l�������
����N�,9��^K������_v/xn��{�0��o�Y[���:���p2������V|S?��E��'o��TO�����$��~s���TY����#	�XlZY^��kV)?7Sc����Z�η��(]�� ,N���٬�zroA�������v��=�i�A���	̷n���E5�QS�f5�ܦ�㧴c}uhzf���W�f��y갼^��m��iF�R��T�Y�[7�
�DZ�$x�|�۫�v5��>:7}�n��,�G �.����p��Ou$�9�ػ�귶��$F� `Q���-/U��H��ܤzz������v�,�����^�ˋ{�H���¯��n���lAܫ���t��Ia�x�����)������0�E��~k{���k4��O�-��Ƌ�6YfD��u �ht}��9�/���xhZ�BO�����{I	
rd�PY�M���I�:/$�ىڛ�T�UGނ{�Iх���B�nm0�|����)\x�Jiz���BdS�fISm&�0��o���=�b{�7���{�ܧ�6�٭�E	�P �\���5������a"�k��~�&''599)[Z����,�P�z�vh�3.Ir�����}Ѕ�?�;�pQ�T��7]��eO/RM�N�mܺA�;���Xmy�Zp�)��+f7jܺA-��q��r�30[p�{��`�kz�Ii $�Ţ���{���ܧ�6D�������ܧ�ט�����~�t���cM ,ӫ_�X_ڬy�=���@װ�&�~]������5u���rTV�gs��|�	Ym��y'd���3��j�Hz�����t�i=~J�WBَ���/�r�S�5�o}�k>�~�Ѻa�G�o�*�����3^�0F0c1���G�Pˣ���8_�;���q��� `f���zW�]�O���@@����uM?���Z,�JTg�h����}�: X��S�ZP-�ާ��aGꂁ@���9����u����b�)7�B����h��#��s�5��Ž���Q�h��CV�`J��z_]�N5l�	��u��Z+9��p�u���h���צ���8wQ�����nPæ�ｩ�Z?�$��1 `&��Xt�d�;�1��$}˳�۷��j�J������>���o�$�\�g:9�Ju3�����Z��z���4��}5���Rmyi�}��nPS�fu�����9��>���F�mGB#s�jԼs�T��W"j��}�Jݔ�ٌc���O٫bzO�M�����^������ׄ{0�z�d�������  �+���"�|���u���`�����T��Ֆ��=Zc�Xd�Z����U��5�/�I�E7�jK��M  `&�_�"���7����6ը�T�Z�����2�n�������oPæ�?u�i�N_��kg;?�urT�Mv�-����z���eM_)Gza�kpBҙ�� �rE��E�k`$�^���?W��ݡ���~v�װ�35%�J�pS7���/Å�?�  @��Kk�R�5u   �ǚ:    01B    ��    L�P    &f/))Y��������8��=K_q�D�   ,Q��   ���    ��u    `b�:    01B    ��    L�P    &f�t����1U���^��>UϏDFFFaFff��?�����⾧;@�N�7�M    ���/�גnJuC��>���������z�����O�    0\    &fOu ,]��"��ޛ�f   ,i�: 	㷧�U�2��   XҘ~	    &F�    #�   ����   ��T��@C�o3�*=_�P�j��G�   `g?PqW����Oߑt�a���    ��q�u}��[
�.���wT8h�h#�   @�4nݠ�m��n)� ���   @�d:����*��P���Q]�]���P    �wn��e��ڎDu�RtA�;
�    H����j?��5e�-�@T��;�H�S�9�Q_�H]��Ҿ��6    fm������d����:B]n���Wz/|��v    �lL��P���5����:9�Nus    \�V��U���7n�G�'���>5�E����f����T��^��qѰ��F������댮R   ����1�S+W(=}n����ٳ�
������46��ʕE�?�T�~��ϝ�P   `	����a��:k���w���+Q��ΟTaav�����$���    ,~������y���|��~6湉t�R    ���   �T?�E����0R    &�H   �%��%τwƱ4�_��i�}���<�3�kKK�s%B   �%⓮:qp�q�զ��I�	X�t}����<ע�Ң�<s�s�    H ��:I��}�8,�w2��1?�2��zn@}���O    �����#8�'����3#�>���:    01B    ��    L�P   `Q�_q}���4~�M#��b��P   `Q*Z���nKu3�o����wk"=+��	u    ����t�   �"�T���N"�   0���
t�   �I,�`gd��$�!w   �$*Z-�6�\:�����ut�   ���^T�k$�͈Y�ؐ&�u    �������+�͈K��H��ʨc�XS   ��B�����r/B   �Eo)� ���   ���]���P   `�Zʁ.(�`G�   �(��~��]P��({l �k	u    ���T7!��Ƈc��P    &�>u    L�s7��]��d��o�n�:O�׻|j���F�   `j��4�tj����ύ8�=:{�W���S���u    � �ΟVaQ����!��w���+1��R��?!�   X"���;/��?��?��f�
�    ���    ��u    `b��   �d�����8�f�+==mI>W"�   X">麠���Zm*+-������熞�л   @�Y�7XI���S��ay��K⹳1R   ��>>}>��|RO�x�l��   ��1R    a��7�aS�
2�Q뇟���H����0R    !�wnS�����sU���ƭԼs[�[��0R   �p�5l�Q��Sj��/B�ZP�j��vD�.ς��_q�r����ܔ�[m)\ӵ��   0\ݍ���?	vy�z�Ԍ�2T�Z]�ݖ�."~�M'o�[�Y1]O�   �4]�Ψ�_��.�@'�    ,rK5��$B    Xj�Ψ@'Q(   @U�i����;.I�w/X<e�h���T��;	ik��$B   �j�����"THe>�`Wr��K���m0,�I�:    	�q��5���h�V~�Gu_���G�   `���5�1��g?Pq���M���.y���[}�!��P
    SX
�.���p�א{1R    a
2j�T��?Q��H�X㶍��^�a�G-G;���n)����/�]Y';B   ���-/U��� ӡ�Ag(Ե>��j�KC��U�QSQ޼k�b�2"�1�   @B�<z�$����?�$5nݠ��R��T������W�q��mTA�c�=�r�������b�    n��jU�����|����su7VH�������P���4���z?Z�.���w�=6ӵ�:    �N�l9�:V��P]�u����))4�W��1��c�Ih��5>�u�:    Iz�zRܒ��B)    7|�-I�,�m*�c}��?�������nX��6W�f�?޸�u�<�w?�4�g,���F�   `��h\��jz�*�th��ju������.�<@s:�re����F����=۫@�؉��z�l�:    ��8wQ-G;հ�&4'MU�j޹Mu�kTY��+CL    IDAT��������u���
��e��Q��[~�_�Y}����	�   @B4��Mu�h��j�<j=~*T8%8B7�����3�^����;/��?��?��FI�s��    $L���n*>���G�P��S)h��B�K    	S��PS�f�U���Z��j޹-��#u    ���T-�ާ��|Is�T競�T;�Wk�~皺勑:    	Ѽs�*��`��ޜ�+����vD�5��f�3�]�pi|Ɵ��IC��+1R    �ר����EP�����5nݠ��5qmL�I���88��jSYi������zNB�   `Y���B�B�.,��&Z�V�����wqX^��#g�z�l��   H����50�3>>}>��|ROo\�Y,ϝ��:    ���`���ω$ b.B    ����X_}�s��P�26�:    ��8wQ��O�q�5n�0�y���O��U$e9cM   ��h�ɛ�,�WS�f5l�Qǹ��tJ�*��T[^���|u�����6����m�ڏ~%�ߗ�'�Ǒ�K�T�t���,Y���[g��P��   �IA�C��6j�-7�Y_�50��?Q��i��	{}���%�<�l���ޘ�'�E�P   �'82'M�H��-�`o���~	    I:�]���Dz�N�|��vF:�P    
2Qo&��q���0�Z�3*�I�:    	Pwc�Z�/�k~��?5��K%��$B   ��8wQ͇ޏ���	����bmZ��Z�r>J��R    ,Fl>    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01{� s����5=�RZz��2?�_#���T�   0�q�8�У���T7e^�/_V mT"�  `	b�%�666����T7#�˗/���?��    ��:bllL�������������@��   $��SZZZ��2::��&    	G�ò�ZT�e�l�,G�N��   +B���4�ʍ��YRR�����a�   bE�    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &fOu��
3��ސ���C���ci�����|�c��n  �]y��+�R݌��,�zzc�k��
=���X
c�����f  `W��T7!*�:,�>cC���   bŚ:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� �P�f�Ck��_Ia���/v?    V�:,�t}�q�%9��   ă�    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� ���Kg\~����v/    �:,�~}�g¸�\2�^   @�~	    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���S�  rm�Zlܗ{aN��߳#��   ��n�������F\~C��?i��%�n�=����\B   B�2qflB����o֐O��   @�XS    &F�    #�   ���    ��u    `bT��i�|>��n��~�l6eff�b���Y   @R�`J>�O���
�$��+�׫��\�   ��_�nw(��|>MLL��E   @j�`J~�?��   �RE��)�l���   K�����)�u�oZZ����S�"    5(�S�X,������D��%�   ���e�X�p8":�������۸�|θ{   q`�%    �#u0����R݌�ݮ���T7   H(B1>>����T7c�ϧ���T7   H�_"n�5�I���S�    a�C\&���-(UAIy��2��_�Y��n   ��:�er�u����W5��    	��K    01B    ��    L�5u �����A����n  �p\��&D�P ��seU��  ����K    01B    ��    L�P    &F�    #�   ���    ��u    `bl> �jJ��o�ָ�:����g:�t/p%¡? X~u R*7=M5��r��c��e�m)l�yџ  ,?L�    #�   ��1�@T�\�*�՘˘�YΡl��������\.��*��D���ONhrx@���2�{%B�k\�?9��˗��Ŏ4��o[���CǼ^�F�n����}�I�Kc�C�>�x��  ư���r��VZ�����+*��\Y�7�\s��ۍz<�(���u�~-��-��<E7����ؤ���T7e�  a)��:��~(�m����T>0���n���oVVV�$���L�C.�K����$��ŋq?o��d�gFF�._��,� ��lY����<���'�===��'�a��7���v�r�-��?�3�p�*//Waa�$͘&8��������&&&��ե���9sF��c
&�%�,������ٳg�D ��-�PW\\����<��?�?�KA�$##Cw�}�n��v�|��r8��H�|>���kddD:y�~�����O?���"�'  0��`�C�xV�������l|��SFA���Mx������!MK�XȪU����k�ƍ��Ϗ;x,dhhH###�����~�;���Gt]���	  �Pg����r��p�je���z�r�\���]�����٣_�V2��4��U�V�G��͛����@ ��VNq�\�������~��_GF�Db��G}T_��Sڟǎ����z� ��Y�.Uk���Ҕ��-#u���x4::�����s��r:�S%�P��&�dggk���)	s��\.}��gr:�:x�;����
"�'  H�e�R���D���JKKKe3�˥��A�^�z��������'�۽dB]��n�����׾�5egg'tZ`��N�z{{500����/X$�A$��|�ǔ��C ��-�!���C���EVV�#u&�~�����y�������D��$�.q" ���z��'��C�f��t4)�á�������v[(��SPP ����ߖj�4�����	  �[�i�P�x,�Pi ������|G��r�|>_[�ժ��Y,]{�*++����Þ�� B�  H�%�6u��ru����K�>������h�|������)�á�7�>�����"�'� �d�,#��E@�mۦ��~ZYYY�	 A999���T~~��y�egg�=���R��O���b~��'F�'  �:B��E@�|�ISoϑ���믿^iii	"��\;  ��	���������T61p���ʕ+<���������Ą�_.� 2���ҙ3g499�={�h||<�y�Vq�?��O  9B]�|>edd��΄&''5>>����ϛ�������7U��4��]�V��������$�.�Ad``@���w�=/� BN����VSSӼ��  H���b Q�$���g�UVVV[����*++Sqq�{�y�N�����9՟��'  ��X�2�� z��'URRb�"�*,,T^^�jjj�iӦy�+..�Ĩs�{џS�YXXhH ��� �q�}���n[������L��k׮y}a���5�\#)��	  f"�����Z?�pؽǖ�ͦ��2����'�H�3�[�Y�&��	  �"�����򗿬���T7%irrrTRR���r�[���{/�����LX ��u B6nܨ��k�O��k����Z��G,�Oc�  �G�K �Ͷ$�X,Kv'�e-##C;w���MuS��f����D^�W�a�=�Oc�  ̏]��b�hrrrɭ��Z��X,���,��V�|>ߒ�����jݺu���HuSR���D������ׯ���G۟  `~��
Kr��|��n�+==]�E�@@~�?�-C��v��o߾,G����K###ڴi��=��Oc�  ,��0�����˗5>>.��#��*�����5�\�[n�e��"��n�q�q݇��bT ���>�/�$��jbq����+�����)������<]w�u*--��>����  ,�P��
r��r�\��wX\���USS�$�
�"??_N�S_��c����)��  W�O�H
��/�˥��IF����UWWS�押�<�|>�_�>���ϙ��O  pu�:$���._����ȝw޹��~Mg�ٔ���իW+;;;���ϙ��O  pu�:$] ��c:fj��v]{��Y����v��nݺ���?�������X��	  "CiB�������f3������:+oKQk"������J���Ѳ��u��]��Q_G�k ���R�gI;�ͦ�˃�nF�


�f͚e�A�|rrr$I7�pCT�џ��ڟ   2�:��R	vf�j�*
z�#--M���Q]C�/��  �aA�ǣ@ @�$#����p(///�k����ҟ   2�:,���<�iq�+--M>�/�>�?�K ��갨�\.��K"*5�/==]n�;�u`���b�O  ��aQ	r��
)�����jrrRn�{��&''�!   )E�â������NA   ,Z��~�=`�w���Y��X��
��b��D��P�EirrRiii���LuS   ����7�����w���?��X��m$�ٚF��,v%j��P*vQG�W�΋�焯jܽ�(�!,��=lv��E�[���L���oþp�C�2��]j_%G�nD'e,%��&��-r�^P3�(��ΐ�~���4���cZ���{� l&r���Ƃ�~�踽�b�
���Cz��I�;�Y�2�eɿza,\�/�ŗ� �@ۙq� �~��;&udZ�t��:"�K�����n�0��,�?�����x��/����u2��u�_���Ů����,��?h{��X��v���Q-�`�K2�Z:��j����Қ��Y}��E���Ç��Ԅ۷o��1���ʙ�z������.ڛ�����8��gB�Nf�g_�_�y�,c:-Jn�:�ű���Q_�	Hh�� S�d25q���ں�k��L�ϬVVV��imll�b��4G���ʙ�zu�DU�?w�/!��2z �^'s{��S�1�����WǦ�����PZ��Z$v\~I��N����Oj"i6B*�*yo'糰r�^��_�k�o����Bu���y�4I��dV���+3������X��EI�:6�rn�m�İ t��<L�X<G*���e�Ւ�d����d2Y��8�;+w>�ٕ����P��ש��@"��<�H��WǦ���Z �U�s�#e2�ZY�Y���8��鬭e�A��Ζ�8���ʝO""�j� ySǢՎ�r~,$�}<���2�,��èK�D�h�Is���U�۷��~I��|���$""�&YƵ��c!��/�%���x�A����_��IH���U������|����<�̧����=""��TF�:��cqY�|�<�wT�GI?��կx`�L&���|��Ge=�����|�t>��v� pr�β��Q�e�̈e���/�˩�1�#jp������e�iii	{��){�W<�|�t>����A���c�,��~I5A�$��P�VWW1==�g�y�t���.�H������/�z<�s�T4�fao���œ눛��<=��ن�_���{��|�'��}������� G��� 89��cO�  x.mm`:}ng\���h���'�կ{���:^ṕ�7�r��u���W�cj�����ف��_B|-�_\�������9������?r���7��Kptv�s�-�#s[����q�?�v�^Ͽ��焫�K�Z��M&n�<u�#��R��ւ$��K�/-J�=�8Z�c��QM��V��������6|uiccKKK���X]]-�y8�YXYY���|E�Y�o��#��@;:;��4k%�{�����\���y\җ��w����7�:}����������7��<�^��$wv��:  <{��mq\�]����9z��7կ��=�n�w���I�u�f�/>���|/����aDc	�[���-�,N�xsW��v�d���x����W����z�����\���Ww�#��� w�͒?�*�ukFF���K�:6�~�b��s���j�,�쀩�{��arr�����/���}��������|fi5��8:;��߮��;ث~R�5����]�(����w5�I�_K!89O�S�R�G���l�;��0p�&����V) `j~!{��G��;؋xr���G�_wtv�7�Z���:�[��(�����$��������]=��ȅ�#��QJy��d���ϏB[ө�x_[MZKQ��֊,c��w��D�I!�N�ʕ+��d2<x� ���wiT��jm��ZΧ�n�Fpr���7@T��k)����-����!����a���M���ݥ���~���A|-��{GIDɼr+j����|�X��7���U�>'³w�u�f[Y]{Ky�+�'gv\�,-ͭL�F��[+�(��l�JM4�� ࣏>���߰��!�"���I���裏��{�5l���|U�����^�g� �ހۛmE���g�l��M�/l�u;{05��pdnK��݅����b::;�Pc�9y����jUMY������E�Z����lC��mDc���BJ}�k]iε��M[5���TSA�:��������7�7�,��`qq�dR�$d}}?��Op��Q�g��_@pr���C!O�n��$ `oi*�9ów�*���)7��X��.�#sp;{v�KUh�f~����S���yy��L� ��f)	X�����u�N��o���5��K�b����Nv��A���BU��_����������uki5m�嗒(�E��u��3�������D"����w��d2��S5��9�����D���|j;�;��4!pr ��H�^%1+�r�U��H���7���F)��I�J���CM�����Dpr�`���F)J�{����եQi#���MG89�Vn�#sN��7<��q
een2�u[��۟K����L��N<u��%��zݴ]c����ӨKت-�N�ҥKX\\l�����
���055���/Χ�{颱��u��=�})���%�?+�U��(��q{�S/��ei��d�ꏲG�X�����rM�1�����-I���N醩�2��Z*۔�ن�<?�Gm���K������J[.�<�xr]�v�sn.��V�s�����J}�Gc	��b�[k�V�tR"Qݥ\�J�.���X,����A,3z8������O?��������|�'p�fիc��&8:;ؐ��'gԆ��	僃��������V�$N�����Z
���E��q�G�mk;O�S*j�+׷��
�:���E��|�':}b[�47�*�� ����RI+t]9˗�zݴ�:�	�R�0�p8���Y�����O>1z8��x<�믿��9j
�'Q��_��M�N�@���-gw���|M15��=�+����=Ww���J+��BG�7ԏ�t������a�Ȍ|���N����Y����t)	���+{v�G�($=}�]�J}����.1����䌚�z����n[Z��^�6�ba��AJ�2�#�mdY�ݻw��3�`qqKKKFIs.�}}}�Z��/̝�D"Q��jΧs�؞(�P���\  BIDAT�)���\z+[�x�Y�#_82���;7;��t�������#�N
5J�M�	��	��4��f*JI�vJL�%������<�_��]R�YS:izLh:�����;>�����^���|C�p9��1�끫7�<����׭�R���.��:u��!��j�j�8�r� @Ū6�H��X[[C[[[��666 I��կ���s����E��{wnWl�o����G^��ֆ��&���u��9���Kx����o�vyy�}�[XO����p>����
�����+�������������/!�+��b�`o���+�!Kd�[��|�'���qQm�����Q���P��w��_��V���,����hH���hii�7��M������0zH{�'��/����ʾ�\���ػw/�S'�f[v�[K���t�;jz����� "�mб��g��X�� �U��>��/�����X���Ckk+�}�Y�ٳ���T�'����Eww7~�ӟ��+�q>kH|-���f4��c������Sy%"jD�\z"�#o�`��L�	�9ܻw���>[�&3% �������B��7��>rP�6:5��{#b��߷��;RǢF���̸W J>��I���j��ޝ�����~�ݻ�������n��	s�\�����'�|�4	Ƚ{����Y�����i��ԛ��R��WΦS����g�N����v|���|�'tI���ID�a���JkP���q� ��rʤ�L�V*u+++��ں����yҠ������hjj������֭[�����\���nA�$�A���E,þ}�jv>�|���z��&�`Z����o����y�Spr��j�o �'������59H������}�`��{N�@��'{.���\zK�$ˈ�Dd.����[�n��T� &udb{��a�Z__������o���|��)��v��N����x���ҎVVV�L&100��,Q4�@<���g��r�O�WTEs;{�9�=�|�\1�ȱl��Ko!��B��	�G����F\�]�N�;Ҽپ}�Ͻ��V|��1�ȜD���s���cSՌ���G F�}<�:2-A I��àH��h4�'�|_��W��_��Tg���v�����~�3�/�$	w���|�(p��p���D4�P�y�7����BprF��g��?r��.�Ԁ��5t���ߏ����lI�k1&�� tX3b��n\�W#f˹q�(��J��I���je��ܽ{�(��v�Ν;����L&������׿�u|����/~a�X���ԇ����%s�{����;�״>>����%�k���*$v-��]VI���R���Licc��q7J�LX__/z]:���b�Ҩ�I�ڵ��bdd�H���UMF����tbqq����*��,���	�P6��;d\�����X����<G#��ڒ$���_K!�,��B��ē�L,��4�$v�s�^��b�;;�%1XiB0�#E���D#Hg2�WCWWW��'�����'�O>�sss�{��f1r555�駟�7��M<��Sx�����Q�8kkk��Tr>wo7�[ng����-�=}N ����b��U�D3t�6|��>�ݯ��H#������`/<}�-�5���ݲ�3x긚P&n����|ϥׁ�F�$"��Y%1�v����~XVW����7�����.�:2Q��5��$�i�^]�������������a�Z��"�U��455��p����~�iX,ܸq�n��h����q�=t�f�Z�900���fD"ܽ{�n�s��Gf�g�K�#��������	'g*��4D�S*e�/4ѽy��|C����9�Mb�Rj7N��1 ���.���b�<�݈�DT�C���3=A�W�|mgƽ� ���FC �F��2:t�m�Z�=�=A�N�M��/�� �J�����u��˶�6����������9Ċ������!<xP�f4� �w~�w��҂��%ܽ{���H&�XZZ����n��n��'�@WWzzz��ގ��ܾ}��_^^�.�����c_)x�Q���c��/����l���`�����a��=p���l%+pr���o��{�Ww���SO�f��ܫ&�J��WA�:<u��v�A�>'��?�������VFDD��2�ɐ���v���6:��k�xA�i��)X�#S1CB��<�;�{�H$tODdY����YEtuu���v� ��������b�ǿ������}�>��3]ǘ/�L"��m��!]$���OeNͧ�b���>|�>��ABWL��M�:GgGv��?e_�w��f�nU2{K��6�5�#sۖ*�A��Dc��؛mjsV	��A� �+~,��xM�� E%���D���nA@ �:.&ud
� `mm��a4����o�z26����ê!������qUc���C,..b5��M@�������AI���:�sS��Y	-����=�F82�m��lC���o���t@�b�v���Ec	u�`82��tD�`˾�z`D���jY�F>�c���<"2� �9A�s�q�77��*��dRG�cBg�ŧ~�O����֍5H��t&S�18���G��e?���~��}�6���#����@ =��.y���S��Ep>���n�[�89 [U�7���_�xo]n<GgGիb�+�|�yO߲����D��0����߈ʕ��e����VM�}?
��C"z$&ud�zI�������o=��-xʰ���_��aߖ�#��8���(V�W��많j�4��M�g!�X�����;5���bGg���������*B�x7��^Q�2K��7���@��k�臈�:2� �$���ՊL&����F����ެ��T1ng�#�Ԋc�A�z%t���-q�J��\U;���Tٿ�r�!��7�`oiR�\��S�LIGgG�^�Qg[*��Wy5�Y�L��,R��.�߉�1�.������S7�ă�3�7���s"x�8��?�M�n���FШ����\U;�����lSv刊\�X�n>����;ػm)s4�@pr�n^�"x�8<}N�g�����I���z�5��]��=��9�f���}�M������D��_|C���;7��*����	�8z�hL�j!�S4�LB��� D�c��fXͩڮ�&�LWw/Z�h��TZ���*�ĵ�x�����9���8�Z�J�����s�7< �� ³w����X��Q�2�ZO�#�\�~8Q଼hgG]$;��~�G�!�C`�Ɩ9v;{����K�#�gD!Z'�~��TϷ��"�{�������c6϶T��*�� x���:}���۾noi��ϩ���~���^�瑲�AY�`o�m���^1���`u�
�YH���F�n4�|O���A&n �S[�+7��Ύ���t(u4��c���j����_�6E��O�3{�����MGt��f\#*WFV���;eI�N�.��3�*,��=z�>�#�S:�j�;؋���}�u�x89�k�LIr<��R���7���^�c�ów�9�mń�ϩv�՛+?�����f&u�+�ł�����;GD�|�}��m#%		��<|C�e߈���[Yf���;���@��M�JN��Q�j�j��r�\,v���I�J�� �U�Bϭ����X�X�����v�Ճc��s14�.OL�4��� L�y\�������͹��_���S�!�֢���oX��k&L�Hs��$1�#"]){E
-G�7G�~#�v���P<�bdoڪ�߬q�H��L�]�]��>�z�S�u;���P�Z]Wx��w�S��$W��٥�:�+�/�SϑT~F(U�����ȏ�z�5�{ng|C���sh:���F��	&��z�;ث~ �,�MG�+66_�s3&uT1Q��(�2��4R�����r�����rtv pr����_���zc���ܛ&=؛m�A��.u9dprF�O����/�8�ju��FLGgǮޣ�R%�_���q�i����4�k)�.OTe�Bٓ:}b����t����^/��_|��
��]{�������h,ϥ��9�.�ԓ�G!��=puw��ݕ=Sts�|��[��}�m]�`�*�q^}�r[�֫F�A�$X,�AH��l�,�2$IB&���$.�� �J�����u�t��(b�?�����vS������>�]N�s`w)��6L��7�\�u���O�7<�h,���}⮴�w9 �7)1:�"prX���	RDc	]MSI빂��܎�
e?[�+�
=�*U�|��l��Ko�����<}N�g����U�yV�{T:�V��7w�`�_�QX�����2��٣V���H;��|�o�Om+Y���tz.��pd�����g;�uv�]��v�d+�U����N�����}Z��3"&��B3��ԃҡV�_֣��N�7��5?�^{��6ڛmp�oG���sh:�=Ba��g5��V&��z� �1�#"������P��ܮs�P�JwKe����U��[pr��5=.Wi6�׍��g/�S ��<e���/�Sa�� �����+��_���wt�˸�B^[:?�eRGDD5���;�޶?G��f���;؛Mb7�f�S����B|-���͓{�m�YO��3�:(���Q�J(dj~�>'��ܤ3�Q�I�R��=���O��~v�2n�Q:��/�����.O�庺T2�|$=T��?r��~� �h,��郒�j�`�[��N�S���g�s�<0Z��s�'�y��LUc���i�9�������Ҕݧ��Z��p�e�Z�k�܄`RGDD5J�\�$����W����-V��(�l7��	\�	���j�,����ϩ�M�!�@v��w�WӤ.K��YT^_4�@0�:���P?��՘�u�����S[�+���
θ�k��F�O� &uDDT������r�Զc�����vـ����-M[lG�%��^B]���+���[�##�#s������Mh�D24��x#bc�9�z��89�P?B��޻�˸�h�����J$�~Y�x���r|C�r@�w���c��!ttv`�� |��[����&s���e�o�_������j�é��TZ�m3"f���T��z\>���P�V���.O�t�q��J� &u�bRW�����(	�rV�B阨Wg7�X�l� ���%L�����|C��l��=�[��4�<@3P�*���qT�2n�)��L�t5??Q����F �22����+�eYF[[���ˤ��teo�e�gy]7j��r��;��٦&����S�SL�`����^�r��ۆ^�3.��j\-=*������?62<U��?��Ƥ���H�0.��z�J�&� �$""""�0�ƛq�lv���~IT3d�daRT���([\� ; �-�3h�DDDD��R:�I���2�ɐ���pq,^�Ұ�l�㎽�Gd� ��DDDD��R:�I�)�2�eɿza,\�cSǢ)   �vf�+��������L�LE�,��/�0���-_bt<�n�0��s�QG����O�����G_ȸ�˸��5J��3��w\����������x��AU�~�k_S�<�9u5��s�V�&���2��ɛ|ul��'*`��q�1( z<?Շ}ˋp����� �2���D�c���#�U������f��f�1��A�t�,�����u�$��x��饌�ƅ���*�r~,�rn�m��0;""""s�4����j���Ts+���ș4�)$�[�_�� d��XJBW��&���M1�#"""2-:�I��$�3���CF����2�H[$���|�WǦ���Z �U��DDDD��V	� Iݣ��E�~{�Y9?j?{�"���nH��t:���	��={�0.�2n����q�;��L�J�ؑ��2��\)-�ۭ���0�QdY�Ç)$�Ɋ�KE8�2�G���q��Fi�yf����5�:����O?�4�{��w[!^����R�k� .���3�>Al�8��A��bEKKKE�H�_�V�uW�D�q��Fi�yf����%=: `[F"�2~��85z�Ƃ2�0zT�_����ʸ�˸Տk�F�gƭ︕�+���B���c�4z T;��E��/P�e\ƭ��N�h�̸��\z&t@/�$2+H��7n/]��(�H"�ЮY,V,..buuuW�>���(�2.���m[��3��w�R��LꈪOF��!�J�:6�~�b�S���)���n?����q�v5�<3n}�ݭj$t �_U�,��G<��M"""�ZW��`RGTu�(��C>S&�DDDD5��	��������H3�N� &uDU��6_Ǔ�C"""�ZcDB0�#"""""҄	�����Z�p=�|�$����IQcRGTef��	����DDDD�;Lꈪ̔	� ��C """��X� Q�1Y�rn�%H�0zT[�v;���vumkk+�2.�(�Qm�����:�*��}g�=+��BF� ���5zT[Z[[q�ر��J����ʸ�˸�5J��3��w\3��K"���)������ڊ��8��V�'��˸�[y\�4�<3n}�5+&uD|�6:�0zmgƽ���v��_��r�2.�2n�q��h�̸��̸��� 6�L���u��vA�ŧ�!Bſ@6�@v��2.���(�6ό[�qk�:"��3ro]�U��JG�!�"�V+b��2.��X\�4�<3n}ǭL�$B��w'_��f�}g�=0Z͘T�dY�Ç�q�����q�;n-��:"	@�5#1:n�V̖s�.b�Z񈈈�H_L�&�k���j$v-��]VIs�%Q�`RGdJb�rnܥW�}g�=L興���`� jE��q��U��A�M�,��/�P������ͦ(�CG�����7��O����v�e\�58�Qm�����8?jH~Ťn���Q5�2�eɿz~,\���
���C�����
0*�c�K"<g�x����k2��r!\��汶�q�^��#���Q�cRGdb�����uX�c���k��0)*	��^'�� ��p� ٠Q�1�#�������G�f��DDDD��/w�ҽMDDDDDT�d׌�ͤ���i��@DDDDD&$`ʨ�L�J C="""""2��(��ͤ�˙LPF��������C�q-��+u5��X\��ݡ�DDDDDT�2��72>{啡��ũl�x"""""jd2pq�����1�RW����f�""""��&���L��sq,���ֶ��������Y��=��/+�v��|� ������d��$��αfR���q{���L�������|
 ,A
��=�|�����I
    IEND�B`�PK
     Ps�[$7h�!  �!  /   images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     Ps�[
�8b  8b  /   images/a7e3301e-fb46-458d-916f-a05c0bde95f4.png�PNG

   IHDR  �  �   ��O3   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���]l��}����%R�(��(�"mY�-?(˃���S�$]Ңht�:l��u����C�m�i˴�Л]�z�a7	$C
�hs5�r��b9�]�ReZ�����"��8�BQ<�����z��s>�o��/S  �laa�G�"⹈8Px� ����N�*=Z�7�7�^(=   ��.Eę��}��� "6K ��T�  ���=�"�E�gC�     t�LD|:���^8z��J ��� xU�s���C      �ӓ9�?>z��ϖ  M� ��������K�      �!�9��>??���C  `��  <P>�R���w      찱�����=Uz  �� �I�."z��      �TUU���8Qz  �� ��ѣG�^D�.�     `�����ߔ  �"p �����8�s���w      4�_=z���G  �0� x �u��#��;      ��9/�  � p �A�"⟖     РO�����  �iw  :onn�q��     �&���Xz  �4�;  ��R�g�7      𩹹��,=  v�� �N;r��#)�ϖ�     PBUU���  �Iw  :������     Fק���*=  v� �NK)���      JJ)���  `�� 謥����;      JJ)�Å��=�w  �N� �Yu]���      Z�@���K�  �� p ��r���     �6H)���  `'� 褣G�.F��K�      h��.--�(=  �� �N�9��     �6?_z  �/�;  ��s�L�      -��  ��� �E���'K�      h�g���N�  �C� @�,,,<ӥw      ��`0���  �~� �ϔ      �R�Pz   ��;  ]���      Z�������#  `��  tʣ�>�;"�)�     ��R]�~.  �%p �Snܸ�LD���     �bw  :K� @�|��      ������  �!p �k�      wwpaa�åG  �v� ���     ��L�  �w  :c~~���8\z     @��?[z  l�� ��H)=Wz     @���9v�؁�;  �^	� �ӥ      tD������#  �^	� ��;     ��?^z  �+�;  ]ы��Rz     @�|��   �W��  `+���zO�[UUU���݆Q��������p'ccc�k׮�3    �j}}��az�ȑ#�o�����C  `�7  tB]ק�z�~����1111>>����v�~����cccQUU�z=A;���<fggKπV���?O>�d�    [���q�֭�y�f���ō7�ڵkq�ڵ�~�z\�v-rΥ�ދ�~��\D|��  �*  ]�����XLOO���t�߿?���SSS�gOg�     ;dll,���bϞ=q���;>���o��V���ƛo��.]�˗/G]��ݺ���C� @�� ���LLL���|������LLMM��.     `D���8t�P:t�����|�r\�x1.]�/^��7o\�#>Qz   ��;  ]PE�������Ǐ�������     �]�^/>�~�sׯ_�.�믿���zlll\��7B�%G  �V	� h����G��ޭ>_UU;v,�񘙙�4     �199'N��'ND]ױ�����Z���q�����,..>�ꫯ�m�� `;�  ��`08���RJq�ĉ8u�T�ݻ�     `h����������ӧOǕ+W��^�������J#��pD� ��;  ��Rz_����8p �}����      m355SSS��OƵk��ܹs���/�[o�5���9�DD�ǡ�  � �;  ��s~�n__ZZ��~������     莽{�ƩS��ԩSq���x饗��_����}��҇w� `���  `��^_8~�x|���     �6==�>�l|��}�C199��/�����=;��  0,w  Z����c�؝�v�Сx��g#���*     ��ؽ{w<��S��}.>�āv�e����x!  6g. h�7�x㉈�u���>}:z�^Ë      ����8~�x?~<^y�8s�L\�zuۯ�s���x~� �p� h�������gggcvv��9      �{��cii)���ę3gb}}��_#���� ��� �vO��sssM�      (���x�������g�Ɵ�ٟE��^^���  ;�*=   ~�������ɦw      �{��x�gⓟ�dLLL��o=y�ر�a� ��"p ��N�      �6�����?��1;;���ҿu�����  ;A� @���x�N_�r�J�S      �eϞ=�O}*�����|J��C�  �M� @k-...Dľ;}mee��5      �������x���o�q�;  �'p ��r�'��k/^����&�      �RUU�},&''����  t�� �6{��="��_lj     @��޽;������9��GDjf  l�� �6�k�~�ܹXYYij     @�;v,�����ȁ������  �!p ���q<��󱶶��     �V��*:t�gRJw?�  �	� h����������矏����     �j9���SM�  ��� �VUD<������<������-     �k0ĥK���L��Ɇ�  ���K  �;YXXX���[}��W^����|�#����5     �����o����]�I)�� @��� @+UUu�^�+��_���bmmm�      Z���_�o~�[y��� �b�Y ��꺾��="bee%���/����NO     h��^z)����G]�[y|����C��  �%p ��rΏl��޸q#��կ�ٳg���      �s�ʕ��?����7�qO'�����,  �/��  �NRJۺ�~[]���o~3Ο?�=�\LOO��4     ���_���ַ⥗^�ֱ������/��2  �w  ����._�_��W�G�~��111�/     Ш�s\�p!�����������>�S�  `�	� h�	�#������w������O�O<�w�ީ�     �����p�B���k�ꫯ����N��� ��� �:���;��q�������'O���'O��     ����f\�|9.^�.\�����x����  ��  �N��{h�����/��b|�[ߊ�z(N�<��[     ����㭷ފ���������t�R\�|9�n������YYYy��7 �{!p �u��Zl�}꺎s��Źs�b߾}q�ĉ8v�X�ݻ���     F���f\�v-�^�������o��V\�r��������c!p �u�  ��R�ox���8s�L�9s&<KKK�����R�s     ��X[[��7o�͛7�ƍq��ոv�Z\�~=�]�kkk�'���"���  �&p �����^�|��x��7�^�]�v���\������L8p �}�F    �����X__�[�n��������vȾ��7n܈����W��GJ��  �N�9  �Q��������{��^|�{ߋ����bjj*���SSS�o߾����ݻw���x���^     �����9G�9666""b0�����u]���f�����ǃ� ����3d���,�?�Qu]� h%�;  m�Tz�{��:VWWcuu�=���z���\���c����X��J_��W��ٳ�g    r;Dg�\p ���  �Qk.�o���/�hx�(��ݾ~   @+=)"r�!  �NU�  p���     ���\\\\(=  �M� @����싈��;      F�c�  ��	� h�~��z;     @��� ��� �*UU-��      0
RJ���   �&p �m\p     h�#�  ��	� h�;     @3�  ��� ��Y,=      `D/=   �M� @��     �1}�����G  �;	� h���      Fŭ[����   �$p �m\p     hH����  ���  ����̾��*�     `T���  ��� �������      0J\p �m�  �FJi��     �s��   x'�;  ��RZ*�     `ĸ� @�� h���      F̱�H�G  �mw  �d��      ����ѣӥG  �mw  Z#�t��     ��Tz   �&p �5rγ�7      ����  �6�;  m�;     @��  ��� �6�     4��룥7  �mw  Z�رc�1Uz     ��I)�� @k� h������      F�� ��� �
u])�     `D-�   �	� h�^��;     @.� �w  Z!��;     @�=����#   B� @{��     PH]׮� �
w  Z!�,p     (dssS� @+� h��ґ�      FUJI� @+� h�     
� �w  ��w     �r�  ��� ��p�     ��;  � p ���8Tz     �� �
w  �;r��LD�K�      aK�  @�� �v�-=      `�훞��*=  �  ������      0�v�ڵXz  � (.��;     @aUU	� (N� @q9g�     �[*=   �  WU��      �� @qw  ��9.�     �8Zz   � h�;     @y�  �� �6�.=      `��gKo   �;  m p     (,�t��  � �w     ��\p �8�;  mp��       bbfff_�  �6�;  E9rd2"�K�       b||�H�  �6�;  E�z���      ����gKo  `�	� (*�$p     h����  %p �4�;     @KTU%p �(�;  E�u-p     h���l�  �6�;  E����      ���  %p �4�     Z"�|��  F�� ��\p     h����  %p �����      ��;  E	� (��k�;     @{�� @Qw  �r�     �U<�裻K�  `t	� (M�     ���͛�K�  `t	� (M�     �"9���  ]w  J�     �H]�GJo  `t	� (�駟�{K�      �/�z=� (F� @1+++��     �L��w  �� PL���     ���  #p �����      -�Rr� �b�  �$p     h����  #p �����     �}\p ��;  %	�     ��w  �� PL��@�      ����H�G  0��  �R�*�     �16==���  F�� �br�w     �;Tz  �I� @1.�     �SUUӥ7  0��  �s�_z      ?*�$p ��;  ��]p     h'�;  E� (&�$p     h!� (E� @Iw     �v� P�� ���      -T׵� �"�  �ҋ���#      �Q)%�;  E� (�رc�""��     �	� (B� @�n��_z      �I� @w  ���zS�7      ��  !p �����      �%p ��;  E�     Z�PD��#  =w  ���J�     �^c333{K�  `�� ("�,p     h������  =w  �p�     ��RJw  'p ��     �M� @	w  �H)	�     �M� @��  �;     @��u-p �qw  ��     �ޡ�  =w  �H)	�     Z,�t��  F�� �R��      �]M�  ��� P��      �&p �qw  J�     ��� ��	� (E�     �b)%�;  �� PB{K�      ����  ��� и����J�      ��  ��� и��I��     �o��G�]z  �E� @�rΓ�7      ��]�vm��  F�� ��	�     �allL� @��  4N�     ���@� @��  � p     耪����  �h� �8�     ���k� h�� ��      �s� �(�;  %�     : ����  F�� ��UU%p     � � h�� ��      �R� �(�;  ��9�     �A� @��  � p     ���  0Z�  � p     �� h�� ��      �R� �(�;  %�     : 缿�  F�� ����      ��;  M� и���      �s� �(�;  �s�     �3��  �h� P��     ��'J�  `t� (A�     ����S�7  0:�  � p     �]�v	� h�� ��U1^z      [3���  ��� ШÇTz      [SU��  4F� @�RJ��7      �u9g�;  �� �(�;     @������  ��� Ш��1�;     @��� @��  4*�,p     萔�� ��� h��     �C\p �Iw  �;     @�� h�� ���)=      ��K)�/� ��!p �i�      pO��^  #p �Q)���      �'w  #p �iw     �n� ��;  ���Z�     �-w  #p �Q)%�;     @����  4F� @��      �s� ��;  M�     t�� ��� hTJI�     �-{""� �h� Ш���      �R-..�;  !p �Q)���      �7u]O��  �h� �4�=      :&�,p �w  �&p     ��;  M� �4�;     @�� h�� �F���      ������  �h� Ш���     �{\p �w  �6Qz       �&�,p �w  ��;     @�� h�� ��	�     �G� @#�  4M�     �=w  !p �iw     ���9� h�� �&��      �"p �w  3333Qz      ���*�;  �� И~�?^z      �.�,p �w  SU��     ���  4B� @c�      �%p �w  �$p     �&�;  �� И��M�;     @7	� h�� �Ƥ�&Jo      `[�  4B� @cRJ.�     t�� �F� h��     ����  �h� И����      ؖ=�  0�  4��k�;     @7�N�>=Vz  >�;  �I)�*�     ��y�W�Ko  ��'p �1w     �����w  �N� @cr�~l%     @GUU%p `��  4�w     ��J)M��  ��O� @c��     tTJ�w  �N� @c\p     �4�;  C'p �19��      ؞�` p `��  4�w     ��J)	� :�;  �I)��     �]w  �N� @cr�.�     t��  4A� @��      �%p `��  4�w     ���Z� ��	� hLJI�     �Q)%�;  C'p �1)���      �6�;  C'p �19g�     �K� ��	� h��     ��RJ�Ko  ��'p �Iw  ��ha    IDAT   �����w  �N� @��      �R�(� ��� ����Jo      `�\p `��  4&��;     @w	� :�;  M�     t�� ��� �$�;     @G���  �� �&	�     :*�,p `��  4i��       �M� ��	� h��      �%p `��  4I�     �]w  �N� @��      �%p `��  4i��       �M� ��	� hJ?|�	     �ew  ��_z��Z^^���z����ґ�����@UU�1Q����R*��-�@D��Ǜ)�A�y="�kq3���s^����N (f}}�������g      �MUUM-//���; �aUJi<�<����kWD�RJ�rν��w5"���=�9窪V#�f]�k?��r���^�wq0\��_��K�w�"��}�K_ZJ)=]����HD����"b|0DDD�9""RJ?�1�u���V?       �v9�^���Z 5��~x�c�1��v����v㻼���"���nD�\U՟���W~�W�7�yT�w�o��o���깈x6">�r��  �w�      �)�9g��Q2O�������:""���W#�ň��񍺮������_����6����Ω�ҧ"��\D�� �j���     ���ATUUz @������^UU,//�DğD���9��~��^,����[�{��{677&��3񩈘+�	 �K�d     ��s� �f#��"��RJ���|!"��s�r����������:A�~��[�����?�s��`0�k)��қ  ��v     t�`0(= �K�"�SJ�86�����R�������7~�7^/=�������9��9����l���G  ;@�     �}�� `��"�r�?���������?�9��]�v��_��_�Rz\���#"眖��2��Ku]����(�	 �A�s����}�eg]�߳ϝ	I�$Pe����ش�VQ���"(-��ը���ҁ{�3#Jr@��9�d���j��"�6`*��,|c�l�4�,�$& M($s3q^�~�G��I2/����}���]k��������^��]:      [d�; �XT9��F�s�9r�`0�����f�d3�������������L)}M�<  ��4     ���� 0vgG�����8~�����ѣ���׼����2��<��녈�ќ�9��  ��     ��w ���g)���:�+���[��:����ҡ�6S����_\U՞�h�҈�� 0K�     �Ϟ ���~�h4z�`0xw]�����sK�\M���{����)�+"��J� �E�y      ��= �Fu"�������`����~fqq��5iS]pEľ�����
�       �V��t �Y�����}0�^J銥����4)SYp_�Rzm������\  �0��      �g� ��/�9�`0��N��waa�s�C��T�{������WD��s��� �?��	     �~�Ѩt  "���l4����:�������C�KU:�������*"���v �m&�\:      [d� ��rnJ�ʺ�?9_T:̸�~����r4��/+� �S��	     �~&� lKO�9�w0�nJ駖����t��h���s���F���v �mN�     ����  lk/�9|8�"�J�٬V��������9�_���K� ��rΥ#      �E&� l{��i8~`8>�t��h]�}8^RUխ���Y  X?�<      �Ϟ @k<?����`𓥃l�\� 뵲�����9����Y  �8�     ��w �V9?"���F?�w�ރ��G+&���:��M�� �R�y      ��= �VzY�ӹy����*d=�}�}m,��qQ�,  l��N     ���� �Z�����u�����N�����ڵ�@�����  �u9��      آ�hT:  �����~0����՟��zGJ:�m9���o|����@� `z��     �~�|  ��ڵ돮��'�r2ۮ������s�Λ#�y��  0>&�     ��	�  �!���cǎ}���?�t�G�V�~���)�E�SJg `�L�      h?{>  S�))�?ۿ�w�r�mSp����>����8�t  ��w     ��3� `��WU��~����A���~��;���xL�,  L�i      �g� `*�L)�z���]:H�6(��=)�k�C  &�b'     @��� �ZUJ���`pE� %/����F�J�  4#�\:      [4�JG  `�^7�*�X�}0�.�T�? ���     �~�|  �_�y�`0(6ļH�����"���z  �c�;     @��� 03��u��x����2�te�� �,�<      ��P# �ّR�r0,5}�F��ಔҵM^ ���b'     @�;v�t  ��?��+�����6yM  �w     ���� 0sRD��.x#)��߿���;#����  �~,v     ��= ��ԩ��7����k�b/����\PU�{"b~�� `���	     �~u]��  @9�s������I_k�����]�N���I^        �<C�  f�W��ͽweee�$/2��{�9u:�_��gL�  ���N        h�g��ͽ#�&u��������dR� �]�     گ���  (,����p�<��O������-��I�        (C� �5o�9���ྲ�rAD�fD̍��  ��	�      �g� �5U��k���x�'��zU��y{J���</  �g�     ����  p\J��UU���덵�>֓���w#���<'        �=�u]:  �HJ�[�=�ܥq�sl��`����q� ��b�     @��� ��RJoX뒏�X
��]w�Y����9�� 0},v       �T�����3�����~�ȑ+"�_��\        ��T�u�  lO_}����8N���p8|fD,�!  S�w     ��Sp �TRJ{����z�-ܯ���9�GĎ� `�)�       �T���_�����-�R�}uu�?F�3�r        �Lp ��y���Wn��.�_s�5O�9_��� 0;Lp     h?w  ��u+++l��M܏;֏��7{<  �E�     ����  ����z�f�T�}���ύ���E          �N)���:����{UU�#"m�X        ���. �vHUU]�s�p�|���`��ƍ �l��	     �~�|  ؀��n�m��~�7t"��7z           fKJ�M�^on#�l��~�w�<".�P*  ���s�      l�	�  l�����d#���6�}�F @��;     �4Pp `~f#S��]p��;~0"���H  �<w     ���� �&<u׮]�a�_^W�}mz��l:  3/�T:      [�� �f�_��I?�u�o����o)  3��*     �O� �Mz�Z'���UpO)-n-        0�� ؤ��|���p�����-� `�Y�     ��}  ،�ҿ���g쥟���s�=�H  �2�      ���  �UU���-����\/["  f��N     ��P�u�  �T������)���>77���1�T        @k)� �;:�Ώ���,��S���          ��X�9���S�8���D        Z�w  �����N��)�u]�|2y           �a�쪟�����/�X           f�K����O��I�v�zaD�h$        �urΥ#  �~�u]��d����s�d�y           �a'�?�����Ή�N<           3)��=�~��G���������1�H*           fN������G����{J�I        �Nιt  �DUU/x�{�|#���<  lUJ�t        `�9� ���b��
����9���          �z�`0���xX�����l           f�N|Q=��om.           �,��-'�~��~�7tRJ��|$  fAJ�t        `�y�7��9�⡂�w��8�H$           f�y��v�3���N����          `���겟Xp��Y           �a)������g� ��H)��      ��KG  `�\|�UD�u�]w^D��bq           �UO�ꪫΏX+�>|��0R          ����;w>+b���*          �6��6b���R��e�  0�R��      �i�s. ����k�����f `�)�        ��Rzz�?LpWp          ���+++�"�+
� `�yT%        p_y�uםW���=�t        �6 `R>�UU]�O* ��R*        �ƪ�zR�Rzb�         @;�� ���u��*"�          (�UD\P:           �-���*"�Q�   L��R�        �6�s~\�+        h��s�  L����;           ��㪈xl�           ̼�V9�sK�  `���JG      `��  0A�V)��S  0�,t        g��J)�,� ���        ���*�l�;        �. 0A;���+� ��g�     `:�� `�vTq�t
  �_UU�#      0
�  L��*�t�t
  ���N     ��`� �	:Z圏�N ����	        ���*�l�;  ��     0��  0AG���j�  L?�      ӡ���  �^�W��)  �~
�      ���  ��R�b_, ��g�     `:�� `Rr�_4� �FX�        N'���*"�_�   L?w     ��`� �II)}���ϖ ����	     0��  0)9绪���t  ���N     ��`� �	��J)�Y:  ��B'     �t�� �����4� �FX�        N'�|Wu����J `�)�     L�>  L�h4��ڷo߽�w��  0�,t     �_Jɾ  ��}���[���T�(  L=�      �g� �I�9*"���H)�U�8  L;��        ���W9�O�� ������_     `[3� �	�ˈ�����Y  �v;     �Ϟ  ��s�h�Z���ѣ�DD.� ��f�     ����  0!ynn�ck�}����.	 ��f�     ����  0!���𥈵���[
� `X�        N����P�=���2Y        �60� �	���?N,��L  fAUUg�      ۚ=  &�.�Cw���w��"�`�8  L=�<      �Ϟ  ������_<Tp��z�RJ.�	 �ig�     ����  0�����g����<  ���        �I�ɉ/Vp����� ��Pp     h?{>  �[J��'�~X�}yy�/"�F 0,v     ��=  ��s������7VpO)���F# 0��:�      ��� �����:�9Y����        ���;  �s~�#�{T�}uu��#��F 03:�N�      l��� 0.)�C9�?x�������z��w  ��b'     @�j ���߻������j�k�y  �1
�      �R* �)�R:ig��-�����E��D 0S�     ��w  �!�t����?�g'm�z�C��&�
 ����     �~&� 0u]�{yy���}vʖQJ魓� ��Qp     h?{>  ��)�ꧼ�\\\�����$�  0{L�      h?w  ��o�����Mp�)��O&  ���锎      �)� 0oI)�S}x�;Δ�["���# 0sLp     h?w  ��hUUo=�N{ǹ��xWD�8�H  �$�     �O� �-�����)��3�|���  0�,v     ���F  lEJ���3�����?>�D  ̬�R�      l�=  ��楥�������Ѽf�a  �q�y      ���� ���|i]w�^x��-� `���     �~
�  lҧWWWߵ�/����K/��V��	 �Yf�     ����  �9�_��z����u�q��Ͽ#"n�l(  f��N     ����^  6*�t����������[F�_~�є�U�� ��Sp     h�N�S:  ���^�wd�_�P���O~�/�?��L  �:w     ��3� ������[6r��ZF�^z�(�t��2 ����<     ��P#  6"����/���F���g��}wD|x�� 0��     گ�锎  @{�����=h�R�/"�&� `F)�     ���  �)G�rJiÝ�Mܻ��"�77s,  ��D     �v����� `���~c�s�a����z1"����  �=      �M� �u8�Rڳك7}ǹgϞ��9�a�� 0{Lp     h7w  �$�����Ż6{���8�;�k"��[9  ��w     �vSp �>>??�VN��;��/��hJ�#��V� �l��	     �n�{  8�c�c�_~����[��\ZZ�hJ�ꭞ ����tJG      `<� ��t����Փ��O*w��qeD|b� `zY�     h7�  8�������8�X
�w�>�s�ш��8y  ��O     �v���ԍ  �.Gs�?�����8N6�;���古�^7�� 0}Lp     h7w  N������q�l�w�|SD��8�	 ��0�     ��� x�]x�+�<�X�8{�^=�~8"�0�� 0Lp     h7�=  �����.����8O:�?�ܻw�9�E�X� �~&z      ��'� ��������{�O<������SJWN��  ��O     �v�� ���v���O�������Ɯ�oM��  ��O     �v��^  "�w����4��O�3���:���['u  �ł'     @���͕�  @Y��ܹ�R��&�0ڽ{�}�N�E��I^ �v0�     ����  ̴{�~��ݻ��E&>BsaaᶈxaD�?�k ����     �n�� 0�H)}��={>=�5r���vo����Q� `{��	     �n ̤QD�����MM\���Q�۽1"~,"rS� `{��J     �v�� 0srD��Z�����v�o�9���k �}X�     h7�=  3g_��}s�l�����|]����.  �UU㷟      ����\�  4��nw�-�0Z^^����ĵ (�D     �v�� 0r΃n����.6Bsyyy9"^_��  4ς'     @�yb/ �Lؿ��.��g�۽2缯d  ���     �^UUEJ�t  &(����v���P�O*���WRJ��Kg `��     ��^ �T�)�奥���ˋ�#"���)������  09Y	     �^
�  S�X��'�����Dl��{D���ү��^��� �dX�     h/{=  S��������_)�mSp��XZZ�ú��w�� ��Y�     h�����  �;���n����AN��
�{��e�ΝGćJg `��     ګ��]� �ͻ���|ݞ={n)䑶�]��ݻ�޹s�wD��Jg `|�     ��^ �������maa�s���̶}n��ݻG������)�AD�H\�    IDATU:  [c�     ����m� ��9�s�.//�b� ��-'��hyy���ƈ�t�,  l��V     ��aF  �R�#���۽�т�{DĞ={n9v�س#���Y  �<��      �e� @k�x���g,--�T:�z��A���7"�w8^�s�>"W:  ��     �^ss�� ��"b���t��hݟU.--�+"�6"��t  6F�     ����  �������m+�G�����vo_]]}~D�:"VK� `}<�     ��� Za5"^����M���]:�f���A�^���kWVV���t������ ��yl%     @{)� l{���v�����o�ݻ��q�`0xID\O*	 �S0�     ��� ��;#�U�n���A�ajF�n����է��E���y  x4��      �e� `{I)J)��F�����1�O���E���W_�ku]_?ST� h;��      �e� `����,,,�V:̸MU�����Ż"��~���RJWD�K#"� 0���     ���; ��������vo.dR���~�������K���3s�?��� 0�����     `�)� ����~vqq��K���h---�E<XtND��9�8"� hXUU�R��s�(      l��; @���{"b����M��4e&
�ǭ��}Ɂ�Z���r�?g�� 0K����hT:      �i�  �9����iaaᓥ�4m&�:>�:p������҈xUD\T8 �L���Sp     h!� &��9��r�Yg�e���w�S�L܏[XX�RD������9�����.��F�Y�� L-�      �d�; �D��߫���C�}���ե��3"�~>8p��c�����e���ʦ �.
�      �� 0V7G�;v����Y��~2�:am���Fį��D�Kr�/N)����� �"�      �d� `KF9���RzOD���vo/h�r�yk�8"��`0��ҋr���_V6 @;Y�     h'�<  ��������rο���|O�@m�s����=�x[�׫�9�g���=�������xlр  -��x(     @�ر�t ���K������СC��zu�Pm��	k�h����s��k��꺮����礔.���"�ܢA �!�=      ��> �����9�RU�MUU}�կ~�_��r�`m�s�~?��󶈈^�W���_u�ر����RJO�������'� �L2�     ��<� �AG#�o#�o"�orΟ��O���}��{����Jd�:
��������<⳹��?��ǎ{|J�	)�'�u��qVUU��9?&"Ύ��a
�vw,"��.�9?����D�h���	?D�߯� 3�ȑ#�O*�     ���9�N<8� fI'"��:�:᧳��s�{;"b5">Q #�s(�r�联���u�ň8\U�=9���??77w����{w��;V �LSp/`��sk?  3�.xgD|�      l�[��֟���?�K�  `�U�  0s(      �����P�  L?w  ����      �qw�}�}  &N� �F�-|     �ϑ�8V:  �O� ��=P:       f� �F(� Ш��Lp     h�C�  0� hT�Y�     �eRJ&� �w  �f�     �er��x  h��;  M3�     �eRJ�Jg  `6(� Ш���;     @˘� @S� h��O     ��1� �F(� ШN�c�;     @�b @#� h��W     ��=  �� @�Lp     h�C�  0� h��      �c� �F(� Ш��	�      �c�;  �Pp �Q9g�=      ��  �Pp �Q���w     ��Qp �
�  4j~~^�     �}� h��;  �:��-~     �ϡ�  �
�  4��[o=��9      �C�  h��;  %.      �1� �F(� P�	      -�s�� @#� (�(     @��� �
�  �`     �ERJ��3  0� (���      X?w  ��� @	�J      `������  �lPp ��     Z����7� �F(� P��;     @{�{���  �Pp ��C�      �n�"�. �٠� @	&|      ����  �
�  4.�d�;     @{��  ��Pp ��     �C� ��(� P�	�      �� @c� h\]�&�     �DJ�`�  �w  J0�     �%r�&� �w  J0�     �=� h��;  %��     �K  `v(� и��	�      -�R2� ��(� P��;     @K�u�� @c� (�P�       ��	�  4I� �ƥ�Lp     hw  �� @	&�     �DJ�`�  �w  ��tLp     h���Mp �1
�  4n׮]
�      -�RRp �1
�  4��[o=�J�      ��RJKg  `v(� Pʡ�      8���Lp �1
�  �r�       ���Ç� h��;  ���     �sssKg  `v(� P�	�      �_���~���!  �
�  �b�;  ��ۻ�9ӳ������n�7Yd��,k,Y���@H��D�!eI@BBd�a�r��d�'$�x�v������~� ��C���y��kg�]��޼���.   �w��ҲG  �>�  dq�     �w�  �^�  d�     ��N�   ֋� �,��      �J.� �Tw  ���     й�� �Tw  Rx3     �����  ��;  )�q���     ����;  K%p  ED�     :�Z��� ��"p  ��     ��5� X*�;  )�q�     t."�  ,�� �.�     L���  ��;  )�      �s� �e� �b�ϲ7      �r�5�;  K%p  ��      ������  �z� �b�;     @��qt� ��� ����w     ���� �R	� H�����2f�      ��Ο?�;  K%p  �XJ��=     �:���z�= ��"p  ӝ�      ����  ��;  �>�      �d  `�� ��;     @�"B� ��	� �$p     �Tk�v�  ֏� �Lw     �N��\p `��  d�     t*"\p `��  �i�	�     ��;  K'p  MD�     :w  �N� @�;     @�Zk��7  �~�  ����      <��  d� ��w     �~�� @�;  i�      ���w  �N� @�q�      ��A� ��	� H�;     @����ogo  `�� HSk�     tjcc�w  �N� @�Ǐ�     �Ԯ^��Y�  ֏� �4��̛�      }�[J9� ��� �f{{���Ҳw      �7�  ���  d:*���     �� H!p  ���      |�� �w  �d      ��  �� ��w     ��� H!p  ��     �?w  R� �&p     �� �w  �	�     �#p  �� �T�5�;     @gZkw  R� H�      ��;  )�  �r�     �?�8
� H!p  U�U�     ЙǏ� H!p  ��      �y|�֭;�#  XOw  R��(p     �˭RJ� �z� �j6�	�     �r3{   �K� @���#�;     @_�  �� ��_���     �/w  �� Hu���ǥ���;      �w  �� �+�      �� �F� @�      �� �F� @�      �� �F� @�֚�     �w  �� Hw     �N���  �� ��;     @'�  d� ��w     �~��(p  �� �t����      �֗����do  `}	� H�Zs�     ��.]z�= ��%p  ]�U�     Ё���� ��&p  ]k�V�      Ji����  �z� ��@      ���  �z� ��;     @�  �� ����X�     Ё֚� �Tw  �-�{���;      �]D� H%p ���      ������  �z� Ћ��      ��8�.� �J� @/�      �j�w  R	� ��~�      �u���)p  �� �.��\p     �������#  Xow  z!p     ��z;  ��  t��*p     H�Z� �N� @/�      �"b/{  � �BD�go      Xs.� �N� @/\p     H�Z� �N� @/�      �"B� @:�;  ]��
�     	� �� �.\�z�v)�({     ���q/{  � �E+��&{     ������ @:�;  =��=      `]mnn
� H'p �'w     �/_�|�=  �  �d?{      ��r� �.� ��      	Zkw  � p �'w     �!p �w  z"p     ȱ�=   J� ��;     @�֚�  tA� @O��      ���� ��;  ���)     @�k�  ��;  9::�     $h�ͳ7  @)w  �"p     H0���  tA� @7�ŽR���      k�p�X��  �� �+�      Kۥ���  J� ��;     �r]�   �� ��;     �����  �sw  ��Z�     ,��  tC� @W"B�     �\.� ��;  ]�     ,�� �n� ��8�w     �庖=   >'p �+���     `��� @7�  te�     ��p�X��  �� Е�
�     �g^Ji�#  �sw  �r�ƍ���{�;      �AD̳7  ���  ��z�      �u�Z� ��;  =Zd      Xײ  ���  �h/{      ��p� ��� �Nk�w     ��� ��;  ݉�;     �r\�   O� �#�;     ��� @W�  t��&p     8{����F�  x�� ��D��     ���K)-{  <M� @wj�w     �3��  �,�;  ��q;{     ��k�meo  �g	� ������Rʭ�      +���  �,�;  ��      g("�  tG� @�Zkw     �3�Z���  �%p �Wײ      ��Z��  tG� @�j���      V��|>��  �� Х��<{     �
�*���#  �Yw  z%p     8;�f  ��� Ыk�      V�� �.	� �����     ��� �� �.-�{����;      VQk�r�  x�;  ݊�y�     �UTk�u�  x�;  �j�	�     ����� �.	� �ٵ�      +ho�N�  x�;  =��      ��~�=   ^d�=   ^b�Z+��� /t���rpp�=���ѣ2�c�    �Rk-E� @��  t��6?<<�]������׳g@��Ey��a�    ��/}��R>��  /R�  ���֮eo      X5�V� �� �n	�     N�� �n	� ������Z���      �""������  �"w  z��      �
"��Rv����do �� е����      �
��d�  ��� е��V�     �U�����  �2w  �VkuE     �<��.p �kw  ����     `DD��;  ]� е�l�MV     �S�$p�8{  ��� ��=z��'_�	     �[���������  /#p �k7nܸ�;      V�/J)-{  ��� �)pI     �-DD��^��  �"p �{�֭�      S�����  �*w  ��Z�${     ���ZK)���  �*w  �7�k"      o��Zj�>s �{w  �7�k"      o!"������;  �U�  tocc�W�=     `�"�J)c�  x�;  ݻr��^��a�     ������  pw  ��E�N�     �)�����G�;  �$�  L�V�      �)� 0%w  &�����      Smss�g�;  �$�  L�0���      0E����u;{  ��� ���yDdo      ��Z�G�  ��  L�0��     ���(�0|��  NJ� �$���Ok���w      LI����x1{  ��� ��8��ne�      ��Zk���d�  ��� 0�q�     �)�����ٹ��  NJ� �d��Q�     �)q� ��� 0%��     �$"��Z��  ^�: �ɨ�
�     N���*�w  ��P 0��엵�1{     ��Z˹s�~��  ^�� �����zW�w      LA�u�ʕ+��;  �u� ��a~��     `
�a�Q�  x]w  �惈��      еZk)��w�  x]w  &����'o�     ���w  &G �������     ��axx���w  ��R 0)����Z���      =����ҥK��w  ��� 05���Q�     �^ED��~/{  �	�;  �DD�     �.�P"���;  �M� ����Ok�(     �<�0���d�  �7�
 `���     <_D\��緲w  ��P 09���G�0<��     Л�(����  oJ� ��\�x�q����      ����R���  oJ� �$E�k�8     �ak����  oJ �$��~$p     �]�0|o>�?��  oJ �$���'_�	     @)��g'���  oC� �$]�v�r�u?{     @/�a(�n�  xw  ��E�k�H     PJ)�ֽ���f�  ��� `���     �����RJ��  oC �d�����0d�      H7��J)�;�;  �m	� ������#� {     @�Z��W����w  ��� 0e���Z=�     ��Z�a�ǋ/>��  oK	 ��E�{�0d�      H�䳒�d�  �� p `�Zk��;     ��f���Rʻ�;  �4(�  ����݋�0lg�      �Pk-�͝����[  �4� ��VJ��'_�	     �Vf�Y���g�  ��"p `���     XG�0�r{{��;  �� X��� {     �2=������o� �� p `�vvv�R��V��     ��������7�w  �iR  �*�9�Ͳ7      ,E����wׯ__do ��$p `%Dķ�a���     `f��8���d�  ��&p `%���܏����#.     ��"��f�o���}��  N�� ��Qk��l6˞     p�666Jk�w  �Y� �2���{��̥     `eED���������-  p�  ���Z�+W�    �U���qw�?��  gE� �J�����l6�u�     ����c�  �IDAT6C��/���v�  8+w  V�q��/�a��     p�Ν;�㝝����  gI� ��������s��-{     �i����Mk�OJ)��[  �,	� XE-"�l6���     �f��݈���b�i�  8kw  V����s���iq�     ���l�����{{{?��  � p `e���~kss�K)7��      ��Z��l������������{  `Yf�  �,-�*�|�TJ���X=<x��͛���:�[Jy�=  ���ZJN�Ν���͎�����f��8����儍Gk���x*��g�M�^��~ "�k��[��Q)�=��G���q)�w��a~�5#�?���Xk�=����s�  �v���R�y�L    IEND�B`�PK
     Ps�['�Y��  �  /   images/4bf63cb1-3675-4452-8ab6-1403298522d5.png�PNG

   IHDR   d      X�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  SIDATx���KA�_�&�Ҕj�PZL-1����?�7O=x��[�ދ'�{�xl=x#"�P"�ɖ�T�[b�&���ݢv��xa��o�;o�f&
I ��ё��v��F��5�M������Yj�ۧ�����ZZZ��v�����$��\�v�T�)�Q�Z���?�;r�V�B�x�1E����� &M6���������FM�0��UUu���[�;<<$��K�Z�L���B�@�LF/_7Ft�o}<YB��.��Ȉ�8��p�\�b�hY��|>D�A=�\����l!�>����=�����y�ϐ!v�[V�������ѓ�=��a��ò���;�\��)�mr.�&�277'�A,C�d�����ƉpF��F)�uI�
f�`���(_���X��N�ǐ�v�����4�q$����"�q�	T���.�[�$�F���E��:MdW���a��n��4�'�b�to���f�����<��.�1L� �=�%n ���r�F�I�wQR�V!��{�G"[��Zbh_+���Ol3$����%��;�'���������(Ϥ'�0�j�����U�99��Xf{Ƕk�Cv�8����
�����v� ;;;����W��t)�x�D�ֱLmll ��PX���ښ^����.�P̂(p$mP!��/eqqQh��!Fk�\��jX� 8.1�d�"��{�n��Il�~�&#��r���>�t�z�JE���>��-��ޞ^�n�a<I��+nDE#E������O�[V�0��T*u�pZl�k'���UV�R1�n�y0q�<��>���$���I�"�t}�4���������J�u�    IEND�B`�PK
     Ps�[9&��ސ ސ /   images/b01488b3-8551-4b4c-b09f-2812c4acc168.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  ��IDATx��y�m�Y��=�s����n�$�I��� �1���0(. U�D�	W���T��
�+�JR�#�B�Bʩr*�+�	6�6�hh���o���{�=��o\{�s�{��H�}��^����a���^��}���p8��N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p��h=��?���0>"�����0<�޿T�fS���bߔC�S��)�P��� ����e�C����0x`(gu��]� �(�X�_��y�����<�����:�=B�6�n���7�k���S�#�F�����S�1-0��!$�n<���!��`(���x~��'�����'�G�iX�s�q�8����:��q)v$7���GY4��1@�a�נ��?`�3��`�G1���3�����|��(��P�����ʢ⯥�(e#�]����eXq���8�W��&��n��g�^6���"t�����fq}�4��/������;�M8ٟ�瞀����O�(��p�$���yL��&�PA���-BꊠDO
����La(Z��g<�0Ȝ������I}"ţM-�I���\�C��x1D<���ؾ�,�"���U��_����>��W�7O��'��W�c7��－�y�������� R����g�H�7B$֌���fd�I���*��@�7%t2�}��|�W&��:	"!j�X�c$~���(�#l�bn:n��kuh�$���y,g~Y�����?o��oCc�F���YBY���c��pp��5�[Bo�^��|�vs'Oު7�/��>������?�R�UH�oA*|��Ȉ��;��0G��HDM��3	'}T�v:�lRO /o�g���q"�ٕ7���Zk��'�]�z�����>�=u�*Y���(��TAQ�ş�Y��+�>9����x��py�W���~z�Əݽ����!v_��Ư��T�8��:�e�����P��'mQfDr�^��L�l��0�Kll@��,�&���Mu�1$��َ'R��ь��ND[&�k_�Ch���{=m
��a�X>���D�.�-*Mź(ʋ0;x�<{aYՇЬϡ]�C}p"���w��.^䟛faqt\��_X޹���߆��N4���؟�l��)�u����	=z���S�(�a��<�ؓ	�I=�p{�|�\�b����d�X�]#y_¦_�r��
ϵCR�c�z��MQ�]�i�Ԋ�ҡ��B�d���U������>��!��������~���~i�6_��)��;��.�K��O"W�����ߌ���)��}w#v-���]�$oB!�3� �g]�0���zg�"Z�� +*�&�_
���D�7E,���dGeO>�<{�˘�b@��|�Z�->�	���2���3h��iQ�!��$��ֳ�����_����� ycI�8�u�X�7�N���g?K����N��=��au��hѾ?��si�n�^X��"7�B�L�=��T�t�2�ĉt�
�&�υ�)�moz�G�'���}�B�Y�MS��-��;G}	�8�[\�C? Q� ��hU�P��]ࢤ+ ����:̠�j<���&4q��0o�;��{����W~����?����O���_���p�Ʊ�l�B^-�����G��}ٛ�z�����}�M���[#-���S�dN2eM��@Y��q�o�U��	�D�!LB�&����׳+s*/�GCf"/���*���ҔD/(8�4�ʲck�,��>��~����
��?E�����^���������_trl/��ާ�Y��)Q�=�������8��Cw���+=� ;&Q
��ԍy��.T7�2�q͚�LD��1�<yF7�����~6�ϳw�>Ç�cH����Bo���*{�$�t}M۲�>�WpPԜ�W��y��Zz���",XC���� �1�z��_~���������o|ӗ���_ï�*@�� ���|�����c��ɧ��}�bx��x�[/����E���4ϴ�͢�܁�d>��B���OT��s�|������T{yޡ�� I=Q��š8LeQd<��s��)M��v`�<���Y��c��kfܐ�-J1�3=Z&(�Bq���1��W���Q��A�gB���a�������������z�w�m�\܆fyN�z���n	}u�.�G7`}����3T[ᤆ�����G���}�Z�5S�ؔ���i�T�2�坑�w�'#�4e��N�d�����Q���s:�l�����A��c��(���s�G�������5�����=���-|\C�⍞�u�x�u��妄��jg�c��?���4|?.�_/����o�\U�G��ߋo���!�m�bq�&8��?./ɥ8}xx���bh\��{��~�����v}�n�7�A���j������	�4x2RzT���e���8T�Q�D�/�EٱZCs8��CR��A1G%H��rb;��l�d	[ϛL�OL���А���E���/�}�(
s�� m��#��b�F$��*�j���gc,�������^J��1�Q�'/��Q?I���g f�NN��}��Ї����'��_V�_xk�^�N��}kHm�3�'�h�B��$nN�	�svy�y;2��K[�r������F�<�t��B�� l_�&��ߨ��]��ʱ�4��;�i�Z|o�E��P���z*_KhŇ�-��H�ҕP�ڢa�K���b����g��{CQ�VY��)��o�bY-u��Q8�AY�9�@�7����ڥ� 	7�>����n6'i迹o7�o��˴z[��<�6�e�������	z^)���G�60l6h��Tw��xǖ8���F?�Y�%�n�A�$�Y��s��4|���i4L�dː7b�g�C ��Kz_�qx�z�� �TbB9E5C%�������v��墨>Z��C��̓�%~�N�i뻟���m����S��$��K����@<8^\���7�����o}s�̆�eDm�Yr�h�V��G���K�ʄ5�dYm��YcM����!�v7M�8M��ɀ/�y
�&|O��k�U�Q�je��"f&U	��r�kv�G=�.UH��hS͵�TO�%��~#�E���))Ѯ/C�>���7T��+c5��b���P����Z�Z]U/���;�=��Ւ�+�����.U�5���
{���E1G���gp�[����a�~6���0���$^�+$�5��Hͮ�'�S\����f��ް�=�h��:4С�,��Sw��s�2�
K�� �x�2����4c���ו-{���L,�P�����Q~����N�1�8����$��
�����TTo��_L}�eU}b�����8T���'O\l���3Y�A؃d���_� �,��&4��A��g!��*RW�0�Q�S�Z�du)��u�gk��S�q)M����m��+�l���
$�d�v�ZP6�'V|B�.���Z���J�8U����)X����.�"zVf�R�D"�Ԅ��ǥ�0P(fhЮGB_�tX�(V]�Gl�B[?W_�ٷB��nS�ˡ]��jV}�(��P�m.���%
�ri����r8�]�..�Cc�������e��ě�Q`<>��������ƾY>74�[�YU�6�@"�e[��_Ė��+�=Z�d t��54���{�k��}�V�F���뇒������5k(�K��U�q��'Ƥ\<&��Ul"W/F�}�O^�Tc�e7K��*s���à�����!s��9�/�e��{YY*��G�}kY�~��_[����Vy��G�7�������?�g����˟�xYΟ���c�o2u�[ 6���:��Բ�(RBG�fR��g��6��h+OB�2��Ěφ�Y��^׺�ǔ�L�di��4���L�$|Mnw*���D�F���E�"'�pգG���"��H��S7������c��E�`SA[́lzS<VE㊦|�T�SE��[U�R=�J��M���P��7�v�X����r�D�s�������X8_�`9�K��-���m����OR�^?�L�>�$�o����Ϧ�����9.�%�힓l{%�8l�:O\���wQ���m��(�sȑ��{������oт/��·��K�P����#^!�%O2��v$�6�[y����^N��CN�R�~�=���
�gCk�X;�zM�KB�C�R�}a�8��q�}E,���B�+G��_��x�O���J���߇/��y�ʬ�����	QǊ�T׮~��6-���&���)W���Q�b	���q�	��p��P]�{+ήnQA�N���dr�4UR����̭��&�WRIZQ
i#Y�r=��]at�U 瘞C���v��.���E��GQ (�G��0��.�es���^��t=��~��$�7AW�	������������hj��)��Op!�A�	����⳱�s�֗\N����1G�5�hL��m/��"\\�`6;�cjGIM9�)��NZS�Ã�r*���5
D�o��G��J.iLI2x#E���H=��Fi�"SG�rhg�'b!U��"{)�K��(�|K��<���*���Z'
}	%h��%T�+��J!�!��KK�Z�75)Ih��4]`F*$��>pl�M3���1� ��nA���ֽ�3�:��v�SCGCU�ۋ{Э.��7Mz:����ͧ���w#�7����U���,���q�yG��� �w/G��m�����^�=y�^�	�������.=�A$s�)u����~J���.�%�'�P�D��c||�7$�')Yk�7��ŉ��ҵ�U�+�x�HO\�(M��>Q�ܩ�m��B���Oԭ���j�]�Q_�_�V��b�}�ŋ�?.Nn��o���]� �W�.}y���Ot��?Em�CH�i��^<�nٔAK4̪6�[<F������;1e8�~鉻
s&{&�4#}�b�*��	lY�y��j�LT��Ob�at3��9穓`\CC�*��Nϑb�%�コM#[�ȝhus�	+ 2�;�̡���Հ¹9�*q+�������f�~>���jTZ ���{|��Me��T���^@��Xӭ>����������"�#���>��~���o�!^`���?/�"h��N��-h%�o���p�f����};��ia�p�!A7����T��,J,����8���������3��JiV�+��j(b���yR�xW���*<Ӫ$������ U�D���Vt��X�&8�(�K��	L�ہ��}4eT���� E�Aˋ��S��L�'�n
�q M>���}@8�%4�X��8�ė1Ц�������!K�8�����#�@�%#�p�b��CH�Z���[�D��Et������OǛ_���m��%8΄�������
m�F)���(���X��e;	Ք�Q�����y6Yش6HK�y��vu�2hv�Ϋ�(��?��|G��Սjv����Ko��zG��[`�<�Fǭa�c��s)J���*���"�@�5$�~#�nlq��C74���$ �+�*P=���\�K�i%lG�[P�-*���ch0�([P|���l�	�4b�Qz{�;<�2OM�mgeU]�v����L�����0Ns������
c�R49B�U7<XI�2�4��������x������/7����۟��7�^ox���hKU}p��\�5��?����C�.�A\O�ՙTlEP�S&�MD^�,���gU��L��q�#���u��|�Ŵ)ô=�	b�;%i��x(��z��'V�P����WE9M�R��9��Pc	J$�|�K0�ǊZ�ThTs�[�V*L�����S��'7`�EBm���p��[�(����CYm����(6w�P�����S�� �t���(=5?8Y��@�n�$�i�:P�O.I���@{�T����gI���+��^vE������t��~��3����|3/�^�u3���F*��0�fժ�JT_�<8���}y������Ev�HA-K��Ʃ��yE�j��!�4�5��B�d��%]���i �<��YJdr	����F�sx��-I�Q �E���j}F�ވ�2����.=��.��=N)���+���ŀ����ZS�d��P}�Cw��g��l��lx�?��Ռl�A�][�����csA��k0y���{.m���E�0L-�c�ln��uwq����@B��r�Z�7qt���i�c$��YH}U��H�MV�X��!b�M�"o��K-y۰E^�0�͆Ƥ����mN�|O�z�r�<{sHq�{N��z���<���th�]���b���J��Ē���s�˱u��EӺu�-o�O�{���4d%+�B�%�E��vgҤ�|ҿU�/V����-4qP�B"7e��!?���U��74է._�$?�fx=�5K�tcW�}HV�Yt�����8C߀��,����5�g�O #tB��'V�ul掹jLf��>���.E�>��t�M�&�������QH���ļe��r�6�
�Q[>D">��9#�flٍ�;�%�v�,j��1�GKl)8��-�9����dk��Q��l������([3�W������v=J���k���`���;*!)��)2��Z%�u�h䆢���] ��~��ۣ5CjyOk�%�p��ف����ʒCd̗����"�Ч�bٔ�.6Ų�l���k˾k��l�ȁ6d�H�&Uz��"�21�j���z��I��J�t���xYx���w��x�B�4��l���ob�?�d3�?�<4����s}����(��'ǹx��5yTe��R��s.�K(.聆9#�;[^�ǁ�5ȓӓM%͐X��yE���Ef�ܴ�<=����0Q2%:j��s�A��@�'T�-B�J~��N��ZU���J�ޢ^�Rg�70�ȑ/-g�8$�\�x�^W��ѲB�'jr�5(p�0�RoFT�bI���X�{����(�ltD�W�V�W͠���kMu�%-��#B_�E���]���g�ZVG��X�ְF�=���C�A�_�Vܧ��,}���9��H�u͊� .�S�t>��}]��NaDjޠ�49�Fu2���&��4�Iq6Y��ibq���ۖ�p��gV����s�$���-��2~�䉪>�ţ�����۟�q���o��^��~�����p���?�ͱo~.��/A���Nz�v���g0�1h�7+	��;������?u�g��>:���6�uu_7k}"6���|��C��,a/���F�Q��g�`���:	�����2Ֆ�G�u�J�2d%s8U2�q�R}z��Y��G6�uZº?��>�cΔ� @��)ǥHj����\Z�P���λ/�%�$E�=�Fu����b�V�*��`=����B�r/ǛJ"v�[�Ҭ:8�����{�Xb�s\?�h�[�鉧C�FAn�U���8�7��"eU5̩�.�nG�pX6<�7�5{�c���`R��G%1O33�A����{LЎm�E�~d������Lb�8����\B����v�g�i2�3�HF$}����1e_Ǎx���	I�<���k�y�(g8��8<"��<�y�1 �I܂v.��c"�w����KRmjua�d)����L�)�6�ԇ��ј��A�I�.����������V=��q-�R��zb�ʥ�jΉ�I���y{r���GŊ��΁C�(�ig>-y���]��;e��\�:�~p�fu�2�����i�DR���
�x�2�*y�E��bY�t�87��jr@�l��"��UPi`v5���x2�M�=~%*�ܶ�G��,�8��ʃ��u��CC(���?�w�N҇/�K8��'�����k�YB?��8{����L]��C�|'��L�"(8�&%jZ�6�Z�I	r��u��f��<�B�j�$�C��]w�|턩sm�������7����ط6�2�(�L�L.qd���:�*�P��d˛�v�GV�y'���=�2%������hL��!��(#�f)� �N�0E�6�,o�&`�{�W��G�����x�D�J]&l�d[ઔM<%��� ɉ}�*���� �h�������8�'NR�y�)o�	d� �h��o襱�0��)q�
���0��f�r��Ǆ\%�����vϓv�ں��oד�u�J�L�{g>�Jҕ#Q~�6��X����y �q�BB.`J�L�ڈ�:�u�ذZP3�R"!k��p��Ť�1�2�#��<~�bmr�&��8�e;�n�+�ΪL�ۆ�*d��*�kR�C�
�������Z�c�N�?)�9��>������	b�2M���i�6�߆L�����$I�a��A����;�CCV���%,p<o�AlDAExݒ��Ĺ�"���&��h���y�D��d�o��ɍQ�]ޯ-����0����Q�C��U&�.��Iw��-dW9I��_yi�e#��0Gq��������+��#��C��?Ã?7�y���$���6\����=�u��5t���~�+����nZ��y����!7]fi����u��!+����ֻ>l�),aG�ؙ`�<oBhT.$l]�8)IB��9�}� �������vr�L���g�8	���X�d�r����Nr��Җ�k|�vu�mZ˨J���lM���}��vT� �$&�tY`�.zV���UL�)1+@�!��Uכ�|�����|)$5��0h<�h��!������Ȥ�K̙ȹl��9�n���:��,��+A�0�2�HH��P�<�u��<)��nv2a��3ӕ�9�.�_}�x�т��)�۱F��.��Iց(�EI7�7Z��
u�KTA�6�UC�=��� �y��Y�cR���2�6��7�f��%�ާ���9.u$J؜@�
�h�$>>%0����ш�5mLĥ���L�ٚv�?��37�ƍ!���5��O��}�9{?)�z�$L1���B�A�Y�Y�4�1�5)U�;0���\o�
E��>�آDc¢��������̲mQY��@e�I�^>�y��QǮ���#������&H[�����<�V��g��D�b��0=W>Q�#~��C�����-";�Θz�UF�KF�!��ή���s�O�{p����~�f��{�����=88}^�x�:�(��w�C���ط5vm�xs��\�����Iv����4G1���mR����#׶j��aO?��8Q�h�{����p�b9���W���fVi0˗��Iɐ��%���Y�|�<N��PE�s�Rd_�T���-WH�����K�����P`��	���/ �4ٶK�H�E�{�QY�1�@Vq �HQj���+��� �|�t(m��k^֯_H�v�����
�yݣ$���:�wڵq��,IXr��ĻSq}o�jr�Ib�t�d�(<gh�6�@���*H'%,��%]c�O��qlǡ	ݬ��3��ᔼ��:���f�lW��9�M��ǆ{T:��+J$�}䡠d#$�yGLJ`�~��$v�:Eb*��(�q]s~G�]��2�{$�~]�d�n��/D�`y�doX&����׷eM���"0�$m2���a�l.�4~?���]	Ƶ�Q� ��Х�T<@��`
}��<����2��Η�}��#��u���z�U�=�K$���ƷCI��0����`���q��YwR�T	�J�I�@9�����DCi:�Lw���ԟ4Z�F���`��'�w���?��(�ā����4E�����<0F�9��e�)o �9��bhP��,����N�������S�-\�{�_�h^s�~��'䗪|��=��FR���9���K�XdWyT!i�y�u���}��'�իߝL�f������P���t�B�d�T�C~�]C~~!���S���ݎ���=�ɽ{��c�x�cB�7P�%;p��ě����k�E����s<�,����I��}�ǭ���6��|-�`�VJQU��r^B)K� ��qU�`u�I�ˋP�n�D�Z0z��0�:+�]?�}� ���]l��͠��������.��;AÀ��J�`�I�pE�>�"�{{�ٮ`�lН�����;�V��Im���y�7ޜ�i�ز�NpK�n��晓�se~eRR�@���&B�F)�� �p��F��T)����LHj����x��B��ۥ*�B8�^ݓ�D�³�A�`���{$�ް`'��f|�d�R�!�.�/�Jr*f8�G|CJ�)Q.T�F�0��q�ړ�7{�tM�ˣ���[G�*#9��ǁJjTdC#��$f�\�Z���n��%��>*	��wI#oܜ�Y� jؑ��*�EI�B�����~]!7�\m�K�-����oI��кR��G!wAE���ْ���e/�$Ĩ�y|�
�K���$1EP�sZ^�Ī.t���JGCP���Vu�����`
��+�,s0�m�\��s��c��3ߏ�NGd/N���P�)����,�_�����?�6��x��5E�ͽ�x��>׵���������Nd�Tj2��%id���T1J5~���
F�hIJ�����,[J��Z�8
L����M6�r"��%��k޲��T( 'k���#Yδ�6)]+�})*�x��+=_�Z��,x]l��IL#�r�_@�c��ڈ�����ńD@��d��b&��"lT�l5�R�/���c����T��O��d4��c�(��Y36x�{R�B=	�_1��!˞c���7�&�Q>=���f�ӸQ)$�"h�����ɅD�Q]�����Ċ!9���R��f�U�T�;���z�Y��;{��Ė�iĪ�R4�%_�xL�{=G�b4�F6��*�T�T���D�;ϱA�օPeO��X ��G�b��B٢`�)y����-TցK�&L��57[@���0�D��I>��N�Y����4��n;�q��_�,k[yT$�l����MB�1�_?M�5�a:m�&:�������R�d]!+���Fj�ˊwQ;;;��2ޣS]��^�ry�M����1��������m�u�� E���7
+u�(�h���9j�<+w,K��8?�B[�Oy�<s�^ks�5>yЕ8'cc�%������a/�:���<`	���l�S�����t��i��-����q.�7���u'��2�'_{���f�nD{�e�f��zy�7�n��}Sp�����c�w�z��MsY��MH��hxbL,��X�8fB�>'G�J�c�2�V�D��1̮��v��Ӟ�q��4u��B m���^k� �[r��SsM�E�D ��z�->�	-�ܩ|"���8�nJS���,��{N�+E�%�fn9I���P�`v���s����������I������4�Z)��M���}�������tTW/)7d��TaP-s�,sj��콒$"���(�%O�E�DN�&�����%Jee�x'�|ÄP'�G�U�{����X�%K����O���)����tUm% �͓����=�<_�$9����=�2@B)��0���m��n���B�����Q�M���$e�v��4��C��^�($a�/vyvY֮ t�lO���{�	�#�&I�N	����z��k�pDi����.�CMbp�+~����I!-�8�k;RH�H�TvF�c�a�4�|R~����@�����8�/��]�?kT.���v�H��������۬��S�zY��^��&����DS���|�܃�(&.x́���)��c���C�=7@��c�8�01�tE�Q^�g�r ��is�K�Gp��������b�����^��zp�f���o���� �͇n���l�Z�nȚr��e���(���M��Td빘X��\��DI;�6�ѻ#�sc��l>=�}����������Y��.+U�j��s�09�-�(d��(�rW<�a���@��VzB!Q��~�%5����s����V1(~�wgܣ��ϵ�!7�$���4�萳�U�N�����o0m];ř�`2�\�+{O	1G���H�G��a���$@Tb��J�8���bΨMb�Df� DRP��Vt-�?ML�R#�O��j!��-�o�����t��U1�٠36k��r�10�%�`����kdKx�8�(㼘(SI�N�:�dd��#�LÐO��f���Wa�?�4��#�QY�<�()	���ce�TE��5���d������\��!�I�l��%�I~�����X�۩I��\�@�_1Fr�!Q�>�����\S~y�����*[W'&�җ���6��#�w�����j.�a1�s��r����c���]=���Է�($�Y���mzQ�Ed<���`�J�G;��4giz,;�Ȍ�呻�}<���J���HBoAs�ݖ�)1��`�n��R�F�5�h��#�!\���ǎ�^���p�����ٷ�k�:���w��\܇/������Y�x�g(�F��ҌAk�q�s�{!�s���X� �$�]�*��t���D����^����f�I�qb�G��t�Ԯ$t���&��������[=�vۇ4�,`V�udbˍ]TI[В˽�ul�Ak��]-�k)�T�f-�,�I��� ��X�n6Ht�l�*ۻ��a��X�`��Ⓡ�'j)bN��C�R;kA� �5[#�5j�^�GU��yǥ)m��
Y�I��iY8[7<NG�^tb�S���%����(�@�f+%p5mtC�XQ��`�QJX6?�߶��D��57�LR!mϡ�0h9
S���jc!�dR`'
���S~g&�a!W�tb1S,���Cz��Ф�ˬfR[]�|��<����v�N�<!�M�I�6W���Uyͅ��!_��r�ZW��b���I=�)�Y��N�y��:c�rS�t�ɱsK�k�@��g״�W6^�A\�F�D�k$݊���Y��Q{גI�Y�q�%����!�z��BR��з=,GLt]��K<�j�\ӆ.��o6|�y�dx�뮥nN�qx����ֺ�~�I�*Iv<�����!��v^7OȘ�d�J�@T�9d���C�ׂ(�A�6�{Xv^l�g��&ޫ��w�ò�T�x�p�̛ᵀW����/����E�'o���?>��o�\��ɎBd�s�$�q7�(�7qU����Z����	 �I�:�^���0�|��ڼ�xcn�|�te-\�I��+�8�K��
"tr����ރ�8�~��2Liܖ5��!M��T5W��%���h���!�����QM*w�Ӥ;w+��3N����	mbB��]����l��h�Pn��G/~G���[-]c��>���bΖ��:\P�{����4P��>�$��Bզ�1���Y������e;�>�Y���\u'�Q)נ��8��+������ܘ$5U?mNZhŬ�Qh���Y�[����?m}l��f����x*A��!���D�Ĳ�8ւx�U��L�)�1k�@)��FY��j�
Mw3�I��3�j�y�-C5*�3�&��L����`� l��0,��d/���'�S��Q�7��}O����w�LTe��S�y�͎P�#b��K"qT47���T�V��.���	�ᙧ��'��{w���y�՚�?O{�d��B��:�i�z��3���Y���.���d|�qMoW�����7���'�P��jχIb��3��d�e��њt-��dI��/5�81�?Eq�.>�o��2~�����o�O=w��[x��w���W�Щ��ʃ�o��woo���o7({�}&�ȍĥ�V]�Qj����8��,�rm�X
�\����Jj=9d�i2�¨�e�|2�R��_�l��oyH��X�K`�m�N� mX+&s\�x=U�r�<%�����%�e�_���(��L�n�8���5��%�[6j�V�D�ԝE�QR&�1�M��#��"���P�7meK���v-��ɯ�ތ�}�ݖ�7����Ę,f&_3��������"'XQ�{ ��A�=c�-I�q�2@�޷�\I�Z�=
W*]�{��-
�
')�P�6��(�Fʯ�-
ZY1�����3Q~䦎��}�rL��5�ig�yQ�[bʅ�-��5����g/j���9�e��鐅ɒLXN�
<�Dh*��v=��(�$S����[���EU`Ұ��?l��y�Dɥ�1���b�rh�s���g����QT���є�`zOG%i*���J`r���[a�MY����P�fL�D����pr�&Z�K� 97�l��ԭ[h ��Z�=����3���{���.��p�\q%G�JYŜhG����RhF�6Y��ES���>[÷c͇��c�<
���d��=��M16��{�c*��c?���`��Q��Be�$5<l>s� y�Iߧ�L
�7D����������'O��^x-�U#tv�o������m_�5_��RO;�Q�f'�M��7�NpA��<���G��jN�R35�tڈ�Z��L[�����/�V-{\C����[�����ld���Z̠;D��s\"i�����O��UD"/�he�`1H�N���UQ�1�'�&�c�A2ԣ.�a����%Bt�lQ������aɄ^R�
7��x�k�AA���Q�(���ZT7����\qY���e�"@�ՓUGJB�V5�)&������1�3��I����T�D Q-�������J��VT��������ٔ %4od�W�jz��M��,xR��ͥ�~@W�O���x�m�C���%}'=�A�������*ق��mL�]�Ģ+����2��Z)��YK�y�=-��X�h�&��������F\�4	!XPG<�O�X�k��LjB��vO��(�<`�-�9�ӝ����)A�[����\FK��4����� '�qITUq"�Q`	�A��҂��ě�|mZfv�c5���1O����w�2�]fǯi�Q���笔�=�s�5���8V䵛�`�cՓ!T8�y������§>����wh�p��!\\&h.py)�>��q�KN�f�a��=��������~�%嫝3�D9c���O�	J3����M)��@!�v0�WY1���i����@%�*��}���j�76�O�Y�_^<��Η�=�x5�Z�;/�;������b���D���v��`z%���C��'��\���8Y�r��(�f3J�#��Qdd�2Y�-�h;NH�W��f"��=�	�+���6&�lZ4�q_!�N.p�Bk�B�po렞�$q�a����$�ʽ��I��uAP"_�;IR;���%4�x9l���P���v�@��%o�BǓ$2�(H�uM��cCj�e�m��kzKpduJ�a����L���&&�F��%J���-�M���v��ڴ�EU�L&tRU�8[���H������*o()Ǩ����#nI���\$8[Gh��̯�cu��i&�:��X�ZrBT�\��m�e�F�+3FF�ºB�cP�5E�@�Y<�kŕ�'��{v�Ǚ䮔��{����9�y9Ve�=D��7|��E/)Q8��+�y��l�'�QJ�����c���L}f�!L��S���2P'@�܃�ʥ��p-��(�SE 4AQ��wjmZ������$���������td�^�8��
��^�g��R�d�/8�������{د.���I|����x3�Z�4��,�ʻe�cA��HS���:똃���7k�����k�V�֘e�H楄3��Ys��cE�$�a?U��y6Ie����ݑykk#��p��S�Ǔ�\J�Ѐ���*�G��-��O�x�/��w���pt�Yx��zsvNN�~�� N��uH}#��P��h1r}�F���8�}�s`����Q_�w	�Ɠ�'�����p�[JȵưM#4!�b�[�����F�B�R�7� j����L��6)�2y��UKB���5��� �orC?�|-�5�)�v;�C��5[�}�HW5�4�-yG�4"9�5�lr6�kK��H_	a���&�D�a�5,����B�Z��m�v��1}�Ĺ6u<�en@$��ErCJ�m��jVHz.]��I��8��cŊj�_:kᅳ _zZ���E�q�z�t�/�UO��7����2w= 0n���jb\���|DZh��-JAR��֪d��G�G��[�!}"�.���$;���95H�L$|���������k!��S偽7Ɖ�l�p��8�2 g�ш��5��nZ����$�ܒ���~����nP�=7˱n��a>/y�ɻq�8�c��ɫ� ɯ�+���a�����{�����P�A��ީ�%XR�=��R(1fz"�
]I��Gͫ��Z��>okc+7��q]O����ŭs�[�%�Pb������W0S�Q�x���~�o����'�O��77˗�o�1� �^B盱�B�9{��.�o�7c'�9��i)����Jyw���V�FBFw�#0�~�q��ݷ^)B��M�T�Oj�(��7���T �h����Y �WJ��h}�E�Y9���
s�r�`��	��� 	.I�<m�B�z��*�|��`6�Z�Գ�w>��ۈuS��{A�|�E�F7t�^uɤ�4�
&�^]-f$����ȵ'q�f�(j�M���7!��J�B���Υ�!R5�^E'�Uڝ��������iܼ��2�^z�����}�n�"'lKD�g����2���``ۮ�G����5�$����1L��
6�7���8�M����/�t��9���lߛ��R�V�J�R�/����"����(��܈֧ݮ!f��zy��B��غ��eO\�$�Uz>�M����څI�O=OI��^&�����[��N��� JIp�g=���f�
NN��`�d^�ť�w@��е�T�6dE�&��b��_��h`�l��ym��� smnM����d�sK��9�۝���������5����W@KC9	���310���"c̰�r�Ʀ%�E���J}�U�Uku�S�|��?���~�s�j�N���]��>K5̧(x�߬�<�:[���9��d�jKCޓ{�^����7QmL,�.Fbe�MҰ�x�+o`��R��8=�� ?�g�w�W VhT�膤wS�5�$K&I�iސ���9W��.b����ӽZb�e�b˴�e�#Gv'M��K�:ơ��s)��삋��Ye���Y��uÊ��p�tL��J��y���Dr��ܥ��d-��Z�K�;�d��F��j������0�OJ]8E3Yon��q׾P�yW��(\�o��O$fg
�e�@�m��v��~5��h�
�]�`�����&!A����JMi�Z,tS��Q�n[2_C�X��e�=|��4��1����⍽z6L����#Xמɸ�\����Ҵ�_S(&��C>.�<�sV� _��� �W�=�&vlK㧍@�gcYƿ�9���1�
��LZ[k$�7�+�-o
!=��㰘��Y<�ٽ�R�f15�w�`��o>�a�Y絜� ��\P�6<B>JF~�y���^Qv��;߷�I����5z*���VVԜ�2��B,�>I�d�=��Fϱ(�]�C��R?����ֿ���\��=_�M\����߮��ˢ]/x蚿�7���mX���ZXw?b�,��d�=\nA.@�`$B$׹�G�\ՌU�]gAoY1��)��?�zVi`���e����R7��w!���F�t,g�X� �	iyS9�� �z�`�B�]�TW�}�E�������Jv"���8�t���s�%�4He|��D��yC�$�,�Y�W@ز�L��b3����
d��`�2oՆ#�/fg�{�Ƌ��8�4�D����,�l�XJb��Ś�X�i k�K�vڃ��3xжp�V��&�WD���5V�5�xW��Cf���ˎ�%@�H,�ŻA���Nj5�2�˅D-K�d:Sd�e��}[����{�P��M�A�zK�"[^V�8Q�lL���9���Zq��;M��Q1�މ1�vW}�q�5u�5�M�� ��=����=9fP�6D����w�w�	���)�Ԝ�m������'�C��%~��jV��Bߺ����{3,�h �ӎm�Iߴ�����D�Ъ�]��E�:O��t,�*�Y1�fM<��d��f/%+!��^J�r"��� &���5�ZE~S�]��șh.w�o$;���M�cE9�����W��V���?;|A	����7��+a6?��]��Y>N��ҾɺI'[�)�֨bK�BIE� 6���Y�[Hٕ9�Y�	Q�R��mvZA�א����i�^���n�3)с�C����DpqM�$i�媺��ؔ��dRW�-��I�u)[��ЙЭ_�N��]R��.uqXs�$MBt���*ĬJC�w���7�'�\�㉘b ������A�D�f1+� ���Ж���bҽ�)9���&���b�Iw��)f��'*g	��W�]�pѯڄ�v�Ǽ
땐���lܵ��<rz>z�N��e��Io��22�;z�;��=��u3
g���[�׺J�����>�"(9!e.5��q���Q�*��[�f������k���My׫�Z�6'caT&s:�T����7(��|�jS�y2�('.xs[v�g/����
��bG'��#i�~�ʣtB�F<5�[3�..a���=��S\gN��ٽy'�'N��=�,8==�^�FZA���p��1�+��	����d{�\�&��^����Vr�����+%6M����ż�ܹQ����s��8��,T�q�GjPV%{�����>�۱��Aw���܊Ο=�`��>?�A��^��'C�~>D�s1u��7,�j�LV	b�V$�/)j@�.A�����`$�m-������B���y����W������B��ꦁ||�V��GGv��Y��Fi�ܩ�O��2�M��g�'�&)����ִ�]�T�ɼ��7m�J�mM�`�voE)t���D�����nd��5O}M�U��h'�<g�j"|�u��FO��_���Kq�L����ͪ���~"̙��$�
*y����8&��"��Q2� ٤fVע0tH�\Y �O5H�ڑ���6��yr�u�ǧ�E�T��0q7�5��O:)eK]U��9>��޾�z�$.֬�ۢ��k���5��%��!RzO%瘃�:W��k�֯��A�%:$�G�'�v��C��{-+U�,���q�U���my�;��߯S��ؓ�ܾ�w�J�A� "_��>�
�ɯ�s��K �1i�
��25�s�|�V���N�H/���baW|�e�{�̏P� ��/pXpY��l��U\��� �����Pq�Uڿ��R�k���ԃ�L�������mu����2�?���J[1�Za�'��Jr8�\$�p�y���H+�,TN�ᨖy*R�\�;\Փ t�,H3�����ۼ�o�-g?�V��yo~z
_(|A�k��(@������6�ݱojj#)�C�G���	���ٹC\��9�eM%�����ė�T��4�['%��Xr����c���[��M�W�9d�`�����抓�"�Zgk4e��(`P� L�)�ߣ�1��&����d�S��
� Tiꓩ�6�����k��6*�};.$�.¤5�J6��R��JB��5*=�6��v�|�Il�ܠ���}��yF�\$�g��u�㺃YAЈ�*�</Q;k=
�V��ӆ+������Q2��h�T����-슊
)�Qq9�f���D��Z
|��엲���x�"ߚ�6S��+��0��ʓ����
��Ne/}��,Gj�K%e�Pi+YY���d��[�k/��O�[�&�?��i�YҤx���AjV@���E�	�����Ī��xt�,�q��m��.�O���#v~�]��\������"ϋo� ���k=iR�y���pl�ĭ^c!q񪬳\x��Gp��-�=u�\5��ڼ\�f.}+��G��ʧ�D2�����qP'�ڔMf���Q�޿�������k�h,#��lyu����'
jV�B���f�Dm�
�*�*5x��۝;�C<HR���x���>�+*y�0/M�p+�Q&L�~���z�7�����������i�����З�_�yw���OR��t��J����	]���i�&s���?�Ŏ]����.�	�o�g4Ɍ�����N"u���ͳ�29N>^'�Ð�n�ט�	{�)�SD��,K.���hЉ�GڧE������\��r�*y�t��C�lx����zr���U��_����bw��������ըoG���j҇5�:
L�fJ�uϊ�.֔욖x�w�;+��%g�����$q�8.�`����� �^�����>�H�?u��`���h�L.�d�G�,9�}�~[� �[�+��|)�Ňg8.sn�kQ�	����c�,?�L0W�Z�Q��H�5�G���S���G�C�Tyz�enϧ�u_��re.��}-Wb�3� 6B��c��#���� ���|~]����͛�m�۩.Jj庀�>��x�e�g��g�>����Ƃ�"Q�Z��y�PE����5m�u߄�2��M��'�}u<��e�ݞ7�Q׍�f('�'a���޺?I� ��e�
�;%ҽ�R�ް�j0�@U�+jo�BwL�
k�-�&��6�\�[,� U��{�;��o�/߇/>yp6�w����S}���خރ��[�Z�݈Ƹ9g>�eHY�-�=�7�)]�l�&�.!�4ɴ�^d[�G�u!��Ab�����Ʉy���nPS��/��c-9͍����^��kRO-�:��7ߦ�,�YE-�Ӗ�X�%u��������v�c;�)1�'n^!�ȅd��wǥB�\&l���Ucۥ+c&��B�t[���fz�-�v�ޟ1S<�X��M�t�EA�čt8Ӏ,sj&�.*�!��G{r%%���RuA-�QXPc���A?���N@���޷e�?I'�2.�>+Y��w�I=deI�ħd��)E{��Wf=p�y�����1Z���s�Q����i��@7M2덟S�ݒ�)�����~���Rj)AQs�NC�Ӷux}B�u��+�r�q��W��%� 3�ާ��{1Q�g�1�l6���S8����//6��@�s"*�(��n@�@����-$����N��E���1�y���5u>��:ٟ�6	�U����z��l��0�E>�=6~!+}��NtJ�ZJ&�V4�}ˊߞ��S�>M��i�3i�6�(�v:�0�9J����l�I	�)Q,�PH;eRBe��5�3�;�凊�����c�m._�����������4H���tެ����.�J��,b+{�Ԣm1i;2iB[��5��|��F�m?X�%�+Y��D���C��n�V��qn�kH�:�ݴg��191X&1�d
ŤDm��0j��ʠ�\��;$�%���)�Ei=��-��ص�m-So� �~�~�o9k�Hb� j
���]`B�=7[�V�&�3�a�����K|�V�uu�E&W������S����cS�<�<M�A��x�s"ur�i�R�PgŪ{К�pQ���-���a�1e5sC-Q�K� ���G���X��u�3>�p�I*�Fg2=F(]���Bھ��q��9�X?�q��ǿ(�2�ę3�r���&��6��p��v^��a!����g�'W��z��y�by]��nb�+��QK�aHJX�6�)��Vб�(�3T(G5�Pt�>*_�f�!%<v���|
���H%n�wy��3��U04�,����@�P]�}��r*T��v�����{f.E9�+s�����'d�h�)~i*���!�,�Y����c�E1GB�>�A1���o�I�5v�g�G<J�;��εC�a�7e��+����'��v����z��z�\�3?�볗�v�ڿ�oV7c��d�iQ,\݀%��>���F�����Z�$<��c�nJ���Y %\�qڍ���B)�1�ʎQ�u��j���D��:(�O��>*x�#%�¦s�꒝�QM�n`�.�I�Y�gy^��(=�Ţ�ms+�$�`�#W�}ZpB�ԄG%�"9�Js�b�m�9�{ ݞvz�����l�̇[@��:�J'��}�>l_f���y0]�����g�#�j�������}�%NJm39���#�;]].�J��
Y&d�RNӒ�"�>���:�"]���u��ļ4ꉹ����&�8�����G������,`Io����QP[�#�r�r�X�R�'���%�T��)����v��Q�񑐷�aK1���n���&�]"�
��הG҈������V�����T*q���^�Q��I��QJ�+��XN���]]Wp���a����K�Z���vg�
�K�G�5`��1oDĝ���!�~���Z9I��W�"�v݅���V�{-f�|bi�c���� �����x!}�֕ +p�x���mu.�B�&[�Vѡ�
"��̶(
5Ri����V�?���_���~�fu��x��������i87�α��h���з_ie�����s��\wXz�Ķ-W�J��Q�y����}_C�y���Z��H�8Y�6�f&���˙���da�
��s���2��S�`\�I�=��$I(��B밂U���A����3�jId��6R��>hֶ�֔`{��-� �h%��Q��'� G�"\7��)5��M:�!>J L?ÉA�|n�h�.4S�̃!���p��JmH�dT�8�90� �E�V#��ą�(���yAU�7:��I�[ɂ7 ��r�Q+>��Xm�!!��,�_�� ���[�}�C~�k�:K�s�5���CĞ
Ʉ�.M��H���Z�Ie$�[P���;,��T �"�6�&��(k�Qޝ1������:���*���6},�I��c
��\s�#n�[�V����8<>��%	�����/kr��PłyX!��ap����T� �d��|t졛�+VVc'�[�S�MFXZ���m�n�n�C&W�ǳ=/,*����#q��{���D��2U� �*�p�o����HZ��N'y:�U��$�����bQ侢����q㙏w�;/�N�y�g���B��l�8�<j���f�]�݄����n��m[zP�}��2�\����s�JY!�,�HDDL�5�
�1JIb�D_�<��� �)�A0��/�!���*����9���֚�K���k����?�Z{�S�����s����/�����F��V��t��ˋ"�A#�"���鑹,��`�̈́�[���5��������B��x�_�z�Ν���|�	�l��([�"��mܒ�5g&��1�f�S&a����_RQ�<�����l5O��؟;�vW~߇�٣�n�;�)�+� F��^`��T�h�=��Z�&Ώ_M��^�����_Rз8t�G҆*�mc$����&4/����^�eD@�h����.jW����%�	�� �ѺJ"Zsƹ�o��]�4�De��V:݀�-�?Gk�"T����6y͗�`���Gl([���\��*�B����=�����~���:~�P�=��FӨ���V�W�B���ԁCa$e%�aj'XU	��U14D1���7�o�p/���#�%l��Go^��ڝ���F�H��Q���t�TP�O�F��/�"���t���h���F#�J�� ���Wo�p�Z�23ʴ�O���s_U��P,l�$Z=��}�WD�u-���Gn�Mw2��yvs>�mn�"�}���_�_=d7�]�WFțu����ϑ?�^5�d��0_�ޡ�es��)j�3ݨ�>(��K#ǳd�D�3`m>��)$�HT�V��ΒH�-��^�"��~|������������*�]�o�B������]�@�?|�����_���ﱰ4W�� jq׼(N�E�Y���̳*`���*��m1��*:T�
dw��gIQ@����ș�ur��.�"�TK�L�g�^+Y���S�Yy�r��	�!73P��q�o�[�MY�,��N�^�*�8�ŭ�v,@X�c��>�5QAU#�U���Z��ރ���š	j�Q��
�&�tcg�:Z?8j?ۚ�O���M\P���M(4�� )>X�:R�*�ܽ�F_�����c�vV�MiOh���J�v2��q̨���#�246��L&P�����6�$B��a�9�vC��4,e����=[Ӯ�B������|��{on �J����\�2�^�h:�C���Y�綞'+"�����b=9� S�^m!8�,=��� ��ת}Đ5_1�V���L����v���LD��se����^Id��^8�Љ�\��ֺ�y�M�����tu*T�iȑ뱚�x{~�PFQ������Ⱦr�e���ʔy�/
����u��{a�D�ߊ�����f����ve�޾���\<�(G �޾�<�b8==�W/��U�z�F�W���x�z�5-���ES��!��m��|,Z�{�ϛ�����&��!J]e�+y�׈�hx�]��8w��c���
%�\�c��5��]Y���P�����iz5��O_�~�W�?����{���o��SW�K�������/��ߙ/����R���3�7�ޔ 9Zz��zG�ඉ}���?��-�[�p�G�Q�w�& Q��<Y��Xt`F7��z���b (�ZS�@3��j�m�>�/4����ۧ����ůy���A��O���=R��ٵ: ������(.2h[tC���{�gI��X����R�#O���v���?:�.�7:�:��G6zv���E����X��5mg�k�>SV8f��E�=h`x�y�2�	t����vʙldΓd?�#"���z?^�6�Q�эk?&��@�E���Mݷ���;0��~�*�J�%��T���'%
�R�m䳃��d��1M�y:t����~�Zm����O.ج���ѱ�3n�B��k���	UrC}���=J�1�}[E�-���{I�Î�	E���E�V���uAWCx�b��(�o�J���ûw����������׋vYC�1z:�z������|��ƛ���z�����M��n��V����qQ��
;��#X��6��:I�y��B�-K�o1���嫿�k�����߿���@8�SU��E�b��:������r}�̝[��܅�k�}1���ҼUe�F��& �WK��׷�z�2�|�/�����;�ë�)��ټR��x���k��My�R�!6����#ú)Ѫ
~�ho�G�A(�zz�t���$��˸�!� ��Hκ�RC�4ԑ��}Ԯ^��T^�jJ��Ew�w��+(K��kZ��L��*��պ��7�$����@���?l���[��\�^�� �Δ��Z��j�g��^"6}� %��QI��45��}?0���:�1��-�y��d����q�۵�\	���Oϕ��zG��j���uI���^ڌ��Τ���e���A��OƓ�C���Y]u�S;oto*��B��ί1XJg�d���ߎ�����Ɔ�����i�G�KΝ<�11����=r����X3x��:}�x6���u���o�%����(E��(��PN{���=P3{ʾ��Fˣ����ʚF��3ӵx��� ����_��*E�5��,��g��=�*���֢%_�O�����q'��uq���ֶ�A�Q��[�I#�̅F�*̋7p6���	F�$�D&�5���0��y���X���oǽ��:e���)���տ�L�j�>�3؞�����|���eQ�y2��W�����j�ӲP� Ǣ�K�	ia �RʂF��p|�J��3��<�R��Y?_d�슥��D�e�a�bļ��{jA�\7w0���k����s� &�Q��~-�I�C/j�x�E�>�P61�i(q�ﾐ�fDn�^B���E=Kg8�|%�v,�j���^z4�'U {�+����^��N���r?v�|��~�c���"��"�n��]{�k`��!wc/ÞܱEj��[�������g�/�t_�6a'Y1�1����ӱr%ͼ|����qS�^(f/c��hG��U��y�ݼ��a�n��h7��^��n�
��
�j�f�k0"+g�5���xM�%R����y�0��>����_��b�X���k�n��m���x�9�˽��qel�M���wX5Nξ��zd1��q@eBGE�j�B�\ �
��G��OS��4�e-fI�ā������2���y^}V���<͗`,�Z�ʆC��՚^}�u�v�.ݙ�]4��V�	���Q��6��'��%�%�������Dr0�-���4R�`�"���i�?��|��v�ǿ:��/M�~ ��?�S�����~��o�ݛo��e�������4=�}{��������
|[<0�B/
	 ��V�3������;�t�,�l�╏P臷���J�{�M&0���T�%��f���z��az��ɽn�����k-�^��I��[m�m)�ħ{J���f*J��(�L+zW��(�=x����Rf�UE���Q�'Q5 ���Q�6dw��
��>�x�;�A+�cإ���i��S~3�)�~/�#�������/��]���~���gi�`�z��+:5�)���Nb)~�F��cW� j��L��W�Z�0/s*F�j�0Pj�g�yP��y�A�j��`Е���,=�hu���nê��"�� �vh��>B�6{ġ�S�3�Ҷ��e#�:e�yVj���{�V�+�^���7A�o q��v	~B��7���=��Y��s�[���o5r��������xi߱ȴ"�v�����	��ݴ�`0�e�"'�p'<z��PB��2���^�O4���^��q�R�2���Mꮽz?Rׁx�[|�0Ѯ��~o��Z��Z�k_�� F���ϕ���VV
�WC�H�ޟ��Y��,w�X���\�����g����*O����$���)�߲B�^I�w����[����z�3����M�'�Xh/j��f����K8�}1��̛��
��-���H,�76Ў�$j�w�P{�H(�I&� >A��La�ڊ NrJWq"�`�#��/lG��!�������Cs���@�4�@M��|����=��y-�i�g"V�adi8�!4�he����r�����ʹ��Q��=�VkQ�4tƇ�ܳ�uɳ[�7��B�aý�x���Xv�~��[�@���g���ES����]�Mi{��+J' ��\C;�"?�Ctk*�=v�K��f5C~���Q���� |ٓ���5̹a7�Pn@v5�Xg���nAp���:�BGs�?�?�7�ɦ���9�sW��Z6�@:�ixI�ui�yr
Xc�����f87�҇��{x)�ѯ���|��k�z�O�Vv��9[�IG�t1DNU��6�M�GMљѢz(2�un��
�<��1�9�n�F��D%4�gww�{x[��I�����E uw,��`�P��\���R#>Fm,_Zu.rۿ�&�.�w�g~{T��H�&�� _t�m�~��"�%s���v,��]xv�b�5���Z���1�xw�����O����q! �G�|??7]/��\O�X���S`]K�g�kW�jW0�Ek�/��nu���H���T��$��g�B5����T�Ҹ3��Q�	�T���������<�Ӣ��y~g�3ⓖ��v>[*���z2��������NĚ�d��$:AMyy�>����R���R<yx�0��ё�Ex�(o�����X�v(w��G�n���RPϳ���Pc3�|�I\Y�:��g�/��7��nKy��%X��^������s�G6��yR�O�d�˂9t
_�9l�:hy������G{���<�*Dd��Wu��B��(�#�����1#/��KJ��G���*�j@p�Gq=�߶���#�#`��5�[����a����s���oU�Zֆ'W�5����
��@@%�=��iP��h���j���c���/4��X�j�����`�o7"��]�d#01�یZ_OU��� W�E�2�a���rc�^�v߮��#Ǒ���Ԩ]�GN��=����C��g���쳢�Sq¦yV�6@��"��tY�S�-�E�i�(ݛuy��y�u�Y�i�.ku�;��~zA��I-��m�]N5VMRq�6�5+;L�$�x�&�^�s߃Y�����'q\�w��������X�~���:b�����y�\�����?��O������I����r:���;����#C����^��MTDs�)�	�dJ3��-d8x��=��j�pn�gXwP�×�f6Ҳ-�lԖ���#��T@�D�d�T�gm"ϜJ�'��`�	�fq�`�nf�*���)ن�Z���� e*�)�{eIT`h}KWB7���F*��~���BN���I%E�3D���d�|����x]��ˇ��	H������Ť%q���<?E�7a�	��|k������)Ȗ>YjL8w4��l�o`��톻=|�ݩ�`4��|��m5���E��"����Ma^�߆��/4��;��e��t�Eq�ky|(c��F9[s�`����]5>_>��z�^o�|0!��V#�ټ�Z�`LF�\���EԨSwpz4WN����)�1_>���hl�s���ma�c�{�{d� *n���Y8��M1��"�d�31(����JȪ�*��.���OU���;Ԩ@Ȟ&0C�*1�qI�A�
	�X���F&���솲�_�4"G��Vͨ�=���@)�� _PE�.w���Z`��*��R<GI��eY^e��N��mr�|�^I>��V��:O]e������`_�����(6��~N�?��iT܉�0�
��� h�<��z�� QE&�=�!4�����f��ʎ�q�ȏ7�b��s���c<���K��-ʗ���)|{v*<������/?���u>������
}z���;����g�z��G���o\Ϗo��(�f�o�n_k�9�hiUT6=��u���
�M��Wa?�Cnop�Ml�:H]h�V9L�ʏ����?d�S��u��z����_/f�����)s��7��s�}�5LIDds���z󰗻�^r*�bi�y'sQ;����bя� ��:��z)C?�����ߒ���2�{��N�~$�r��nA��z%�����`JX|C�}��C��2�O���>&N���ۼ��|;ߟ>��
P������15t{��RE�&,��8"�l; �]����A��J��& ���=�Z��Z��i�Li�̅�_�?u?�z���ކ�o���Wf��n�m���TC�7�^�lS�Z�f�3Y�,��x�����$���uj���4�^/�k�j��ag�[�}��-�S���%r[bթ�hN�hk>�����f��;^A�������ϋGC�`pg$�	�H��?ʬ���P�����,?S��Md��{�Ҍ���2X��>���]�~�x޻E%t����>��e�fP����nJ�fpVo�0�Cu�܈P%O�!V:�i�#,��e�L�^�-��r�4���\�J���Ff���^.���5�a�%8���5�c)�U���$��_����Z�5�x1"��?�B�ݡ�҃���?���;����r� �j�-$kɎ\�ε,�D3��ܳ���nl�G~�؀3n�s(�k�z�5�����TA���~'�~_��P�����pS̛UG����������<�I`����ьr���-
���܅;PHI�g2����/�,S���{Z~$OO�,ro������^����=�q�N��p���b	k�k�8��7�v�K�*�AC~�4k��7k�!���y��>�����><�~�.��?d��z����ƶ�])�qP�3��M����Q�e0J�P ��΢��40��B�^��؟�[�}��
�l[�7j�'�b3g�!�[�L�<�Q����sg^����W-��Fz2�ޑ5���t�Y%S�p��Y�_7&��6����S7c���Zq%�G�|��1���H��ӏZ����^q��P�5�^�s������
!��x|(:�c����6�"J���W��g�q���g�(F�8��*熕k�
7�mܶw/�6�V�����T��!�������Hw,���
��(�=�[�*�\��4�F1Dfᑣ�eV��:?	*���, F(Y*����=���m6�=�q]��7�s�+{���F�����������G�����_����)�����Nq9?�����/ͧw��KٜW�6S�vX�Y4������>�j1�:Յ���E����6��=��� Z�����ꅺ��+h*��}��·�|��m�^ͯ�3a��Ԭ��1��6
�C�Xl���CQ��������l�}��+
�5=x��\e�'�J 2������[?/_����Y�Կ
�i<�c��S�X�.wd�4:)�0ރn�$�_��M�JáG���`	U��Xނ�^�O��S�Q��>Hj��X�K�ȣ�N]���y~92u��2L4wYv X����xO��ˇ��-�ZL��mpٓU����|�$��.���YM�er;�������]�|��#kh�b4V.��0���Մv�HYt$;�C�0�R"���HY�R�Q2��o���j�U�����ߩg��ٔ��P�^���{��cp����������K������ah�`�'�����Q��=Gy�;$�eg{���9��k�*��2CM���LK����(鬕;���U���m��aE�`.<�a%�����y�-oU����wP��+%�}i���9�7�w"���R'X��*�H�~�>�ax*â\��s�5��<rR�l�)֋���*����=%d�_�9W���(u��)ʟ\b��������w��<=�H��>������|щ<�-�g�\��t~���ǯ�Z�;ԙG(oҼNT��$��y���@��h�Xzu�&��d�.���`qԉwf��
�#ʮ����X�Y�fx��͡},gۉ�vM�b��ڭ��N��=���P�*�VEUlQU�vo�8��v��+�Rm#	l���������}W޾�L��b�;��>�I{G>V|*w��vh�`���R꽭/�=5T�B��z�~
�U�] �����龻v�����dyҒ+��C�Fs��:ۅE�wr�������E��'�;$,YS�g,�R��j���|�|������V5�7��C�*�|M�#Z*�yD��Հ�T�h��: #jpr�s�AHF�*�g�v<gO�ʛ��(�\��p%V.���#'�	��l��>k�q{�.��t<�9�܍C�>o����о({�ES�~���VC�5�Η�pxQ��f �^�7<Lf=Ǯ��p�� ����1����%ˈ�'��G�����zQ��R����ƽېf�9�_�7�S�l���`�AI�X�m�0KG뫆�6�BE։�@C��x�a���gȸ�V��HAʈzP�VR ��4F��K�� ��V�l���;��7�7=�wG@�4�A�p;�FS�
^oE�;{�a�p�2�)#�o����o��O���	w��Ǐ�����&-���r�����_�>�V�� �?+9�D�����Dn���P�ތ�J�<���}���B Q�1z�C�/�v���LD���D]FCZz82y��L�%k���Ѽ��� �k��A�u��9�F�l�+�2?r0[,g����Q�~�/9\�P4j���g����O�$���坻�����x�����>�s��r?����!f��A7��;=f��թ�r����7o���<�	�m��	�7E���j!���N�UE�^0�=�]�0ʎ�xWzp Ѷ�ݩf�+Bc�.mL1Ez�#̡յ�xnU�o�Tz�ln�^��z����.u��v��Ô�y*�w3�=��5u#�͇�0��a�����	r��X�EP�7��4�S9�U;�dݧ,�,��n�WȵwOE�T�\2Дzĝ� w��_B���+bvy�/מ�����i_�V3���9�lQ�\�/n4@bM�Ziٮ(���ӎ���l錸�ދT����C���~�B^�AK�H�؁�x��P������^���A�]O͢�9T�0We��h�H&�<�8�X޳ WCJ��u�_���P�@|_�eO<�G��X�Gp��j�]�G:�����`�y�������ȝ����.���9m��8�}nʹ����z�f*/��#e#�rT�	;��_ᡫ�D�M��~���B8��?��5���p�V~��)�ӻwEYܕ�9a�~�x�n>��篧ޯ��妴-��֯�Sd
�kiU.w�PK	�]�}�]>-�p��<DW�����db�&�ڒlK�hf���D7�O��?ف<ǟ{a�B�.�*,�1��|�<�gR<��X�Dw��jݦ�=��r�E�#<�{���@A���x�&:��C��x�k���*7���{E�iX��Q��r���G������o�#�h���hlT�-U��{� �(z�\eq�H���k>f��?��j��"���c2(N�/g�3�!0�נ[���Ƶ�&wE���p����r��������{ �s^�<g0�0�*;<�1Ve&R+7N�KG��{v��`�Y�֥�^e~����������U��e��W�a���$��^Z-�9b�A���Ú��geAiL�����4Sb6�we�3���_k�;���-�$����]�:�òq�ۯ��$���o=��R�7n<6�C�>v�-O��i�{ Os80����{��Ľ����@�j`��dW���[��As��_?��.���H�w�a�^&�,*Ӯw\ټJǭ君���)w��w�am4bi^jmuٺR�g B�)�"�"���T�����i�/:	e|�����gU=aE���}n�Ý�C�Y�tb�<��JW+m�]n�՛��c�������NW�@�fݪ�oķPw�m�9���YC��Ɯ���ǿY�\R�U���M��U�yz�R!�����ݟ-��_ZO?z��w��IO��fKN�=g״�rP�"���:�ⱆ�����Oͳ��F5�-�����&ر i"�K,���w(�Sq�)p@�;/�G>yY�������Z$uY�b��R�ŰZ��޳�n#X����+��:e�/��-���� ��+�,�c�w�5� ������;I�b�.Y���o�)�2V@ǿ>|F �~X���/ ������읟�����E�5M�	(-xS(dHKk2	X���ee)HP��i��])\���e�]O��VHF	�\P<g����Y]i���n���;֍=�t
Z�X�������#�	���W>E�G�W���2GE��/�\�2v��/㶔�>�c�OlMH�J�-Azu�l�1�F����k�^��pC��4T�J�[.��c[�c�ߣ�j�@���(�в<�j6��!W�&�����|�����W��zY�F�ʚ�F/(u��G%A}��%��ٲ��T��X�W�n3fl�A��V~]��|��\�@{�ym���|��:�v�U�r@�#��6�
v��16 ��<0������y��)G�o^_g|M8���{��@�T����^�N�^�Q2��j7ID4g���I�5�e�6�>I.���0%a�:�M�Ր���~��� �	Q�M<��!x� ���h��u��Ɖ0���i�(�U��p�J�|(J�]��ׁ�]�L]6�Dyٵ�����~��]����`z�S\�=1""�bK��QvEE��%��x�����ͯ�ӣ\���oV�6~U��y�����|�{���ry�3���'�R//`S���^�{vK����ۉ�{ܿo�Ym��|r��������jZ����P&XЁ�D��}C�Z���NoF$ӟ�<��Iw
��T��c��^�]�+s���p�Y�~����s|�#k�A0��I.E8^�<w0�t(J�(��0f��JA���;�k�KV����Px ��(��;ʮ���Kf�����|b��N�/j���roZa^�-�"5���^�OE�(X����dG:K'�(��pZ����֮��Ɯ&��|�B�y_ky�%�s�j��5����H�I�}(61\\���f��24l�7��ml�T0�_��-���kϏ�U<{O���e(�����]_B�����uL
����|�`�+���t�j���G2��	 �aQ� �0�M�#��%��������k�F3��/�H�zu���^��"��ЯG���G����J��(wϻQn�ѽ�u�������)�8����׮u�5��Th,|�M���1�t���`�Q�A��}���!��8���@�3��G���U#�u��
9U�ƣC)/u洚A� e�����@6;(sz�@�f���Q�2	�@RW�h༃�;�sU�����Λr8�Jl��/�?|G�&��J��n�����t�Gv�a�l,}9�3�Ǘ�vr���_�������7���w�vΉ4x���Q�$��տ"ǻ����r�!����|_~�w��w.~����ß��>|��H!�S����	�k�CPC�#7�e5A�7�k�xc�Nw�=��Y�l�ia}Iئvj������
EA{�@]<��K��Of��~���7 �&W�F�ҶP*6��9�����@��(�����;��ϏT�;@��%ɑ)t�Y�XD=����xG3�3�b/J=�1@ɸ��(�VTeƼ(<*�1� c[��B[�d\�
�t|Ey��cic��@�b,(*�8�T�V�<u��aC��������_�9���>m���B��(%�2(�����#�zܰ��Oh�{�k��cUVַhƗP�[��i�/��}����6�'%sx�QwH��[�u����)����Yk����W��ο�_-�bD�ƙ�%�g�_����&D�D�*��9�S��g�0�������K����_���E�0ʳ�~��fS��*W���u-�Bv�o��90!�y�V�}�����'�TY𖵁e@9	0HW#z��ޒ�#Q��ma���f^�T:Aw����Av��F9 'Hڲu@�JC�Q��L�x��]��'���e��7 ���\�SJj5��jm� Wp��,�Ψ���#��b�5
#��li� ���Q��'��7�]���d��e�$��r��xqGE���t��G����FU�Jy���LGd��pE|���~��?���ez�O����cw~�������3ǻ?F�������o,O��}�ˤ?	�������������K�:��ѿ6_>��r�����,��2��B�����(��#C�z�B����.d]�>_��Fl�΅�Y{o�;(�����`ĬV��֖�6��j�Y�͆ͧr��V_7��jt��w>z�t�|�m���P`�V����0T�r�e<�1���/x�j��ɱh���:'-J��<� ژef�|����>�G���ͥ��Aٟ��6Z��A��$�X7�_S�p�V���"S4���깣.tz����<&�����N�p`e�)��z[�|���{p6���<�����Buؙ2���T�����QO>�,h���&"��'2���	ePF5����gZ	Q 8�y�T�=���k	�	����h��B����~�`+�%i����L�ԑ�Ӵ���v����a������������o%|�=	o��^Fxxz�AF8�i�ծ'{�ޒ�S�6ɪrO��&�<qk8�X5�4w��֛����;�:��:��g�M��L
r+z*`o��ͤ����7I�v�ow����Jf�s���� #��a���SLf+�|!4�R�mQ{��U��){РZ}��*�C�s���a	�N��\k�=��(�E#?��rw�A��� 5�+Y�"�(-�bmR���̓M�{�<��k包�s����z���ȍ�����W� 	�X�n����7����������o��Q��Kx���3?.�w��zz��/������E����1�zJ���^}�����b��_^�_�L�~(i�uU�����)�\�0{2�sS�J��)i�o0�S��k������^�M�3f��2��,����]��Y��j�XRi��f�<�`���E�F�Y� f�H٨�q�� w���$��@�X�z���+n(�u_'%��%B�k���|*��*��H�v �����S`�:h-��� �b�6!p�،7D�`D'�i�]���N8�����N;�&'J�"㜨�I�h�6ʺ�TA�%�".4G�ܽ�����}U'O��(�$w���RKn�S̐c.�6Y`?tr� S�y�>�^�b&�x�	��\��\A\���U//(�M�?�� ����s���&�B���f����^W�c7��-a#�
�V�x�5����=H�'�2k�hDyІ�@�Q����[�3��B��p����hshƇ�_h��o�����'?2p>n�N�j��ޠ�#Z���j��dЎ�����o��d�\���2C�l�F��|]ƭ(��q�^aZ�*�s�>C�"�F1��tb4c5cdD
o��l����rN:��#Д����0p�*���)s���aΡ�9��K�b.z���i6�mvc�@p�ph0�|
�Z���&�e�@���J6��=�]��3���1���^��P�U�yv^<R�Z���h5��q �^�kz�'ְ~+��������Ç�����c<��7��.�Yb��e��\߭���^NOO�qH��,oW,��D��JT�U�B�8W��JD�є�hyg�vӺI\��B��J�6*xcguk�d��,��J�7҉꥛'�JK���o+ָ���Nݕ�e�m�l9x&��WE�vޠ�������M��P��=��_�sQ������l �@iڒ�J7�/. ���w)��t9��z�R'q"�@��:� �̆���\b���0��m*�QK��8�k�`"ܰ�$��? ��aEe_5E�C�჆�%���1�"F*C��{܊?C���B/F�Ս��q��s�xkY�D��╧����6H�A~��4[F�?�x� d��HE����?x��y{y�yA���h��Z�����~�=�E�Z�pg�D~D	>�8�}��lmO3�(����%�:G:f�Ww���YY9�G��Ywo��.�E2�K�����@pl�a���<e��Sj���؅��O��kn��κ�9���E��^�6����zѡ���F�2(��30

JvFU�Y�~��B���ܠ���d8�S����Ho����B������T��a�g��7��N���̢eFW�!�2�.��"Vn��R#�ڼ�;M�e��˼�^��3�k;���׌��Z횃��#�H
j�qR?�K��̈]��p��;�u�#N�Aκ*jȽ�_nijX���^�Œ粀�?����,�{w|�_��W��K����o�P&�nW��8�e~?~��0�{w�æ���7��&Xsò��Ր�W�#N�-�.�Ym��o<��+��m���t��z���!��O�X��W�UB������h���ϩ���\-��_b2/]|��í-C�n,����W��w����W�v���P��sD��&4v.4�������X�����^	9��bw��?��r+���A�T����k�"(�E�� �a���F
���cK7A�\ط��G�M�;�"���t���ר��qo���I-x�\L��@���潺���^Wh��@ܫ<u��Aq�,�X��t���Y��}Piy��x����.�]�y��6'����R �W���B�\^𸫡ZݠfH޶��7I�t���<l�zC!7Ӭy�����ׄr6�Bx��i��Iz0����#a�;3������*���*=i5�Cv���bƚg��0���;2�4(�f�u��s�Tai{С�U�(��@Xwz�96�	��p��C�l�.K8�f`k��/�_�����W��ْ�)�x'/����t���8 pV�夥���;**�ʜ�0n�FUi��}4åS U�6��
�ZD���ٕWVO��1j8z�^8�/h����ɼ��O�欶�:����c$�Jb=�����!zS�t�I�l{�y�?���� �G.�a;r�����$A<�n�C3��N�ةde��:�Hw��`�����ͿYd�����ey�_N��<}�5ٽjy�1_�O% ����b�}��_�����|�����vd�P���G��X��f��h8!�����n�m�	d�w�j�I�-#nl�B	.�sd^kf�C�D#!w�aRe�,�b�b�?�!9�a��1�6���S+��.=�nl�f�TO��C��+0I�
�<�FI�h�K}��+�B8�X��R,עG�j��J�p���V��{� ����?�.��yf��$�)�;B�#����
*ǫ�㡚���k��-q����͑-Z���"wAv�9�l�Rjq�j8 �ʜ�*^ h��fDqj�ddC�M�	��?���LP�n���Z��	x�����4���TҰ�z�D�fF��e"o��!��}�E��[w#�H&���uvZ�;���u���˕D��A�{9̛r�q|�y�;�W�7�y7q�[p��1�
�P�F}��0��憊ԥ�	���TƦ(��Pq w��5]N���Za�@����'�>�8��K	�*>�*������%kŬC��
a{&70k�q���p��,-]�m]��*���G��"Ζz0#2�yp����� *P���}"�YPB�n5��3����Q)�I;�r���)΋�����2��X�h��j�RW`[�F]Ng�=�d\��Ԩ�<:\�i4��H�Ȍ�[��`qs��	�R�m����
 ��e��F���e�,C����m|e!������fBS�`|d)�j�;k�8$u�$
��R��k��7D[&Ϟ?�LsFkHD}5:�&1�3k�K 8���g��g�����H���S3��,�拲��鼻�}�l�m����U���!��_�K�]���˸N_r�W���EeMO����d���伝γ.w�hO�pe5p�{_m+�{g��C]���6�79��Mx�ˬ��[�+��5�g�{)*1��P�@ќ�#3�.e�3��Z�֬��^T���{C���vv�\=�g�K*|�N�{-��Z�
�s�k����X^/
�28.x��lp���9��a�����bq�z�j��5�I��Z(ڽ�Uw��V9�:Ҕ��\���R58"m\k^��`�	���x�a��1Rټ�D���H ��頣���'��t��{x�QK���+S�k��=�1D���ܤo�4u�0�,{;�A�s(FJ�*�3Il�{�U�^����ж�K��c�O����F�˖��"K~�~m��:=�J����X`�i�d�� ���׳�X8Y-�X#.`B�関p���	4��K�?烬��A��3dނLF��-�P�O�u�s�;���-�"-7C񩣗o�xĔY_� �{n7/^���\���/��K��R��` d%�B�G3�c7��Xj EO���Z�b@�y1,&x�Eֳ��jT�Ҝ��2'�E��4ן�>�zյk[݇Nڢ���,��f�mx���|J+2Lm�G���cr��1jU���eF�y^x�+��"����l����]��~_�5�-%%'̘��J~�٢7�����ڵ�8}�ݘ���/��B��e�v�_,��/��t<��Ӕ����G�Я7�����ӍW�勁 ��b��Y���CUw�A�
]������f�5G�7���T!�usl�)s������7���H��,�����묗����Vt��x� >v�F��v���ϴ��ȊBNū�3s�$��!�0�arS!�[6-�o*�3-t|�aa���f�żj�!0co���	I9�~�Z�fz>l�������
�-{�o���]�E���@V�VU�/��5�l�R�.���8E�ࡺ��z�NAE�ymC������i�2Ӓ>�LG[��:��M,I��iTH4� C	��\�j��<�:c!�����n'��I��GcV���TI��](�5�T�F��-W�^T�P�R\�@�X��M0xN5��k�^)l�R�"�;�S�t� ����+J����e\��I+�ɈA�]�^ۚ/E�.\�2�|Y�I<<H��R����JP�"��t���/5�����9Ϲʯ�7M������;�=�a3HhU��0T�orHr��N�rrh�W�o�ߒ�z�����e��@��vy������Ϣ��e���AT�]Ǌ�մ)��ޒ�0e� O���҃��ү���j��L����X�f�Væ�5צ]eJ�� ����ݞ0B+`����l�25<?�F1U�N!�wa��c(�2n������*�o���&g�Ôٚcjs�Ϸꊬ�<d��p���Y�_��Af�0��N������(��?���!��5��z��@��}ݓ�_.�~x%��t���H�g�s�Y"�<#n�κj�\��j��Z}Zk�y���ÿ���s_�b����b�Hj����p:�a�[����b��l�+]�|7m�Iܣϝww n�$6���Þ1�.�_{\P]P炞j�,����}�
�j�-�= ���"~HT1cf&x�˩x�g�ۓ�,� ���_�lQ�FMT�(�������4Dsa�)�f�;f�R����U)ЋAsj����٪$�Z��Pj�ˌ9_5�5���U�5Pb�^����[�LYU���;�ژ�7ڔ�-3He((��S���|\��zb��z���j,rL��H�c�e�>�fr�{�.r��|I��5�5��r�H[�Y�����f��8��FSp����;����`G��QK�`
0m2g��!ܑ0FZ�;��OD$���`|���aZ=��dB�8�����Sj��������ӕ�2U��Y��ۜiV�R4�w�F;��hF��ٔ�a%˥v�\�eK �^KKP���)��A��r��(��#�qnTc
f�	���:q\w�}U(|�S�e^�G�
�_k��t~z���|v�]Ĕ[�*4��N��Q��$w���=4�&]5���'���9+(5ƀtƃ���(mV�/j��?Z�T����DC,Z«F�쾴[�r�h=�b���2��A�����^,ؼ<i��Ų{�|�?��b ������/RH������rxuW�O��p�6X���n0o&�J9h�`4��6ܢ�;�E�T����$7�i�z�b�s��C����d�~ּY�YoQ��;���� η ��>�ռ�zn���_��$�%�Nj�lY�`���(�q����ղ���ٰ6�8]�����_ɫ�D�k<���<�u=ɮ̻#�;�6�A]����q<)S�7�q��`�W{>�<�^_]�b���F��9.�[�S���kٻW)󟗵4���j�\�,�5���ê����Sÿxл�!Q����Q��a#v#W<��<��,ݲ�0�ؙ�z�ȓ"����F8*VܰA�f,K������ �^k�PG��j�V���Z��k�~�)��G�p��h���H/d�AO��ֻ@��Þ�º&����j�!_8	j(�t(+�)_��>�$���`�,{K��^�>-����y�����)�l�@�*n<t��k�p���w��\W4�{�;jgyoW��N��bH|��f�>(�J��#E(t'a-�{��x���c�̇2�����2�߳�C�=��_�8�\.EV\�ф(�x��[h#խ�>�A�s����^gk P��#Qcx,�O�14J��I�����:C�FK}�hA2'�S�T��,JlFͨ|�]���T�����/��Y������6*:fz��y���>�(�N����r�2;�7�C���d��Ǹ��dr��d:�dBn� ��-H?4>�
ָ�k�]�݄�{в�T,d�5�ja�P����^�:k�-�TE{��u5x{V�f�J����[E�pc@����/yX���zo!KO������wEi(���c�2(����/:_���e�����<�X>��7��}���?��˗r����H��x�[k/rL-��FmF�]x+3CX\��BL6�5��C0�}�J�j�n�[�U�Ì��E��\��z��/j�2�s�2!�˓�	6���  ��(�	�rMG��쵁�iJu� 2�({������LN�'|�!�J!�0k��܋��M]�zO���-B��^,���H*Ą���hB1�wW���~�t��=n'Dhj��H��ܯ�e�~P�c��!�ދ�P /�׈�l�j����TJ(�J�{Y���ԕ��h�l0�H	���F��8YjE�EANq^ߌ�'����?���d#Ϝ��	����u���[�n��O���uͲ���酘�x�^��T��h��S��H_15�ߧ��O_�r~'+�9�1��YRԸ�M�/�{+i�[���S�mܺ�Q���a��"Ug�v��ji����1K�{��C��T�u��'�*I;?�"�CB6��+t�1�^�@�0����Π�"�:�W*T\��%�2~Wˊ���S�6E�
�F3<E��e���;a2� �f����b�9M��ray*�x�{F��#�t�-�+��_2�u��W�fZ�8�?�2W��� �]U��Ԉ	��������A=�Z��r������O��lR���Dj�X��^6�q��u%�߫�s+�ţ��f����G#���_Ex�7�y�B�zF��F���l�f��`��V���
S�e|1��ꗴ�T�M^C.�@�`M��t�K:˵x�;z�څ	`%ҷ��l�_W�k`��0�+�D��Us5��ZUw���ɐ�bv��5̮�E�tRj3_I%\9�E�!+�y�Y�A�Ϻpԇ/:�Oҁd�m�'���%m0Z���9;Qs�S9�u���	�cC����|-�P���,ic�-#|�;`Q�����͍d�Q�5���D�N�g| �}���T�\�����%�^�E�o����S�A�US�̎a-�IM�hx���=�f
 9�.RG��|���LX��yR��e��	�Zd��9�e����<��K��)��,�B���d�Ժjz �fT����x��OGvΆ|s=Ίh
m>��I*7��܊���^$�B1��ӏ�B/��I��;&�~��>X�ԓ������si��s/��m�#�{UIg���4�<�5��q�5:��W��D7R�F�S��⍲D��B44+��:_�5������ƃ;�v�xR�ol|�ը��!�ֵ�K�(���U_��)�Ք���$�������1���[�q��:f��&^�o��e\���ڴ,6��Yǔ�K86d�7h^���YrUug��EZYWP+?c�&��'�jq���6�D-:��m���s��DVj'�mj�����m"�-M�D5�j��;@�7P}�O��n�v�7��(Fs�s�4q8�p�Ѯ��9��L��;pYhZy���4/^>�T�2��M�ZԣKy�۵Eu�1R�g֍5�Bnat��l�'"r�F����K��^�ΤOP�%=D���׉��m�l��mfX�sX6�Z��zs��9\�/��Bw4�S�s��Ra�Z�3���2(P�Q��շbp��]�EC�;4	v��Rk�1�E=v������H�k�>E=�$-�Y�Y�=t�Udu�ʗ:b;�ڣ��x�Rt9�Z����cɏ�� �O�殏�-{�@yG�R� �[�rH��2%b�kxD������qB|��U��%w{_�
�4:Ae�-:j�����U����0D�QC�.�U�j6Fd�ޡ�/�+%ș�[���H(Q?�T���1ƫM�c\�%=���jy�{� o�-G���ʉ��D������x���Te*t���*V���б��l��u�>��1����K�������+]ĕK���,5luJ]��T�k��D}3��1�!-4X�{�Zme�N����Q����~�y�P�����\qЛ:���a{S[�f�����)3x�9I�b�Cgr�#�pP��8	qG �A�%��dT3I1p	�v�Qe�=���bI�GQO&���^ƽ2�h��);Z�^��� �$����e�ު��o�+sg���i9fiHy�4�'�����Ud�1r�-�;��>�	�g��9�]k�]�)6O?�S f{�+�>�_8�4� B�)*�o͚'�.B��a�'�ZiT����kFY�P"�l^�������Z�w>�{h.�]_�sQR��v��M��`����s�G�~�U>6$�2GG-��$H*�n�O��j���rϹy��[d�om�U�W��e*[�4���#䦠0�Z�_�˜����h��O4�P�^���y���e�x���T�Us���g�u:X����n��u�y"������lF���ڢ3��{&U��KD�P���F�0��j�v��,�*�I������bYҵD�\�8��W� .����x�.2�B��K�'-=Pm~�+a�c���N�8nkIjtI�8��=��"iN��yP�i�����|4�1�M�w�W^���Tʀj\+��2��!<E�W��,�>(ۜ5�5��|��ӓuTZ�L�uVC� ��'�2!Xʴ�u}9��۷��o�][��H���t�xj�J�5�orP�����~H��y����������J[�	t���9�����T螇�]֠!��Lup�"��b���`����9K#4[�@*��`Z��Z�c��1���w�t�if�&.���ھ��4���	>[��֐OX�D9ٞh^�vÈx,.����-��{�m/��K(t ������ÑN!l'����$�K�e�����_oy�f����E���u�,�r�,�|fDdUJ&��&�8�Z~�� [nz� Թ�3�c_����{�ˇ���]�-o.��4!�~P�=�U�h�og�XH3%��Q��HqF����7c��{T:���һ7�a��а:Wm.�3�T<�� �������/J�м(��uR�
Q�{4����= �g��%3�@PT\�W��8�d��F�qԖ�=p��2��j=����d��+����[��{��ކYuL�+��
G-�A;߻�.ʚ�S�P�>� %H��A�������1��ԹGid@��9��-E�C��(��o��<�/y��(���Y+]X6������TCY��q�A2V��bڿ��]�j'5
��fP�Z{��[����Z��+����j���a��.ZX�5���an���z9�8�}�5���|p�b_��A}:�Gft�5�:Q['�)��c�Ot�MQ�x(t���5��3k�n�B�^�����4��7Mf��
dd̖re��3�U��;uF���S�7 u�4���wv jߝ=��u[7Ր��Em���X��j�:���L��i7��N�3xogL�*����, Ve�̄5U+�X>1��Ͳ	ղ�&p�y�=��ج�ؽ)�d�bo¯�-;#�sM����oW�z{!:)!wO����J�S
]ﱻyq#�3���o��S���N�u�j�QsE�����Dm4��|[���TVS�k]��pV0�\X���/ ��2�ҟ�����O�G.�����ox�����ɭ��Ɖy�®�\���B�h��y��Us��B�����љҎN"�=���l2�+�vQ�1޼��@���I�hHvd��a�SK��������nH�%;����Y�:�Y�ͨm��V�����O��u��$��/:T�\'/� pѽ��@Kւ�!^�!���ѭ��� �8_����MQiL-�I5��'�,'�����F#=&rVG���޲{��>zy[�3�O�p_{o����)�*�BS��2Ou��=�Z$�ys��>sтqT�cP�~9�.�������|6�G���{y����vd&�Z�tU�;�ᄓy�����F���(5���������{�7U9^���9>�h;R�J�D�����S�!v c����GH����W[��h���-f2�uh��K��/lݔǮ�a�����t��M��%*k�����X$:�,	Z~�����������4%��A��?qD�兼!�ߴ�+���ArM�6ewd�5o� @�e�?�k����u��n�u�&��1ED�mg����ք�ǎO��)���\��V�􎓆m��Z4����»�}�>[��� H��Fp��.Ys�:��	AX��H���9'5�ZAdN��p;���\}��u2��4�:�`�*`-nV�N�kf{�ME�k��ec���.�W-d�ls��>��\H�JO*4��Ž�' �,���;t�4(���,2b$E��dB�Ě��|ءMk��!�u-��Z�?|M4�����s�o�"*D� /C=깷X;���-KW�z����ޅ��bWe�J���3�m00	[U�.��+y���~u������b(ܽ"�BXic�F��O����@��1�8t/�M�on���C��\����h����ޜں�{��ޔ��1���UDIt���ǫ(��b�u���):�_/W9O�XT�|���������P@a���[��c����ɯS�ٍ��1k`����椦�����"�	���|�n�<p:��dS�jWx�7|q|t��'�<�փ�+MK��������p�%Ǫ�=�Ө�?&���tG.�9�b��:�t�rOM��T�����b�FPY��B��e�P�;�<����5��rR��$+uj)$�7�M���ɸ�T�5?%n��{����Yn��d�mYN���o�u-��,�q���@�k��I��j���b���d��5��i�
2 �Cq��`�,e�f#Fl��� Osy�Z�n"�.�թ������7�W��7를��`t���6���NĐ��Z�ǋ��S�P!^T@w�첵�$��)�K��t�vmv���s�C�u�:�ʎu�L�X��yV�e*m4�*����U��!�O�?�yN�7�ej�Lq��&��#����x��qhy�m(>Kjv��ﯼY�7k�ז�:N��9�u�Ϫ0�s�8��(%?�¨Mfg:5&�5�����؃g�Δ	�8h�U�+K����hS
��cq͐�0ߤ*nU�ye�BW���D�f.t웧�&�z�=B�wl�	��@������.܌�.�Շq��ȸQ��\�yY�3x��c�s��B�tr���i*��|�ӗ_J.?������#�]#{+^�ݣ*Tx��v5t�����<�͑�_|�Zt�sp�$�x�7o�U+���Q�s�fD��إ�q�'=�g�q�̽dN��E'����Lu�J��5��l��|Tm~�^$�q���t�ь��YBL��1A����o��.�r}z����s���ւzk��<n���1�������&T�Z[բ�������gC
�pb�u�s���iH��s�m�N�Я�Թ;���䣇O[�yօ���BK��?zv�hc��)[��>9�cQ�.U�^�'�f�u��:@P"o~�>3DO�T���� HaR��*>���A���Q��	���z��d�P�ZZ��^��H�bV O��k��S֒W�L��>6����`
ٵU�� �X�	.�k���T����D��@Y�H��s�S�gۯYs�@�/��uT��}�o�2[<��h��^�	��c+���E�!���-g��x���Bl{D^<����3H=O�)�A��).v&-c%���S���Y�8_AJ�P��!�>�.Zb
Q):��WOO��){K�V-QL.���SJݘl�����g.��q�ѧ�i��-#K���[:��L=E�e���v'P�Kf�K/Yˠ��9o�����F[��lNZƷNgF㰗�W��1D0�2�^)��O���"��x$�/OOdSŜX��л�]s��alo�^���؅~MuQ��}�f�\����a�x�4S�����Y�7j`[�����1���`kC/'��7'��B5���P��?��C����d\V��Z6-�#T%wZ���:��Е`6�ࣩ�c�ܢʧ	:(��$�|-F%B=g9��i��~�xSɄdp�!6!Ѽ�ҾT��/�`��!�=㩛�I^�Zۘޜ�n��p�M�&�:�F�J�dl �`�V�<yp�g��6��ã��}������n*�ȸ����V0e���	9��+����}�e_��+zI�*�Es��*�Ȗ�'6���NP��8/sA�q�.Ve���'礬M�se�^��jW/�}�.�a��:˪�W_T�F���.Q���5`sXC~m�5�csB�.G�i�K��tm-?W۰�jȬ�w���0`�T�sE) b ~�ݛ�L��6��!��fy��$)BXؕ�ꛒ�j��J5Y�k�)�X݆@�OlB�a}�ƨ��F�Q݆�v��s�Bq��wķ�r/�e�O|_NE��"�V��e4�����k���@���l\�B����YEpk>1�=g/uꗈ�닥�1�C�76��e~�QŮH��F��y����vņy-��r�F,(��XΤLV$�������|jb��"�o-���ZU�'��YB9����;�o�;��9?��L�H4��e�����\�����d�Ie=���yk��2jȇ����\/�H����q������j��>W�Q��J�}��j�;cb�r3���9�UYVI5:C��U��6�^��;��Jι!��Sg�(�Zw����ӥ?a��V���^�V�H�"�a�`����R�&\�ʈ�sq_�g�Q(��	�TF(t�8��Ud�z�]TZ�ƌd��x��F��M�ӻ��EK�Ue��=�mq���t�=����{��S��C�i����5Ёoܺk�h�Xd��8���">���٨�"c�˥�+j�͆A3�(�e�,eU�d5|��mDb�D6n��	�Us��J�C�0{NT	�1c`���A��=dޕ.�X�"��3u��Ϳ��0up+���i��l@6����k2wF*
,?J"���b���F{4쌶��ߕ�q�#��7
�f7{@�v���zdqnJ�[��������r�T_˭�OoU�**����`�&�TЈET���=m��5f�J���Ns�'�aqlJ�[��f4��k�zn}4��ހ7{��ą�&B�c���W%����hBY��A����^�t�̧"S�.�r(�X�A,DB�l�>ur�NV�J��RP��|.�j��"����͞�3�g��z!qr����k�����;��? �}��]��:�w�K����}���G����B�n4��W�i��ϛG5����S`&V��й��c��&��YGH��a3�ӎM�d3��V`�<�k+(�w���b6jZ�_HC��;zd�`�F������:�9��kx��e�\߈R�9�' �4x�B�5��ቻ��=Z�=9����s�����t���s�P}�ze�^�NG���~{�\���=�ݤy���_c�p$C��m������<��,r9'|R6$ ����n��d���m��R]-̥u�qc/������|�ڂ�\�y��m̭���Bwo��G���6v/�7���Q���T�,����H��#�U����(�~@/o�%�JAp��,����J��}��C����<�~GR�f/_�O���j%Gv����L�?��-���V���=�����/|���&�������N?����6˯�6���Ssw6�*'+u3*MOC��<�>T�J�����u7�>ro�w��Y?����.g4���)���#Zs�����._���\�/ܘ_�aKm~~{M����u(�y^h� ��B��f�@�����'t�f@!R� ���q��}�B�`Z�k J���O^2���P������J���s��Moϫ�j���jx��KV���[��,f!��}_�D<��/�/g�>q]��C��i획�0l��#Z��E6",���6�QJ쵞,�JE�2�)fӬ�ͤg<��(�l�9j�=��?>���s^ܟőϣ囌|$/��P����IjzU�a�5�7�_'����Q����0|��7��	�ȿ�������]����E���K�D�د��@♋��N �q�snJeET.F���o�Z��DJ�hD�TV��w	�AS�h�{�aC|��7�\O�m!JEs�u����e�q�yގe#q�Ǻ���戊|U�R�����.֒4g C�c�qI����1�^^Gg�W{��wk���ft�<S��~b�ޚ�'
j/I��9�����^Z��k��Y���sG���܌�d�
��IN������+�w`�u]�� ���y2�l���W3��Iޘ�U��d }�=�����V`h�E�Qۛ�J�`�t���C9_��LG�f�"OW���漸�S�,����k������ X�q
�d����E��	�LO��q5,��)����s� =�����W��I�q�ˌ~�De^�q�(l��d����V���\��mc��f��jP�h�D������T�������m�}Иs��9�}����q�Ĥ	�*��"Tj�����_��T(�*�TI�6UUTR����
A!iS�$�$`'q�q|�N��{�}��{�9Y��c̵�>�~�{Ϸ_�1�c��c�>/�1t�B�q�u�=�]x�Ơ_"X�Ew�f�g-#(Icǚ(�j�B�D��c�'��Tv���O�b�9쵵!GAc�b"���u4�����%#��Q\-�B�y����4L.ׅO7��^�
�B;��w�.��+c�M��������1�tḖ��(4����h���'-wt3���F$7��I�#�-�HL�fF�N?5]ł���7[j�T�0��#� � r��q��e���ۢQ�Y3�&�33������y1K1;����Ɣ��\6#� U�[C��T��HQ�@����\w;n��趚Y�r�ɯ���ū1�{g�I��6�u���J?8�]x�}�\ô�]�馝W��YQ��>�f��YX�<�YE�dAZ�k�:��d|�+%�{O�U>������J��,~���ٽ4�a|��>.&ĵ<*�����\��X�2�-��e��51��v�����+�na'1�?]P�H������ح ��N!���Q�s�`�I{�}�X�[�Z��t��3�b��d>�q�>_[��T�[�F��?��5�����/ҭ��ug\Q׮���
NâpW���h�Z��Y6�@I�퓺�80�lq|��\p�i�
�#J�դ�g�h\+��Y���!����mĚ�N���IK s��u��}�Ќ�%�
��ڔP?HEYj-Z�Brs��%�V�n2s��e�_����Q��h ���V�]�6�%e7���� CFٓF���iY�I*�OU�	��
j_�����"`Ò�{*1�=������]�9d|�nbT���h�p�#�i�&�x�c�X����?���0���ŝ_�ĹK����<G*8un�Q��s�}�Y�/ִF�n�axO��vX�;�փ��tӻ�7J���CȠ)Ow��ΩT�5؄08�Yc�۰:��{�A�����fD_�i��2v��U��0�6ޙE~�n�Z'Ԉ�o��7�����`��( #�=��q1Â�|��<�4�[l
{Ũ+5#�}x�X����qL���}qa4Ɓ_\֕�ĭ~rGJ��&��V'.�49���r3 ��v;y�,Ϝ�Z��޵�]ځ̜a69윀7�˝F|��4B_`"n�V�9#�tC�@�[~o���z �����i�=`^G|������\QK�P�CI�*����Q�f��]8�8����j]���^+����!u������%����V�(��r�0�E�0�i�b*��[K���63j��Z�����f�q�dj���#�)ƓX�3���������:7���R6p��G�(�NC��wT��R�u'�Q]L�3Ўj�ڔ��]�^&�ɻ���{�~��ǫ�ۈ���Ns4׉��lD��q��_"��T�j�\���#�������ALk�����Ê
,��̚�!#�2ݎ�W�\ڵhz*`�U�%d���?# ��E�kc0�⸎��ÞfC1�-�H�ܥĈ��.񹷑0��-��dk����]�/��8L�v�<f�=^�\�u}`+�hȃ V����0Q��%
�f�������X^�����܉�ee�|N���z�\d��܂i������V*e��a��|���.w�P4c��ֽ��Uq���l�g�c_m��7���:�=+7[U[\.N+���`����e��V3���͵��AƁf� �@��=��f�p)�2���iܮx���"��Ê�qL=!�X+�3�ft'L�yh*̊�Ϻܝ�G�;	}�cZ�Nk��D� `$@�q��H����q������S���h/}g�W�ݥY$�	�ȿ��Ђic�J3�5 =-�c�Y,W��3L��-������	�f	1+���
XpM���G�o2$�j�|���K%/�k�3(�|�Z�emC{�t46��2���@��׋��_���Y�pQ�ެp���"h�V#`��Ͻ�5bs������(��	�T��F�.�R��@�2<-��<H����=��ʝ y�)&_�ۆ��ݢ�v�ia�YG���o�ڣz!�+wf�e�\�ئ�][ϔ��Ev�4����{�J]P����v���FVO� ~u?$��Rv�ýy��Za��+A��"� bgA�Ҁ�"��royN�ֶE�qYd��#����GAP�JŘ�B�`!2�K���[LZ�a
>����lx�k��ժ��a�~�լ�E=��f����ƥ��L����x�gQT@����n���'� B�!qP�����4�b��� ���S;H�	��him]#.0#�Z&��юu]���ȭQ-�<X����s�>�g�5�� p��fm��0�e:mIr�	�|,���ik��f8h����s	ymqP� V�R�	eM;J��Yk}D�j�a�Ә5�3�86R��3f�=Sk:�섶혠�n"�͓.�D� �����4�B����U�g9]�ok�`/a�f�=6*^i@���Z�b$�"4%H.���NӏM��g��+��P_�9��^(��&J�T�KP%2����s�Կ�����t˛YS}L�Ե;�ۈ2���e����pÐ�t�$uD��NQ���`uŀ�[w=7482���ژ!LfZO@�"�~$Iw�}�Ih����#N�-ޠ�4`���@��bܪ���Uo�f��T-��Y �;���������y�Ǜq1����kh�Y�V
@���,�&[�J�5�Xs�6�y�LȜ�%+{ttjD��>�l�v��G
G�񩠐��|>QUP�܈�(��X�,'q�; ,(]�K	)�̤� �8�.i��pz*|����!�k����œ�j.Y����N�>,����j��1q��x6A�n�r��i�wgb�a�� ��oT�U�����z$���l��8nIﵮω�n�<��}8ϊY���Mg�����q�Mx"2�wD�Ϳ;�i���,^�.pW��NR;�$���Z����I|Cާ���#R%t�@sf��%?H�<�E$������ :u�h��n)Hޯ�н�_w�,��"ť�\��{7��4 �u3����i��d��:�g���ɭ͹Y�/n���� pz���'�o�^�ƚ�BaU�sg?�����n�h���'�6�ӳ�Q���Y�+|�X�`����_Z4Ff�m�*��7�j�#r��q ����w�`k���Q!H�,v�I�aM��f�XZ!k�c~t�Wj��e��j��
��]��ʧ��`��ڄK�O?q$��*�<zw�&V�RE��],͚eh�aA�	=��O�	�#K�k���������z-F�Z�#���|k	O ϠWy��`���k0���7��o��3���y�m�c�f"�r�q斩];�7{��UQډ30RP��������x���Y�Av��2���]Z�oRZ�@�G��rof��ks\>c�K�8=ZǏ��LU�e�µ8W�v�/[.��{��`)�"����t���ުR�����c]���������y� �u�]�:<:�4z>��R`^��p:����b��ʖ�A7��I{kI7Q!D	6^�J6��``�:� ��Wj���y�v͎��>�P*�	mC�j#�<M+_ԿT�!���\sʛ<�S�fĝ�w��%�@!=�<��.T��[Hz��Ͳn{Y;Ig�G��4�M�ϒ�dk�01�R�+� 6!���tuiz��ݏzBր��t���^�'[��1��w��`9�qVeQ�Yc
�����,���,ǿϨ-n��O��2w��dؾ�̹�0u�G��%�$��|�k�
��q�����t�HFk�R"Wz�	�*k�)�bz�����-&]�*!q�m�g5+V7*�J�iׇn�c�L�k}�z�u�F�`aL�k0�.�u�	��x6�^XZ������onT�������T~���E+\��t��b��Z.�ia�Ga�w��o��a{@S�w�]�-Js� �yŗ�����9�������{C�z����.��혩K�Izbh���b}�hq�Vw��P��5c��G��a�����hI�K��K�i��yP;m��LlYT.� @�F��kD�"�P�F�f���nv0���Q¯� !�q`��I�>�a�ȑ�it���������u���&`��_ ���b����|$H#q�o�8� �`U����|����W,]j����q�	�3S:J&:�"��֧!^�!x�y�)\.�Lg��M��߁ ?D %���D51>јM�q��G�F�)����Z����L1O6��0�p�\�+��axI���'��(R	����r����{�wt<�Zh1�	���e���e���h��<�3y�����.���>-��ӻ0b{��0�!�#s{DFg�>0fʖ	��{\��yuL�(,��Θ�2h�S��Z��+�s� ����!ɞ��Ip"�7q��"f\�7P_�iq3���Gm�;K�׳�׻�9rt{o�]v#�����·�Y֒ �-|�/�~���g�^-��[3�O%���F�"�cA '�<�_W�Bꑠ�w8���S#d��vtް»b����� ɿKᙖ�>�];��&���pԤ����E`,��TJu�är�S~��
�6��ถ�ň}au�Ƒ:���hv]|lf<�VR����sN�0��u�Ř���+y�9���L�a����I�R���>"�X�G@f��ū�T7~+A���̠��~��h�04�q6kAIa�֜� ������+ENnù�
���v:gÑ��k��9�l�*.w���H��j;�uS*��^��=����J��	��Q��̆�Q�Y��xp������1u)w*f�es!��Z ���ݵ�)�W�� ���4ֿJms�"����-�k&"�C�R��� ���x�C��z�A`i-}��	�U3�u�y�J8.�u�7��7�(|'q�2u��EF� \�,��Ѫm~Y;�tn����e ��I�ﬡ��j��t��>�ܵ�R1	Z�%@��^�w����J�����f���^�a��nx�E��^��k@�*8�=M�'���}^] �Qg�g+f+�������'wV��TLY����,+�
�P��ӣ.hlV��O��'��"��F��%�yF�D�畡��Q��`\S)D0Fri)�I�=j#�Ј���x�Z���!,�v�;~���	3����Z�&zGzF��:ޖw��i�������R�ŊDHY^�0����
"��1��br?_��!,����Ee��Z�}�x�J�Ɠߒ��.�K�/6{�����A�^JK�+����su;T�����c$��w1����X��� }X�np���� ���~q��D@_}���\lN;� ���I�E��(��{�;Msbߟ�&��-F�9�j!��&��Պ%�>f 9qWᔉ�X�s���M�#bB@G�a1J�]�(����>�� ���8hό8�n��Ҕ��x�6�$;�\��
=�CҴ�b��n����1�gߏ'�ة�w�Ҝ%�� ��2��@Ү�2��i�+ h*��xD�M�NG	��gk޵���PW�q.(��x�.�U;�us�ٳ�k)�E���\4��!����4o���YBd�����2����Z�@��Ҭ�s�֖�m�s��z03
f��в<��6&�Ŵ�6���-j�Z|�u��S(6�1anҶ�I�Ō�C���������t"�됬1/u3��bE�P������ыC��L
�EϚ�k��Na��w�3�� f%!tz��5a��qJiJ�>�&?�Z����`J� ���B��q�K!�u��'�>N�,2��[o�4���L�G�9���m�g���(�16>C��0�?s�0W��ҋ��G�?*KI�uIT&S	e-�,O�7��%
��\w��-�J�`V�G7?�!
��ӄ�C��E�!�=�> �n&r��b4�}"�k����n��V@�}�XP5N���vI�*yOK����������H�ͼۓV�b��^�3x���Ü*x�H���|!O�=�M��s�Ҟ���A��k�^T���,%���d#��W�t���~wRYF���Ýu�d뇔��b>fF?��լ>5���̋E�a}�^�Ҏ���������ʨ��ʄ3>��@�8�\K�����z�|?h�X��N��H?GaJ(l48�:6d^=��s=��	��5h$����e&^sC*�
n�Q"�7K�#W���ERM#���*�g���_����;.����U�pZ�D�X���ղ��,�P�?hZ��|B���@|����	��b�Η�d�	�#���<3w*�+��DM���\Da��m���f��V@��'H�(����3�AtqN��5�~50 �13���c\��Z3h���@q3z�T	�vճD���9,7;�`�V^�1Jܴ���!���hKb����=`N����º:|-"7���[��I'Ɂ֍WA̻�C�;Tfd�M
(ml�h�w�Vl�#����FC{)�o����y�V�o<^K׎b��z,��hu抙��|�6 �[w�h���Pn�e�����Ѿz������b���颦|���O]�*Iv���JѓD�:N����srC>�>_Y�2m�� �8�y�ZA��i�u2�ܕ����$��u��w���&s�Oi��m��6���&�n�_��:�������i�KVә�T�T���~�Q����Y[T֌�ř^C!�0
K�Z��z�R�dVU�X��r'V#$�1���LXXP�X���p.iA�ϲ�;&tu����˖�5h�*IGl��b�{HH���H�ڱ�y����9�:����i;��.U¸j?�j T�Y�b� ƌ��l��7M�C�"'��	Q��ɢh>�dD�9K�f��6	��KB��B�p���+�2s�<p��O�H��!Ee	��^n�KBɈ�ù[�j$d��(R �Z4�j/@�ԗ��V�fl"f>Y�Xh��n�w� !��̓���9�l�g!rZ����tuA�~;]�k��輐k3�ti�5*�ŉ^�]�g�C���tMɓ�SP�M�ݘ����h�L�JD�7AG��t�W!iw�U�%��fL*��H�݆j����a��'F�y��g���r9�k��D]w�YQ�+��gۣ%�1gMٙ��M�rww���z��U8i-�؊a�:e�L����G�kDN� �\�B��  �V�%���t�,�^�"P��O�����:U��r1�s:SU�����[g��')v�4eB��,������k��/�����Q��2�둾�{蹊W��4 �R�"�~X�v�=df�6Բ#��X��j�f8�h��AV�<<Vƅp�����m��A� N�C6u��ꎙ#	����sc�Y�:k�ZjR�gQ���-�h�[�m.���QD�$ؤ�YM�z�d�NXL��WH����_�K�3�̀��ʚ��ֻ�t�f��C�M�mhX�Q�&�s�S�k5�"��\�0�hzE͘RX��gr�*�8J��������C�:���-��!���^'�MՀ_����<��@D�?6/�S�-�6��u�{B����#[m��ќ*�[`�3�Q�^�GlS(�!����,̼r+C�?�_��n3�f����}��8:�AV��<֌��o�9�[+��|�v���Q�+�k��ǯ�d��m&�{�E7�-�;,Iqm�j��M\C�JE�Q08�#��bKp�`(���$�ǵ�ٓ2�������\�Pa��Rm^"����,����#j͢��j�2Ƨ�e��?��6�*,p��q�* 0��~�̼j�k($:�0������:@�-�}	f~���"���P�����g�h���Z�;��"�u�E܌�����ޭ
'Lc�VJ�M��E�L�h��p1���&�`��My�h������-89e���	a�E����_T���T4���1�N)��4����&�����'�m5���+��Ȉ+�8&(C*	�J7[�{���|���K��I(�oG����!���D�v���}SF�+�8BjR����JT̏H�'\L ����[@*6���Q���}M���=��}�N(��T��QNY�`�I^�2a�D�)$��k��]�m- ͥB``�ؙ�s�"�����'?٫H�u��7�{Z6����/q\g�����>�z���n�:�d���U
�2`������l�5�k���g��f
�� �s�5��k���8���/�"%i�<�=2�{����q���p2_�Tw;�/\̭�Ћ���|�#�ό����f��n�`�)�������q��9�a/L�S3c���R���G�S�>,ِ��>?�z�_��[�kz���S��5S;�F$}[$"�%�W�;W	�ě�Q��<��ݢ�	U(}ߛ%H�W���R�J����3&���˝��5yA"z��$^0a��BUԷ<+aBp��ު�#*�vc�
�t�QzFE�,z/�ܣdkhU�|i��S�6}��&��s7��x��c���=��@LH��>�1�FT[It�q�$/	�`��;Lm����Qp~0�<Y���K��B��f�����Ho��7O���tѨ��o���	�1��QJ>t�f�N��:aF��݂3Y�ٱUj&�IX4��L��W�G�:�Uql���R��jz���㾪�D�,i]Y�F��2ФjE)�$�:r��t�u|yǥ�k5Z���\�0���m��\� �w�2"�q_�����9<$n�9�1��И���˵Ҝ2���эg�B�!���
8�&��|U�&{�����̍V�)��R"��4w�=�>��F�K:�^���ٞ�q�uf��-qK�:!e2�q/�u�9�5J���-�ס�"�C{i�
Xo(�����	��
���k����Vz�ݼ!���T����0X��h�J�|���*n�|�\Wdn�=,�U��"��ϳ��U���>�Z)>�%d�i)y�������Z��?b^FܻJ2����ɢK[�&�H�Y^$4�&�K'�W�?ؐ�z�X���\k9=]A!�\c�xZ}]�@�|D4���&o��g�ʈdU)Z
ZkE�h��إ�Xҙ���o��ʠ�Ήq�wS7�i/�R�P�N��0�|��%L.#�����MP�/5�l� 2���&b�Q׈1����@��5"*V3���C���aL�w��7�ڜ�g���]�Hf�����Q����jy��̐�- U��vg�:��P{Ȳ�eI����C%��dyٶ��^D*	� �_D�*��@P�$m��������]C�K"�9�b�u��H\td���+�}4�$б"�(�?�4�:HNO�>WÇ���I�]d���T-�c�,�������L�����T���ր��V��d����/��J��v�@X��?ܪ[w�D�Qud��$�O���"@g�Ʈ4��XL�@|K�)~?�BKf��Ǽ:,��\��C�q��@e�´2_���D&�5�I���Y��Ц������$��|*�|���*kb��/�|��8�N�"~�N�sJ�Hx��>@�l�w�  �h���M�S.��Ϻ0�̠�:�C����K�`�
ģ�c�鉑��t*�K�ț��a��Jeϲ���D�K�j�M_r�t޹��h��l0��{��ӲSŌn]����M�B���bV�I���d�rJ���/֨�ӯ�t���'�m�� M��h͌��7��0��o�ف!D×�8:0�1�٩��#���a�����w3�kXnba����}Y�b�ikSib!E5(��˒���иH�&���H:�Da�,jB�$(m�TP���2�����
h1Z��h��F�����Y1�6��t�ݙz�O���s���F� ����#�`ܢ��B(���W2�l0t����뗙 �oc�N���*�\)i�0�e��tA�ga��Hf
iM���}��X����-�rI�MG��)�-���h�b��dunrҢ){� �>���v�E^O˴)�J<�8LPsz���2����ή���b�K�{�%���t"v��$h����=�D4^��ɜ�W%d.(K��-M�g,����r���Ͼ%i/�N�2��ė�&�;�����J�Ĳ���{�-���>sn����;����vz�����/ݵ�����.���)��&�	A
����a�w�b��^���3��]����L�p�-�)����� #�iy�����*_���	�hc�}O&&dR!P=�&r���x�})�Mэ��D�[�L��Y�Z��YM8*#A
V�R�cWW�#�=ʚ����u��x��U����)�ަ�.T��`��K��	� t��Q��k�����ha����!����L���ʄ�W�QXva�!��jc誙Ë!�6�	Ü��ʺ4�ϖ���n��.� �֙��ސ�V�s�*���r��a����`)`���<���k�$+��������m�1b���N�i��N�9_�-�L��꥜"W�.��ԉ�6k�'��
|6��n0��9,��{���R�z�΢J__�K��#�3S+۬�Ě�*�R�-(��GC=aj��f阭�+c��&X���ʟ�+]wSU�n"�j��&�� �(pc�ĉ�� [��Ť�`��J�.��H!\��7���QX)|�u�Y���h����Uk����(�B��V���Kd�J,�{i3��hw��f8Sc�H��l��r�;қ��#������f������2~z���dy���´������?���|����C�_y韨������������DL�j�Sm�Y䞘�d�^Y�@I��KD6uT*s-�S�S��#���� @k���=d�5#́+�F��muO
�J"F���a1�/Cc~�ya���47��EI=��9�Fq����c�@s��UC��j�z�\> ���3(��S^�C�ZE7N�1b�ܡϢ��&�*8�,)�G�E$��ZĻr�h��T�&ΚGŖ"�BR�K�H��Ղ){;�bk��eܾ�r�L���9�^�1�e�M�6K75[�
E3��Y��*
J����� �r��}�t7.[ʭB5k�/t�]���&���׉}G���w���[����%"��Я�TmJ�y��.V a�d����T�=YM��'��BS�$x��K�kJ�b��Y^U��f�^��̈́VߓE|������}�� �Eq���'o��ƒ�]���AB�v8��Z�_W^)�d��X�i���w��}kɐ��kx��߸)��W��ˎk<����5�9���G����^�����_�ly�����߲,z�/|�SG:�>���o�����/|�7����8>~������~z�l��e��pJ�LC-��ՈnW�P|����)r�K�|F�J��QN3�&Gi7�g͡�(�h�Sr,�6 ����!��|��Y/EMWa- �� �v�ficC��L]o�,�C˯��`�IB�dV��B�o���F�(�Z�M��(6�b5���M���7F���mi3��)�Ѽ^ete��޵��yf�0�>�l|�JᑠЌd�?W��3��Z�ϊ��w���`r�kJ���++"����8����׎5#�����=�z��@d�4�&�w�L��@@�Y/2��g`��,���2��1���Ю��l,G��ަ��\��dX�FBk�pt�+t���c�u5wnZiOc��1�����X����o}~�V��T\�������`�������F��Z�� �.�::
5Ñ�jJ�+��� \�rc���]�]���E�Y�,�b�WǮ���Z����P��f���|w����m-� ,��g�(r�܉}Y�����s�Z�����^��=���u��|������ }����;��a,��ȯГ����ϧ�������ku����������O~O�,�i6K��e<�G=c9��SMkU����I�TS���:yw�D-o�Qt�k�P!#�x}_�O"���,�^&Q�o4� �����'�@�=.
�=$D0v�3L���)-�+p�(#G�v�pDc�9ԯ�F$���1	�I�9��c�c�}����>[(��Օ��&�p��%��!I=kf荎3�	w֮5fuꦝXl�ᰴ\�`�J�|���g�'2�NG���|���Í.���#k}< ��K�^��+]E�mfkG�'f.\5���8Rb')|��pL\��vݹR"��2'L���V����nF�c�}صG`,#��m���k��+���x�� ��8�L�����b�cƠ�������;�����x�ީ�F~<�S{r���XV���Y�9:5b/�����|�`
|��F��5}�v��K���)��w�a�=JzM`���$�o�����4醦k�#_�:��{���\�S�b�m�n�e��7�G/�n���ۻG����O~����������>�iǝ����������K�ŗ��w��{~�/����ѿs��{>>��O��ߋTί� �`'��
z()aM)f�S�lf_  �IDAT��g5�Iw�"����.����~B�����n:Of,NhJD�n�ɣ���y��m ��Q�QW~���VL��]�&� Ƴ���OV����X
����ؤ�ƈ@�hJ�q7X�ð{�`�1�>;�D���[�_|��HCp(	�ڒY����i.��ťЊ�&�-�\<��|���GP�������?��-WU��zT�Kn�5!�f�Yg�0{ ��ī��Xc�4s#'.�J�hoO��u��UgzN+1^ujfAW�iǶ\��U7G�tG8��=�K��3�5C��ٖ�p��|4{�O�Uva�];�����:s�Z�m�:��������ߏ�t~�x�f~������vh�8��ą0�n�h};:Ȩ����
���~��]J��kCBĕ�| m��vzp}ש#��:9Cww�Bj�h���5s6�/R7�f�N�{U+z5Y��y��Go��������������G?���;�&�e�_W��<z����w��^����������O�W~�<����/��G�_)��Tc�d�������v��J�~�Z�������,�O͂!� ���ݸ$.lZ{`H}��k����M�7~��S�p5]E$~�R��q^$>lTj�4t��},&�M/���cg�� ��Γd�y�MC3��:�[E���ta	X\�'�׸n}Ctd�-��	�1o��d��lo��0'%��2�tJB�cq&$���:Y�.��g�w�=�R�\��+!q�.Dmb�y?z��P�����$�(���T�O��}�$�l�1x�~2��rP�����V�-d�1��KORT�4��9R0T��s��-k��#�&)�Y	���kF�2�ofNb��<��Z�V8,V�K|f�H;�ȳ�Z��v�T���۬�<�\�?��~@݉��hF���B�{8	5�1V$���d���z�ƴ����x!̇tm��I-����$�Y,����S�0t���z8#������KQ�Eh�����s�pw�܏������/���Gw��k������6���_��w����g��G�^����Ͽ�ߛizy��Ov�ףE�.��� K*&�����:�y,:�W�ڣ9����k����ڡs �a^s+��n;�"�)ļtiM3��q.&R.��*l���l:k��C4����~�JP�Y�L�lC%AgRdҪ\E��j���;5'��-�ᬱ�m�u�k�(]�H{%sN���W��X�������r��u����z�Q�g���.D5E6���d��VO�W��e���s<�vN������F��v��;��1�� ��,L�̂��*u���ي�4�;L�\ϟ�>�XA+]�~~M3�e�]�JL��#��A��G��I�f~~J�t/=�%���'��{�}��$fQ�M1�OE�7	���!Q�����"-p�Si�Ji��\Z�i��.���6�� ȣ��;�]���#pB1h�U�Bݬ��*H�i�R��@%W&�s���Ȓ�uGf.L@��HV���R�f.M	,��Q�?BQ��|/����	��ۡ��^�YJ��U&""0))5�vW>����m�}��1��d�X3�u������
���*t��7��<S�4M�,%R9P���Vn�L�^�Ӈ��?��w������"��]�NO9��p����_(����z��s��>|x�~���n�����ҝj�&Nt�sa���"���Q7T4�X#- C�'��{����с�\�8�!R۱����5�^F�f��:@��IkMSǇ�RH����?xM��I|�IC3Sd1IQk�G�#��� j�.&eڒ"J�dݐR-%��k���ՋWA܈Q�����2��klנEj����:�b�b.k��Q#�81u]ߢ��o�ϵ���U3?��%Bh�ᒶ0_qk����u� A���5�ɖ��=闿�4[[Q��Fi����S� �	e���
|�<N�1@�C͊�.p�!� ~G�V0#~Քͱe|��q��5�$�q6�\1�㌏�Z�@�F�?�nF�g��@�K)xZbipuh3�֭5%���ZӘ��9��-_yjxl�� !H`��?�րhE�f����ᭉPJ���1�6�С�5&5ܪv�����VN{Rf4X,I�0�i�0	=6��iz��I�)ڡ�����	!�@����x���Zlr�/��a�Ь�_>	]%�+�����&z[D
E��R���l�H�W71<T'LVYꈣ������+�ԥ-���i���Q43F��X���=���OM�y��:�g>�~���O��k�鹷��:d�8��>�������~��5���O�1=m�y~\����ߞ�ﺩߐ	��w��,��� �p��$,5�2@׊^\f֢e����g}�������J�h�*�m�}ۯf��6j\+���`�������@=6�1�QZ�)o@����J���gG餡�1i3QHڄe�� x�!�����e }��^��;��H�Ecl-��w���D,J���FkM*[a4ʝ��{/r�N��H�2H��O�T������k0(onIa� #1�Q��o��a�;������CѾ���y�̤��ᴚ�UH���E�F�iRw��� +
d- B��t-䦾ah�b�# �Ǘb��R�`�Ó�Ǝ�\���X�X�fB�Č{��/�ܩ��*f����q���|Uw�y>/�dc̋y:6m���T(n�ڒ Fi��Y����]�зaC��[×L�#��b����XX���Xp����0�W��Fs�?��x�b������%��'kv�BQBê�@-jYU3��F7���g���^����C�����ߩ���7җ:^C���oz}���ɀ�������ٟ��O�/�щ��H�R���=�������"�nT-i�IT�匉���V̵����+��4f�Nk9�+9��>�i�d�#/4 �h�C�ޑ� ��mL���;(X��77fiOp�}��E�V�
���I��T�Ĥ1��,n�vf�@�B����2UY��'ن�I\Q�z59�7�5���T�l�#��0.3���b<���ML�,�8�U�9��E�@Y��ςQ��^���\0���p����=^C�~6�{q!�}�E�we\�;7�IE!Ŧ�J��s�2؉f3Uc��kK�����cMW4����s|u>�W���]���9hQN���ؕ~����i�Nu�I���`6٣v����,Z$��F`�lX�S|�M��s�ék~t�����V�`����@�]s�X��8.�R:�]	0�Ep�(�Q���횬�ӊ��ȍ�!Q��DN�Oy�N"�Ռ>�^�ʟ$�د�o\lf�;����<�>��˳?�v�oz������:�[g�>��?~��k��2л��}>���i-�f1��TC�z�F��Pr�~SSx��Q'�_�xH0����7,�M��%�/�x���e8Gir�IA��\gу�/�<l��5�Y`���fj	��W1̩��,37I��A�Z���cs�S�V�ӱ'7��6@�Da�S�����
���Ip(��-a��,�:fs7��P�I�'����i>_�n�Z�L硦I�g�+�,&!�#�%����D���,*>rBк�׀Y���d���@(�N�q������dt�
�}�n���P����z�I�'�ps��ijB�z㳭���IM��OZ�L��zeܰ�oY�΁o[���täj���CCW�>�WL�M��<� �{@�a��%��!��0�4�\�FPW`�'�f���Y���݅���?`JҽѮ���)�?�o�U��l�v��-[���
��nM!��@���4"+N�Ч1IM�L��f���;�\�OЭ|/G�=���n���=�=�C���g��7�����_6C�C����I���?�������֟_&����ā2��e�`>LA�c��:pJ�%��޴i@�8Q����&�-d�i����9u�C'����m�C��(�o�.��R��8��c6���U��{�,����TB�NV���"r�t[��O0td����Է��o�2���<L�SM�8J�@*����m��a���!
��1l�f�~:�ܕ�ZE-k˫���7����"<3WL��\K!2֪�q�*�P�>������,2���MƑ�#������`¶���j���4JKYq&�;ES���v�Zz1f%��
@���&"�;?w��`Cv��``��6'�vu��Cp8����o^�^�ԇ1��Y7˷�׮9Z���C8h"�O��B�ե��MJ�	ꬁ�]�i���X��d�v���ԍ��{Pm����?��xu
�`>���'���[Ҟ&M�U7��a��ٝW�ػk�!u�Q����bj�IT{�b2e����VUek2��9�O�~u����������������=�A_��1t��L�����������G�y�"]/W���il�1��räѱ�-_�,
�{���j�U���Q3$\1���Ř�^��h�� 08|>p�6"u&!\2t%�-��͂�ҹn�p���DCԠ�b�E2ӽ0r[t5B1������D�+C`�L�&P��0�*��60A�������10�����h�n��y��LxXKb��Q�g���D��mg��ee��jD��n^76��6Ĉ1@M�]5Jd;���f�ւ j��o�1�J����t�c
�'��/�|��{�#�@��f�p�n�-�F��z'ʹ\��]Ts��ߌ�Iz���&�Ɔ0bxk>�f�o1�/q��;��ۥС�6���P��oԎA�v�����|Q�K�A��Q�z��s��+Vt�3����oi5���m��K1���K�Ef��qF�Gky6���P3����ڄ��j�mX" �r��Y��	�Xm#���;oy-�tH#�Hb���k>�NR����3��^x��V�[���1}��W��_��o��~�7���������ߟ��N���6k�/J���mJ���MӰ �K�D7r��Wgէ�J��ɺ6f��ߊ���p�s>J�w��-��"��<�a�q�2I�H+#/�����̌��hT`�v%2�XȋuSmb&"��l̤�6�k�(I���+��L?�a��&cj���͎��V�
ps��������p4����[)&��)���=������Ka��*��l�V��No��VB%4��"�=�����C�}ݛ��U��a[~?꠩�F6���v�g�B�
Ke0'�ܲIX��Y*��խ�\�F]��^;pM��M���m2ʎ`Ä¼2�����^�������;�ay�!�3q�KL�Y��� Df
�2��|G|�>!�Ä��}S{7��q�a5C(1q��	h,;�oґ˃2܆���"l)�`I*ˑ1�*Q�2�Ɉ`�6�X_��h;�$(/F�{�)��U!��4���YXҒP�ߓ��_��~!4��h����[Bk7���%hV��$���>�^������Sf��,�
#7�����x���o�����=����ߚ���羚���:o\���?�K���_�7���~�����>�C�\�ʽ\��iX�{�\R�J�#m8 ��@tf�B��`� �Vw�bC,�%�m�����6�(��Tb�3V�}��A:/�.k)w�
Y���jK��<Ka'<�jlk���]b��k)Iz��w�7n�`�_�ّ���ݘ:L�	��6���Q(�*��Ã1� ٭!A�y]�y<݈��~_�z��}��r�''��6�G4[`u��fF�0W��veR�l0h�>�����9T��1$s�H���mV<�HB ��f�S#B��`f�IV�5�
x((���� k��V%w*�����Z�ō����JW5#����_,E�TP1��1<k��.�by]z��]�x���g�}dV�i��{�!)��3�'�V׀h�f�h���;�.������{�l��*X��[:O&�j��J!Dv�N��MZ[�|��i�'��M�G�8U+��!*5Ł39����=�6U�90ԒR0��S��Ҧ}&8%��
y<��L�"(�`�Y���U�
�M�?4�u�⸞�	Ӹ�&r�y@��(z�Vt��x��έ����H�;��ŏ:���ED96L�nZ���w����������5o������5�����_C�����z��O�'?�y�腿���]���G���܎sq�KL�yqgʦ�)�}U�wVBքZe"�.`b�ǖ_l������}�#��ĭ����3�0.-ia.����@��'���(��*�B`�Ʋ?/����H�5k����K�t�K�)^��v2f��Q�`�Ed}(�i�6�kƗX����9>��^e�nY<�8��Y��M�x��)SŰ�#j5`�I����h��c\v�m����ʅt������p-(�^3tנ$�:>y'01�ca�����\(�7��/�Z��y��b9SS�\��jvlpE���.�>�	����/�X���t��������!0[�c>>U�K�4�Ӡ,�;���Ǒa��ʐb�S�s	����7�^E��o��c'q�Χ#u�~��[4�t�e�����g��3"��qpl�)�-h ,��t{3�^��w4�بiaӅ���5C�
wF^�/�C�>F�_��%>a']��X�ئ�ۻ)��n~����_�����"����M�����_5CǄ?��.s|��ͣg���6��ϧ�_��!<�)� ��ԏ���R��TȂ�	ȩCW�cD�w�,J��60^��͕���\j3����B����A��#u3V�A\g�cH��ƶ�t&�e�Y�0�cR5� �u���cU)����ѻ܆�������S�J��:��!��]�O07b< D�M�[�Q�fŵ="�R�$w��~��̟��:4+�Z5�Rc	!I��vhx�
M�,�Y�w�.��J �0��)��B�pu����3��iU%(�W&��Uh"+��1Ɋ�_+n�"�ۙ[�.�4�IN5�Ά03�q��H f�k��
<�1	6��s���-=	������ɴ�&U��QH�)�����v� ]�����J� ��kB~�:��O��.����"�h�)M�L�0�A�����݂˧e��'�������H���Ee�is�=�t'R �僀���lЙ1�9;�1?T��C����T/�Ǻ\��99~-$�Sq+���_+<;K��b.��j謼�ɓ�c�l�s������?�����ߥ��7�����:���������2��������M��{��������H�'���f��,_��^"��s�	�(�֦Qded�@��ȍ8ۙF�bѲ��D�m���AW��m�m;'"���#i��@��PQ+���6NaV��b�(��m�֛����΁7��L�	�/$\̳��:%�6��.];hB_���'��}����T�x>��k���C?r�5#�n�%/L���I���Oi3a��A��I��T�;�VZ������f~J�	�ȵV�閒��	m�Y*2�5�f{J��Z����z�����9�Y<�;���i-v���8��R���(Ym�|�ҸV]/eǈ��G�@�3�����k�,�W�>u�̓�lM<�u����
M\�jc��9Z����1���ʭ[#aM�X]9Z�%aZV����<����Z�t�óM_q���"��#N8�����Y����'����4[@"��Ѹǻ�Ňj��� 5k���A�����2�c-d\3ů�E e���{C��of~#���'<M��q\�^��u�dw��ov��S����
�������1t>�������L��l�(��"�}S�@D̈� Dbt9�t׵��g)g>�ɧ��D����?��f��g����>Pd���+���F��pO��5nb;ɾBP� ��Kmq��L�a���b=0^����k���}���ǤxEW�>��H�3�Ey��`͑�tiMd]֓��¶��6�гb�P�<��qٜ�g�{z�����ip� ��a~_��Z���.\'��%|�� !�U����Y�2�Ԅ!�\�"�j�L��@dR���B�+��"��#{j�v�&����R�=N;��D�b��G���GS��0g�a�}�����SR錉�B��]��UK�S�S�紕i��c'½D]��I��nF�+x����I6C����\1��[�E��2�XO�A8u����Si�hV�ЧJ�����V^Եҥ��N�m�O��|�zsG����r�|�s�f!��ZD�!�S��,|f����.��b6K~?���|)��n�Y���|X���[�â��q�kDγ�<��Ks���A���s�ɝ(.ӧÂއ�����{;�r��oz}���)C����>-ƾ����8�;���TΏ4��[k�F0pt 1�����Q�ś-W������8��f�&M�j�(�����ơL��f�	���2	�~͐2qE|��DZ6Q�t�Q��%�EY{00�����inBk�o����0+�� ��1mŉ��W����6�J�q'��䫣d�YC}|���N�'Ҟ�0�v0�Ƒ�������K��2t-�%�a*$g�U�J�-��X�و��{H�pa�L�O�s�u#TEK�� -_�������5a��j����S�9��M+V�����p'V��D��|gBC��T�Uf��:Y�o�&�U0�V#��:N��s*lI�!ÿJ�ݰO3�L@�@`�"�S2�,:}�}���(��([C�a��1���0�mY���Ь@�f;0��c8o��>�f�^��*��.�}���Oď���t���p�Q���+�8&��
du��1
ݛ���	�C��G|�y�=�9մV���3Y�x�k+怏k���A��g13��i����m�BE[�rN:��-L�c���ͧ���=��.�}}|���}����?�n���v�?Q{��K9�!�3�Y4@m�v�ཆ��{�Qw[��Q�U�-��w�`<H��8�(�"R"��R��������e��d6%x�>C�
�o����f�V[�ig.��k}����^}i��x�7R�T��D�:�r� ;2eQ��T�m���4�I���v{���檀I0(���*�����XCkp��nH���i�
Y%�CXh�5Ba��Q�0�G[�3��w�CۣRCohn�RI�<I�O&���H�p��	PY���	�ac�L�`�HeC%:���P	8��M�#zc��N�p�'�q��`�VŃ��3��q�b��pd�EYΘf�{0�UaN4=��������If�]�Me����@`][���f=�S��H����w��%��%ѭ=�JZ�@�%~�n7E��?
0i��u�%lK���gV����)֏�٘��d'��
�0�ݣg��V�==y�%:��[�ᶉ5�YbEK�J���\�
��!�A����%�3��y�����9bs�L��Εv��z����[�9�i��i�)���3���Ci3wQc�p[��R�k��s�Wf��/N��?t��}���\��ks|�:�}�{���W�m�;_�Ŀ�����w,0�6��=�I�ڮRK桐�.q����t#O�r��T�j�#u#��:��I��%��,��&���m =f���0\#@��^C�2�3n��K����kE� ��tO�*V�cWn����R;�?�ӱ�,fR6�I��pMflf�-���+o�Ό��m3��0�4>�{:������r�tKu���l���TV��:��U9Y�C0q.}7�RNU|�'6AΓ�z'��_�8�g��*�˳�
d�S��'*�)�l$��������S�#H�Qr�F|%N�g�
 '֬8#_i�|ޝ�)��	a���5�n���k��
8�΍=8��,=���Ls!d�R);��rLիL�p4ۺϊ��!P��=�2������q��v��CA-DbL��#�{�GE�o�_��.����uy3W�=f��Y�UF^�Q�0��*=\���~6�U�R��|RZ����0ef ��TA0f�x�v�qz9��nXC\��x�1~A���,��%ca������ځfX�-+��|�`�#��d?8#݄�ȯ��͚�?�x�����P.K]��+���iv*�V�OlO���R�2AT�a)g�����5��.�S��p�C��sLVN��v�s�wg��_�}�����6��-��ua�||�'~����t���������~�·g�� _�j`@�fJ��ZE*�4m6 >�3���&��oVŝ��~Bp��^��]@4��/fu��� ����m������m:Q�r6Q�"��?⮠��Y���gL��F���Y�0�Q��I�Ed����H��[�WG 3��0� ��i��/����FR�%D�<V�Of�QF��n������y5�����pAȨ3sumn:����d�n�>����||�Z�M��)�, Z�����E!Pj��)e����j(�,G�PX3:/�5�{�b:H�Ct0t(m=�'�����T-�\��F�Z[b�0_g���Ws|5G��P�	f�Kn�����,�Y=��$�3�G\�~-�u^5O�7y��\��=�A^�I}��0�P��=�Wr�f���๾��4G�x�px ^���+���$Ѡ\�,��X��v��J�����Z=�MȪ�0�\�}��R1g�@3�7����"@����E[��G��?�����{/}=��C����P}�S�8�����X��?N���ʵ�HL�����b�J��˻���$9��Y]�ޡ]���/�	�R�ȓ�Z��k]�Nc͓u�Z ��M\�Gjc�ƈ� ͚�G�	�`�\þ�s����̆ȳG��eW��-����d�r�t\�3�fib?��0���%y.�Z�j钺�5�y���6���*���Q*�b�B�y˒�
b~Nu��eGb�֔���*���<\�}���2�����9
#����}�%��|�<m\��Si�e��oi�hD\3f�p	Z:=pd�G��%����A���T�ӓ�z��&���"�Y��n��#�Q�fe�K�:��[D�2z3�'���Xm)�]�G�Q�"����֝2Xg`����ڱ��f-]_�kꭅ@�`7��>h�aɪF3�b
c��`������Hy[q˙/voע��J?�������o���3�d&��!����W��0��v߸�g[�֣]��D35R�4ձ\��]@��!/}>2S^j������Z���]��ښ ��/��b��[�����eg&�I�y�y\��4�o~�q��~�;�z_7�����E^{�����ӟ|�����g�N�������X�}���v̱v�<�V@�f����"9��];.��f�`�=cK1G`���c����_�z'��[I�d�.��4�ۂ�-�(�gT`�t{�;r6%��h4�B�OR�+n݊)O
�q��YL��y4�F��3CKU��'G�;hu���Cw�;�]���5�D%m4א,������M����س�|^���Y[��.��*~x^㳚yĬ6�J�V�ִg�'8�v8k���U��1�;_�Å@�a��$GF�K�{�w�4\�6�93��L"���)���M�i�s���2�Oiw<��]:$�`c����nX�҆E�>W�f�K�W�X�D�yM �$�$��-.8f�{u�|�̔��	-\!&�Z�jw�x64ʊ)��SZ1��"p�E�Ͼ `����87F�,"|5�:��,{�M�z�h�����(��̻X�͒k��0
O(T�4ǣtZ���JWi��f%�3�kʶ���
r��.J�y`�9�Iig��l���F8p����O��}.���ϫ2re��7'�s����8M����Ox_��}_]񘇎�C������::<��/�O|��,���/0y�DS�E󛔉��=�c�EtJ*�1����̻#4��Gf�L�LIׂy㛮G%�&Q4����iP.�i��3Af.K���׌�ivS1%D�	I�H���,�Nz!릉b#͢��_��!�Z�����"��Ԛ��k/�L��][��v7�4B�Eb�=�w��/w��)��ر�&�[��=�o�ŧ}y�c�&!�g���|߽N���Fʭ(%9@l�bG��F�Y��c.Zꘉ��@�o���5G*C��`d��B�^J䑩)�
`(д
�,�)��՗Xw�f��"k3oO�.r�I;���j!�����%B�n�\<�a����v�ϼ���_�9m}�͵%�'�B�3_=3�:�U&�P�T�G׽�﹒P�q�_�ԃD��^ph�M�5����pĻ2k)�k�iU<��������N,��}��$�a.<s�Jr|kf斁$�M�1�K�}V�h.��n�..]�b{�\];ZB[�52z-��5�"]�!v�D=����ۚ�#xSt|/��$o�q���}е"���w���[��_�}��g���������3�R��>����t��}�//J�?�H��R�6�3i�M+�RA��Q�����s�F��fk�SB��؄>�G)]��`� vg�N��!���\Ւ4�˝��s���o@���cD��,&�&���>Z\��L>�S�N�����izM���%Z��N��E���~9!�
�D9k�V�����bN:��&K%�5���y�:�����8C�p�NF؏`h%�L�5i���qa�e�ιj�^��5�Zj�Ko��_34�/��n���ay���[xҠ$>9Yh'n�"��E3R*�<��!�s�.0�R��dx�H�L�"f�L�ʑ	�:��O�[E5��{*˟��L0�*��L�j�T_g��Qj�]C�u�9�k�m!�^|���-���|�}LAM8�0������&v���I>��*��}��ձ��5@��OӀ˩@���\I�2k�糬A� (-�Z �)�"]�drT�'�vՒp�]q��5 C�V�����
N���"\#:6�)Z�~3����I�j��H��\4t,U��,�gv�pB�dM��#��@�jQ����V���1H�-���N�/.~��ܻ�����}|4t��������ş{qz���D���$��-�XU.� GD�FeMY4SmɝSM�J��ҧ��C���������MߏRY�D��s:5�_CWd��&6Yw%��tj�5T�`��BFLͤ�L�DÔF#]��{��'VN�d�U��$�4���H1I��G"��W�)Ҍ��_K��:�=�o黑�g�/����ߙ/ lMza����r�+�N_�h�Yk�kᜪp,��Hk�kmr��n&z�k���Z�������))?w�㒯���_���:h���'ZI�Mx�hc����7v�:`����nfo��	ڟa�Yk��\[*x*^�d��3��K׸��߰劥B�࡙vW��/[��p�I&B���f��%r��j�����Aq�!�zt嬸`Z ����w��$�Dd"��A+��O��#������-V�C -b=��鄈�"��8'����}�-��S��K�d��R"������22��� H��pݰ���/.�qf��ƥA�a����O��M+�V����1;������gir�z�X.�����H�����u`�nu���d
*ǁд��e#��/�އ���g�������7�����}��׿�)��*��o,���K;�-��0Aʓz�E����),i��Q�U[*�O{������� ��9�y��2�g�G�jM�0�5jRDF!F=�$8�g�5�,��u�!;I��c;�=K�b{�!i�2�RLL���;2��Y��$�$T�V#vB�w��Y>8p�� �SW��ޡ�[�Xl���<X�����a��U�p� x���g!/%*_������ŭ �U�[̘�ҹ�~��+mO/�G���'^N�-4��h��nγfV����wt{7��e� z�	��y��L��L7�I
�D�8��d3�a�B������T��ا��}�@D��N�ST��.m��%H�8��H{�K����r����'Rⶋ�{'- ���t��]?�᧍K�!����@�
��ʙ#�#荿�&8�>�8$m���_�yˉ�մ�N.0�P^,�ք
��kB_��4b#T�fݭX�#��'��1Ip��N��c}�R=��l�d�"���3gr!����e,su!D��X���Ҡ�.A�Uc-��BK��-VDr���p��8W2�Z�L"R^�ޭ%\w�B�e��5�\Cg`t��[
�eAA!P!sf�������<Оb�#1#��ig�G�'�������4E�8}�n�u����������}��7����7����o����/3�N��ۿ���=�����0	2GB�?�(��E" �����������]�V���t���F:�(��V�{W6���U�Q���5k�y��M���r��|����>N�G	�	]h����NBT�@¡^�E'���^�}�������*��q�C�M�B����&�}��@v]�u��'^$S��s�W�@B�+
�d�t'1\N� ����<=��i!
;�/���O�C?�u�_g@I	�Bjs�� [���c�UP�&������ih��Z��* ��@:�z����K��X`B�^���F�k��ɛ�(���V Ø�"���ڔ룖^���S��C�)����������Z���~/׼U��4�5?{��1��'�́������*�t�+�؃��1�$9���.Y�d��X.gv�
�LښS`׺��Z/<b\��ي�0=�ׂP���r �K�,2#�fP9�ߔ�����0�{%���Y�nD1Edx>Y��B��y�
�Z�����iO�u�D!�s�mvߦ���Z�)]p#I5��h�<W�[�w����ǥ���ݳo�������K�:�a��o���/�������O�6�w!i�נ��Y|�-Ȍ=��b�^���AcQ��ms��I���ދRw�����Tb3wՒ:�lML*�eb����M�JLE��lr?qj�4�>��礔_%jKC��jJ\�gl��{��/����)�Q��l׶��[�����ݴJ9jh�q���}��oK�}��z�dF��ˁ�!̳ᓦ��F~����j�F'��!���7R��1ccT|镧�7ӳ��1͂˞jP�k����,n�Yq�~�� �~v�^)��'X�6���s���^"^K�B��E�;׺ꤘÂ�q�̟<a�F�ŒYe�ZDLr��2a�#z�](�&���|����M��YK�1
�B��;k͌�%���ZDB�X;�
:�w��}T��k�ɘ���'�I�U��?[$H-�p���l�?��Q�~�<��$�q�<Dk4�D�Jv�-B��p��� �{+�{М���͸�T=��-{�,{j�Bռ�Lڮjt`�5פGk&�=UXơN��w,)n�Z���bL�:��8U��T_oj�f��A��&�ql��N7���~wf�������u|C:ǧO�4�~��{�������L*��*�`�~�چn�j@���_��i}��FV�k;%dv�L)�M1���-`fi�7H��Y��\I)�j(I`DQTD�I��J�fM�$�eA���⤂�"�l�p�L��$3�j�j1�r)p��km�#��!$�c�5q?i6QTS9�E��1c�n�K�%u�;��[:;�BO8��o��bm����yY�����NZ�hR)R��J م�"���H����/}�C
��>81P��c-ڠ(�N'H��I[I�ڮʖDR2EʒxI�rxn{���c���9�>�v�P�����������6p���{䁅*�%v*-K-�8]/����i��yj}a��8��|o]�S
�H����oJGٺ.�
�̊���@����8Ѿ�F:	�?�?��fQ�$��⮒�EU�7��U.u�$��\���
��[���bN�������>{7�tyy��q&׬�r��2�I[�g�}$ga�I�5��X�ܽ��z���z�e･+�I{#���lU+�L���I��N�dn1�ų�	t�䦊�x
nM��}O�N���@����r����V�͓b�,2��d�9�H���t�7)/���m�ˈn�n�]�D�F�A��)!���Px������h��"��+�~�?�4� �'��y����������n�O�A~,&s[��w��dBD+���4�Wn&�MB�}6�-�{�h��]���C�L5C�u��z���Z�ZNb�Y��X�z��+O�ɜnЄ0����4Z�����U�@��H�ĭ����._Q�	@�y�:��O�����d'($Fb����u�

H�J"X���&&v�21K��>Z��%,i��h�4deG�5��"��X��j����U����8^w!;i�u� ��Sb�Wtʲ�\精JHaz?�'��(��,V�Q8j8��u�\/�e��B���}�FoA�{/)M���uy|i"e[G�vV���1�:�˾�7Eb�<���)E)�����v#��_���ngF�SI�i�{w�%���c�9�3���8ȥ������ᾍYdB�> V����F�S�dI�%i�z��}(�^��ۼt\�Nי5��Uw�<�{�MV�F���Q���LY�<��k6�����)M����\�8^���Q+rg���B��F�$#��JkΣ(��P�B��wx���.V_�����ӊ�?pB'�'��7^�*�ůB��O��?�~�N:�ѠxH��LN���d�0�۠��Sk�֛��	фɁ_�m��[�w\�a
�/�5�sL	��U]�l��?|ә�y�=5�� =tlY}y������U��8Ȫd���7����RӜ'ʲb�m����� ���N[J���3N�q��e{\(�
�����-��.�� ��I��J��A�}�)���Q���[�Î��1QԣA-dxn	)A5��IEI3W�t�)M�+
����-kz�:�ߧ��TASr�͕9�9ۃA��%��S�K�����\Z<nO*�Q���qF�VS�q<K;h����'���0.!�>�s%��� �D������a� 푄�a
yk�"H:@�*d?�"��9Y�B���lѰ��>"���z�N�ٜ��JsOeM4o>���9g��8�@c:�%�n��_S�̔
j(�ݍ�N{�ŵ�?X�w_�L�����}ʫh���?��Q	�9�I��4'ɔ1��ߧv��Gg`Xf�D$�ͳ
lO��{��a����lK��(Qc��$5)_��n ��kxS�e��5���!t�=�~������o)�X��?�J�>Є�*k7*s�)���%i���YJ���þ}:�>J�B�Ek�czH���Ff)���cL泿��!�q+wV!�	���ロq1q��q3f�؅b`��$�`��K�,����Q�T��تC�Iq��T� M�&�ȣ����,�AW��W���e���1g�`ݷT9PT�c�O�)�4
�A�7oѲ��ER�+q��v��o��e��Ls�q��������Ш�ԉ�@ٳ�F=)6x�wܪXr,F�~�0��g6.���I�A	ko]�>��kLi�YQ0���Sᚵ$J�u�@����2��N�D��(��Q�%��8��t�����v��<���1������|�5{<k�C)c��Dnc�#�ȱ4�Ŕ�[�Ρܿ��i�HѫM��`-`����W(���u�"7H\�ŷ�7ރpR�K�\*�g}�S&����	ux[4H�wm`��]���םt/�̙�����X<02.��4�V_�Mv�c6�/����b�n�>���$��ae��b�P��U���^'�%�P�Q���<�`
k1� FS~4�F]Z��MAcE�ǟ��=r��4M
��܀f��������P�a���:'|`�~��	�q!�'�v_�+�[��<Aٳ)QRW�]�@kա���/�u�}����&�A���Xx�A+\&����ݪЊ���$�4`������ؠ*�#���s�=�O)���4!Y�H�If�/���8$�5Ťdnnv!�D��aP���:�>���2@��\S��4� ��,���0�Ʃ��3i���X	u��+���2�J�/�qԬ�՚����6lx�\"�J�4��u��{�D=>u��D�
[}�<��b�(;�^'��$�\�]�Xi�ѩ�P�>�����\l2O'c5iς�z�t���Z�I� O҃Q�X]�U��'�)
Z)#���R�i��|j@҉�d~y!(C:��.�j��Z�J���4�k��g����^"#á$4�^�2$��M}[#��"��Z�����T1���!�+٧�{'N?�Q�$J��ΥRB�����/�_ϼ��M����%���� 7'j�C����.M�Y.����d��d釪!��	���9Ú:�I�Pi=�`���n���z����r��PԖəȼ��M�|jSP����5-.�\�r^��FOTQpJ�zZA�����`�H��h�(fc�Sԁi��/7m�]�7q՛BcW7��P>��	�.b%��y�7�uiHC$O#S��]�z��[��?��6��p>(|`�~��'��?xN�����������/������%��k4��4;�R��u���ZtP�w�ԥ9�V�HW�m��-�؉Uez�޳�
T�2�%����B�Xד�K�Πپ ��]�6��"�k�l�$_T�G,/��`u�r��j��B�+�N��_"�Mq��e��k$�1�:j��
�zu�3]%:B�q?�@E��i��hh��R��,����C9�z�ht��w���,�ɿ��������ٚ�T�#!M�&b�k��GF#�?��y��zL��V�j�\_>+5�(n>�m��b���5��<zk&�s������j��zZ�8Ϙ�o�o�G`e1��wPWi��K��a}MQ*��Qq.��}KeX�m?*@�Xt���\��F�^�7�C�_�ە�\qF/�;9S���g{�ɮ�R�D%>kώ�[�|��Ǟ��'/*�{���L�V�Q��i(H]-�\��p	&y���:$�n'�+)�-Z�4G=������=y�
_�2s��G����ۓ��X���:��B�1��:�q��"<�7f�O=�0��<vz��&���ͮ���π�4��1.}��j/m_�p������k��%�L�>0B'<��S��+�.][�]S�]�����OQ:T}��]cMa����Y�(Y�Z��-y1�����"��ķ�<#��L��L�I���I��_�t���?�U~���X�t��˛�}�1W���u�l�V�е)��I�8&9e0�I�JcYY��4�����[�θNa,	+Bu�Շ�n-C-��� ��Ne�Z| ��B�6IR�n�� �}��5��8��	�C�~�n���>W�]��7�_A?�(Z�`��O�^��FnLS&ƾ�c�q�%Y\�j=��յ4��:����~�[(��V��H|��%��8���N�^�pe$ZM�0�� {
ְC���cix"�iw��̪_�{
�<e�:N��e�d+O��x&��a�TT�P� ���YH=���|-���SZ�Nd�(�V�9QԸ�疆I2��n#��	�.ԥ2�n����h`��9ю�� ���h��dD*]�Z�T:Fqx�����ܰ���u�Öd�'�/�C�S"���d� X��B?�0��U�I��yN�a�ӊ�d�T&��;�%kIn�!������ڻj�9�8�i'7;��?�����o���k�>�C�(G��J�߽ ���l�� ,��nH����D�Ik�w�ĸy�T ��-ɤ��tr-����Wj��q�2��r7��D>jז�P�B��L�畿퐗����f�J6��mD�k����)�
����&=�눦�Q�g:���K,�T�;W��Zƒu�*y"����(j�Y�d���;l��al�i���3+;�X�b��SB���fT렄��+D�[\�MGd�-c��zM�)4DN=�:�µkW����^�訞�]���BCB�
={�����2٫\��J�C���
�btn�Vl�5��k&d2Z���R��t��Iv�F�dL�Y�$o6uA�61W����qtM���K`&}>.��z�4�����$�Irc�׮�#7����o�K	VerkĲ�B�EY,���k�\��O�"�k*k������?v����:��+��8i���p�>�d�B�N��"�i��PO	e�kG6.{�D�+X,� �`�9�A.t�v��kR:j9������6Eɱ���魨���s�s�'�������],͵8�d�q�i�&���5���(��7��=.n�^�Z_��N1u"r�2����_=��~�������'�4|���	�ޏ^����B�^���m�����z�C!e A�8C�Aݕ*�6S�+����%n��'i�g�v�o�)Li���4� 
Q���=����UL�n���O(�>	O��R�M!(.�L�$�I6y�E�f�m`m�e�V��A]��]�J cR{����ikI��$ܭ�`��o$�\˙�� T�ݲe��V`�FژG%�j*�ز>o��EA���%t!Z�⑩$<n�Zq�ry]��%{�����{޹���1���1^�c����Z��b
�2OJ�(D��k�L����I,2�u#-����nl5=�P��"_�z��
��F��M��#���-N��սU��w��n�Jf1��K��[J�/���$��]�:�͖���uI�q�q��Ե%����I	��:�P\���Öm}�^��0	w�]��:%�5H����9M�
��V�e{ۄA�(PRIc2$g�+ٗ6���I�;�f���
�mu���� �$���s\C�O<{c*#\�48y'��;�Pb��佯_\ir��<�������JO������"�����c��(*��W7}��y�ik��ҵP��\/�;�LLCY��5W�<&�@�=��-Z��j���a�[5�p��>4>pB'<�ħ���/|.^x�~���zI�P%�[�LbKNj�ԅ��Z�dnVw|����Wvg����<����w�b�������a�&�=mz����h��cuS�W&tv�Ic��6�r���ꁐזNh|�A�.���V�-]�E
���dN������ř�
��o(Zn�Ĕ�Kָ|�X-ԥg�:%{������h�Z��������RU�f$Ƕ��$��VE!�Z��ΰ��޺��[W��`	yQ�+�ť�9�.�ҬC�#g�q�9UE��r�F��e�7�"5[Hc^ۣi|��w�w�o�dHw�J�.�����b�U��>���zdm�)��Lt�6I���w��MI\�r�)�����EnL�I�~t]��KhI��]���e���=mߕ.7����qE��5�/��A,�M�c#!�����+��1db�Y��}oϙ$�ir%-���ȺF�g�R�d�^�X��4��%��j��[�2��J'��E� �ܔ3= hY��y��~Sh�v�D{496���e6�^�vN8�������d����R��-yF�{o!ç��ͪ��+P��ȍ�̓*�ҵ�*8�r:��.�N��H�i��6�'c�������h���gӪY��>l?��Ϫ�i���\�Ąb��b[/�<
Mj,������<����3w�~�����a�o�2峏6���F尫D���SM9�� ���q���zCɌ�E�#���t��r�*�q�6h�t��l.t��;V���h�L,���Ժ���
eC�3VHS�2�e�A�K7Y�l�z�'�$▭:\�t8C�$��"�r��YZ��O������vKB�*'Ȓok�|���j���a��i�ꦂ&�˔��C�ʁb!�l�,�(<CIpl�I��m�`�ض�H��v�q|��K��d��}�\�J�7:ɫ��B&���}D���S�4�;���ico9K:�V��J�l���<'�*X�ps�ۚ���w�I��&ɘ4;��Awj9�b:=���uP�>s�3���Q�;��d	�Akι�� #Q9+�:��\�g���T@B��F�ޓ*��B�_	+�*W��h�R̝���w,h�"�9,�q�e��gQ�s	C��v�AP~�m�?/疔���e��NVr��2[�{2B >�l�wFA� �7��e/Fk ��|�z9[�q����������:���Q�]p[�]�?�{����U\�_�}/j�U�6r���q��R�f�Rc�,�#��S��'�`ԺWM ���qSw��Q#ڸ�ޔ���12G�0nA�,���1�F��t#�c,�O�Af`%���d�Z�a��*h��J���?N����(2�%���C`"��ǂ��A�(d�1-�k�o��*Q��@<RJ�5����2c�E��aD~h. U)��U��N�
��.���O����f1�%]��C��=Z�в[��v�I��$Yk�4��n����bm�w:�U�B��f1�������a�8��xC�ߏ�	V��ٖ��9�bR��7��ra�1��0�kѪY�屧,[�+7���J�ܼ9�v�ބJb�9�װr�a�Z�,q݁�A�YQ�4' J�'ae�K!�J˱����K��(��#4�Xs�A`K��^U[�vtTN'�9�i��`����,��M�=@�[2[��)%�(M�,�n�*T���AW��ؔ� qd���hb]R�@�pJR۱�T/��хp��H���Cc�����a&e��"��5OĿ�mВ_�K�*]$�x�h.: ���:c�)6�K��PuU��?W;O���n�M\Vc�xI4�ڋ"bJ��f�Tʂ��U�^�0Q�V�|F|N*9?�9Y�0&}N���^7-W�C���R�Zr�/�/��������gg�����n'�V�N���O�+_�2����E��e\��qH���&+I��<��~�Lw*��Q���x).ҏ*��FLP�#�6^�i��1w���ܻ�@��1��ݫ�d����S����-�iK��4�^�OU���*l�w�=���/{��Cę
Ӓ���j���3��� j[�<Y��a��Y#u��뜅r@YHTz� Y{��G,�K^���J֨�-��ф�]	CHc�n?�۞(y�zt,�m�h�JYS�������.��H�5I��+}��_�x���f�cܲ\��W�/��W��QQ��V�3�7�2߯�,�uȏ�˙�"�}�ʥ�\�0�"?W�N%��*8�R���{��@�R'�����V1�<��mɸ@�.��h�K|��ǵF=kV�i}�y/�v�:s�N�b�oUMΩab��Ɇ�\�.Ӑ�=g�'#d�ܕ'��S�똊G)�(:�ne�]=���ȑc�n�{j�+�,��%�R���v.�o��C �qD-YJ@��u��I�Mq�y;;"UR�kQش�,X� ���^3X��}(l_���i
�����PY\�����N5�ԐJ����E��CX�u���r��zE��F���b4q�y�\��$�X�պ�śh���P}�'?����9���x�O�k���������/�*��&}]$Mo�DX�轕j�4ԥب���:l�K��]Ǐ�#~��|����	#�}��V+dn� �{%i�aZgb6W�4+���|��.1zq�rIP]+!NZ�ir-٫�h���l��R����Cd8}d�DՒ��?2�E�!��?k԰X���͠*B�.�����{� ���$$��������u&���z�ԉ�a�Ꮊ�i�A"mZ�^����J�-m"���Xيl�|R���C(��+3w�`8���J��-�
�uގ8��T �+�_�n�.1�~�h��3�T���+��}>]�qK�YJ�wb}$�2��Eʍ�%{���:tM��9u�WAz�GU�J�@I�,T��^A^�P]��-�J�L�+�QsRc�2fA��ɳ��9�|�f��s�dM�������HF)i�:mV�� S#�r���G�^.�dܩt$�FB� ���i$�Ž6�3B���Tz�_�Z�S�j��щ)򽤿���Q��T��<LZ< ���-%���0����Z�(be�q��i/�s9�(��Xʨ�u�S3 ���&cG%֪��}n��` �EP	2���%���Y�W<�3�g�Z=Wt[C9 �+P/1����m��w�=x�����ے�	=����<��|�կ��O!�ZF����u)�I|7K�G�SѲ!�x���N�y��jY�`��;R�7�]1M*�Uʁ5IPE(�N��2����^�o��H].��$F-/r�U�.B(e@��TTg�6f)z�@b+��`]�Q"���*.�����u�ЊF\�M���x�D�CF���R��PVm�l��*4G�{Ɏ�����<=�M�ǣ�@n��uL�f;��;J*X�nzq-���C�1�'j�E��w�v�����x��䚫�L��o�H�b����� w�+XU��ϟ�2{M�-F�FTմ=�����|+�^�q�&�g(Jb�t�Dʺ7�
�J.�rԎx��3�lu��5V�2���U�)�D�٢\,�}�'�,'h��C�3�!��3�f��B"���Rڎjx�n�l/�qWX�%Tu��ƽ6�[���ɂ\����i����F,��5�?d�
��~M��fz�,��(�;��K�,"2�����J���-���RA�����o �A��	��9潑-X�5�H�Ѧ������_&�Q�&���(�%"�=9v�NUVQ�ίT�؃�=���.(�AcI����N�µ�=S�ሢ�{I;r�4���+(6N�-syZ��j��cH�7��_�����6�W�=�p;�%�z���ϯ@����C�?�/���?��gC�|��ǆ�� 
����$@�����֮d�W6�>N4e���ׁQ��Xڧ��m�wy����$��..A;�j�f�`����ԗ�,�`��3D�����*����|
��$ӂ�_�7��SR����͚`WpP��Z��%V�3�CT�!m�-��@�XIR�t��И5k��HV�l�CqMN�IcW� ���hIqRQ]��%#�ѦCa��~p0��t(ܨ��%�d����IHl��Jb��t��Ԍs��E�2�{��PB�^�����\��Z�J�eܧ��L��]g�k
�7���0�F�������ⵃZ6����H#y-�$�8��Ϣ�d��K=4� Ւ�փ�e�t'7gn��� �0�9��K��5%&�Ui֒�~�	���19|ڗ������)ד�,�O��19�^u$����T����j�������^嘵v�:�6���E��	�=,���ZR�j�O�f�	�LT�C���Ʌ��a
o���> "��I�8�4KnJ�� ,��D@���|ǩ�3UO��q�G��fYy�dY����?��-���\���@5�6h��<�|%��cbŻ�F1m�7��vI|[��ڠ���ј��a���7ˇd �m�ۖ�Y|�y8^�w�}.����I�^jQ��HO���C�Ƣ>��?&�$ǉrE��=�荹���d��n7���D����`�.��h��t4�¶�*JҊ�b)�RwwaWq�	���I	'$��͏�Y��5g��T�����,�54H�Q{�S�N�U^_�c^�Ѭ�&�����3Z%<a��W2�tDx�;�噄N��TŁ��� C񺌖7e���V���	.�3��I�Ww�( D���d0Tx�U��� �*B��Ư��O-�0;|��]�d��m5%0�2w���q�P��!�g{���d�۾�mkC�w�ޞԘs�Lً�uk��F��6I;��Z���{b͉�����L9-e�"�n��HP�ӾZ���Ui��@�A�#���A88#V9�zck-�Ӊb�`��i�&͸&�ǀV�M���U�v6o�H줎X��������D�Ǜ��!-0/Tֽ��}���G	��-�m���j�35�$\RI�'
/� �6�l��x 7��v�B�9�aG���r�q�*J�8U�?a��3 xhL��@��A	m���P}`J�����X�)7�ph��qw�����XVc�>�J��_�\��e��be^�M޳h�ǦfoFl�ȑ�c���j��c��w(�^�f�����O}nWܶ�N�z����P���֟�ׯ���M�#A����EU7 Iz��%���Y�>ђ/�]i2�%�A� L0䱄l�v��k�6uф-b��64 ST�byۈ�8r��q&�;+Y�pbA�d.1�ʬi����c�f���$�O I���$�
����3H�-�zm������ɪR�z���3�*Q]��#��e�o��hw4�ɯDC.J"t"\��G��A��*����RAM%y�mwx.����h-�C��H�ڎ���p�~ 3_$�ɵ�h���j��!�۝�}��ys48�u�y�<>�|��3�D,,��NvKj9������
E�!�CY3]Iι�V=�<�i	�*REԵ�h�!Y�e-J���F��B�Z,`���A۱��B\f�myźi����Tޟ�J�z��2�%�H����� ���b�ɉ�3iX��QL�a3��\�O��'e��7({/G\^OϬY�Q=2Y�P����
!�\ͻ3�sȹ�p��DJ-�zɌ�G���˝�}j"e��j��=��{�ۭ��P2�%a���R=�$����/�+X"m�Ŵ[�I�9��b	�lR���;}w�+0z�FQV�h��M������cA����>�0>є$�Už����TR02W��p�H�5��|�z4W��r�B�.�D��oլ�/:$�\U˟�Cz�r��nw�քn���O3�߸�\���g��������!4?��Ie�S��#$Gc�<���9�b� �U�U�2m�-��!Z�n�ʈz���Y7����J2vp�;&Vݧ�c��ц"p��������~G�+'j�]1���A\���k�߭UI	�5Qc�Ԓ�s4��F-
���!n�v��V�����غbwk�b��+{���'P��.^��=�q],ީ�0��ȵ�+ֳ�ܐ�̍I�\7H�[��\Ԇ�h��.�0Z-Y�H.�Z=��s���`��jA�׀\�76'���X-8Y�d�w��U���%T��ג��sE@b����"-��Y�GgP9�a�e?�d�h@I���n�0�=6Z5�	�L<�5���ֹ���s�xr� ��:ƽ�
�j��O-�$|?���Ru2��C��FؤDp�ZK��
�J��l������ZA<<i}��׮f���^k8E�kU�wH��a�~�C�!/�hF�Bk�#�2ds��W�ְ�Gr����V��\�����Ӽ%S��D�y���I�,I���
g�:Vd���Ǧ��G�RP�]σAHq��O�q��'�-�V�m@{8�~$��C�A��-�r"p��̳0���kv�x�H~�"4��EA�KaHN��*S����*�n�TH>����LHk\=�&+��
���aYD�?�"?�'�j�0�2��]Q<���V��Gqm��\w(�i�������	<��!�	�#�@���g�����z���C�Z]���B��'��-����J&�����"n�G$��PmZ�.��`�m�\�<��S����jYVy.����r7�:���TTy;ZU\sJ�6j�H�s�� �vF�>)�UK�k �:r������l���H���G2'�Fk�}���9���X��Ζ��Zk�Ce�N�����oL�Wm���X;�B�AR�
��E��p������.��Ξ�g�(�q]47�b�~␥��NvN�oT���5s�k�ъ	h=-�^���.q$�6���E�B䤣�	$vj��F�v|�Z>xz]���^Q$��T�E��zy?z8��q�,��Q���e[�1����p�)F�R��Qq��~��ِ�k_�U>��t_�}�d������<��T�f���M���O
MF�A�"�E�t�%O��uK��-��r-�w^�>[�k�Q�q�k�G \��Xq���Zs��4����j��p�����S�9��%��W�R�{1w�ZH�hl'��&q7�hw�bFY�I��d��6n��^,4�Uh�u�%�tpB���Ǘý����!i�y;�%�����Xն/���|Ơ�"Q�[i����r>J��
�j[��Y�:��CDJ����l�C�|4����=U�%ᶳ|v��	W:i�f�QbŀY�0�H�玨S�Ԭ�gMA�Q�{Z%��C�a=b{!��G/ʤ�B��0sJ�kv:{���5؜��j���nu�9Y!RWr���]��l˟�o\���{o�'��?w
�B'<��O�+��[p��5��ۻ���_T!��!�3�.rS��I�[�Q�vu۳�*k��ˤ��n\M"�Q���z��c�C��E""-�,�m�V��e�ns���� h�%)U�M�� G��I��c��JL�W	�H��Įa�~Fb���fyJ�9r�#*�X2�7p� ��~�]���#�5J�.����]6�Y��D���c5�HDQ;�|wH�<�hN�(Ԯ�G���jl7��k��*�u�8���u8IC7p"`�y�(uӲʋ%~�~�3�U��9��<Z�QP���w&��A&�H�Y����Q��E4�A�Ȃ�e��(�"�����mW�t��G����l�Ӿ�4��%�dE�p^���t�0����7���AY}=�(�.D]�&�Fk0AVV��aZU0L	[���1�(�$��p�uv�C�l��5D�Vl״��PO��!-I��Z-�;�pDb�j�"*��rW���B�ˣ���2�Y��� ������#!$`�d&P�~5H.^'Zbʽ����Q�V����U]m�.Ħ���#�-���)��7��v��+۴��Ks_]�����JH��Lu�vx�jT�������TNH��j���zsX�sV���Ð�R�V��W�\.q?��=4�q1�:=�\�Kwy#����Q41q������ቅ�����9���k�.�-d��iv$��<��*fu�P�zr4���H٠�<��5^a�B%��h��F\*��(x�{�ʆ����Xvb��.�ZF)�g"���J�ь.{��g�Wb�V���Q��Q�X�bY�I|�+�BI|!^�f���,����1}�������ٳx�"t�C��,o�7��ē�_��O��V�O�e�yLÉė��Q��q��D+Oba|��Lgس�'km��PJ
��Z�Z-��>Z�&2o]�&��nQ�p�8$��e��]� vF+}�b��#�wx���-#J<�i��sſsc��<b�H� q/���%�Y����Z� '�v��AK����+�~R�e�[�����n�����W�p�����5\���/���2.�U$�׸G���]�X��B}[/:�h@7�Ӵn� R�p�\��U�w�C��v((��t�׳�;��.���>���������^v��� �n\l�M�����nׅaP7"+����!^c��~��u��w��Y��M����e�J��A'�U�S�H�BR[��s���a���FJ$h�C���z?Fϥ��xS��ɾ<���$Dݖ��&�
��޴=�yy�=�+.q��?A�B;$t��}�V�uw��D#��<`�/Ń�b�-l�lmqQ��X]8�;T���0��AJ���G]\v��h[�K$�x�kz��^�k��P�����2��w�ڽ�_߾�� �u�&$X�qs�r��'
���?h=�m���u^>�_H�[|�v���&S|��^��>8�͡AM�;�Dhq��M�Vx-*�^ց�N�~�q��H�UN;���5\�}� �����ݏ��}H�w�НG�=���p��Н41w�#��q)���%en�zt�ā�Ns��Z�T���z����:����{��w�No�c�Q�5I�,T�F	u}�D4�@�X�6�z���0� ��!�� �s������h�{R��n
�O妍O����js'��Z�|ܰ��(H���Ԩ��2��k�ѧ�iE��2G����-����x�?���7��y�ﵗ`��rG�9�#t-�~�wP��p�Ƶ�;8�s(L��������5�!"Yǎ����L�x&$Q_�@B9J�hr�es�I���d�����Zp��y�S3�\H���r\��[��	ʞl��O�to�X܊�FΐM%Q�c�<@�e�)���>�Qk���J�
��@?j�pnyG�#~7���Us�(��j9���oT�����[H�#���/���U<@["�����W]up�{�׿ԟ�A�Qfi�K�_3��?uir��iK�5�U�<X�Yۜl�dr+c��%���������ݠ �"4i�^���~l�K��\���~�#$�����n��l6��n 5���z�����1?�-���q�h":_��Q������M@	����|�1�
:����n��Dj���Mlɶ�f���py� .��.Ƹ���N��,[p���~�|�;�] �P����:U�m���&��v7(�#�B��琻���b�"j4����6������q�9Uזg�_Y\�pyu�~'��o�@}3ԋ�B�ڰ�ߣx�f�}Ŗy�4^�!���R1b;��_L�K�Hx�,]r'�����Ac�T�-c�Xi�m8����w�F�;��&�L�{AO.���UؑK`��:���Dq�ł׏�B��h�{Y����vp������\�w��߷�ۑQ�ˇ�Ck���=y��:�wᛞ�ϵ"�?���,��!Y���q�d̮ǟ��S�n��c����F���e`�@��<}���ND��a�{�q����[.��n��Jz���u��$<�Zb�[��l^'%s+k�����v������}WNy��W��/+�r;��V��Wi����Y�F��پ�󲺊���������=���O��w��HB'|�G���߅���~m;�����PX�d����Ń�ڡX޲�=R�&��(]��еW���K6�KLJL�=nM�y��ꂆPb�c��>b"l��*��)��ޟ:`��6�a���
�#�A@�l�d���[�*J)	�&�Y�4U�������A��H�0J�_��K�a�d~����g�:����VF��hӄ�JU-�@�~ַQqx5ٯ���Z���^����������HG���hli�~��m/]z��o�	��ٿ�����ݖ��+W�c?�ɗ�{�꿼z�$�a�D�ۊ\���=���:,ֹ:��!�� ���dǡ�Y�f��F	�A¡(o=�+5K�0>�+[��*�'��"IV��K0���4b�>����R��R�BIh�i�D�I��`$T�2��p�Bi�X��}�2O��b�\���d��B�H���ˉ�(u�'i$V4Gc�3�EB�#����;���v�:i�o��^Ajg�8�:���7^�]?��uj����Q
�uj���9o���~t,m9!Z�v/g넚�7p�#gҺ����vB�r��W�n���.�;6*���oO���z���owpR�~�a������Ο��G�k}/��9o���_Ev�P�n!+�t���aN�woK��q�\�DbC'������͐�7fb/�8
U2���w�d�G4j�G�J֕�E���Yy���%�4��/�p~���I�h��_F%j�ʰ�%)׭J'�`�K��?N>b2�ѧ�6��L�d��߬���@��+�t�R�g`s�;��	w,�z�3��W�
���`5|#�.~%\\���
��>4�^�?��8�Q����<�O$��Y�͙���'���2�lOg[Z��ru��%U����"�ٲҿ�	���F�����gPK�̽Ρ'���.o9�k�VC�5�T�E�	:��)�V�~�R# �Q(!d�u�H�+����� �����M�x}h���������U��.�on��-
��,W��/����?��
\{�X<|�¦�s�>?h�s�={_E�z����ۗ�f�u<g|�RF��e{��1��������֕����Cv�$��H!��Ą#I��=>A��k�xf�'j%�T�eXw`�&�Hڿ2T�I��Gz����m��%>ߴq�*�K��5͠�1��F-5�*�!*�\8�2��@zcw�M�7�|J�+�DCjC�6�ɐ6'h~o�t�z�h7�]}m�߻֋���$}���,shW�w#�k{p.��:}�����/����+��e��[�%��
�~x	"��;���������;o���Ґ�7��sz�܍js�2Z��'�6��u����G��?��~�nG�P����r��2��8ԱC��lJRd]��N|��4�r�* �I�t�����6��dH\���k��l*��ȵ�垄F�)_V��:���b����J+dU.UG�=��O���!X�t����K$��ߝ�KnO���m_&$�o���l뿎g�J�!Oȣ?�����;��	?��q�~#���W��r�8�%H7�L��O��~.��n�f-���dِ�HIEÄ�7�5�3��57�F$�U6�&Lc?'*�;&⹲֖�
%�!@Bo�^�c�t���I?�	l8Q�`����T�R���)n[hK�,R?�0�S��-�s�sp��\::8��^���ֿ�@|�^���f����=���܃�!/�5,P8����gΜ�����>��0�k�������j�.s~)��K���%�N�ڲW���TJ�n\`h�M*��U�'�Q�"HV6?��9.��a��!<�÷m��?��Ko|�k)�T���1�_�����.n��a�1<���~�$�\��uX,Z)���$���8�N|����u�Է�ݓ"JCZ:ɭ��J�c��IR@���Gi����q��km����3H�<�+E('�-e�e�����H>�(P^�^GfPJ���_+�#��i$Q�t�fGTy�8�8���"��b�:�T.7������t��>Ń~���쳴U�ͻ�����ڍ���t��:}	�"n�� id\�H��Y��u�41���btO">Y|����ӕ���!
��՗��jާZodͷ��fj�X7�ȷ${9�PʤB�2��ي:�5�*����w�"m{�!�Ԗ�X���$-O���s�5�Ggw���}$�g�����h��[��~��k/�CIM���
.�}8>Xܩ.@ǿ:�}���{~��Ǐ^����w��/��������'и�h���3�$�����Z-������D1$�b�b�Z?*\TRB@y,�X�r�k���ٚ���+�d��/�v)�L^+�8���<bd��h�`��`Wy��r��1h5J�<k�]F���,L|Z8�]z��?�FJ��f��|9�����Z��̣�l��yl\�;�"t�O=���<�?��|��+9�r����ٕ����>R��'q��萺�����4,�Щ�$��H	]\�b���&�b�2�hY�v�K�����3ژړ�T��5ר���j�r��~♭�ƭ�7{��ó8�x�")d������$C�tc�8��ษ��98���s~���K��w��/��ڷ��wp�O���1�;w��ӟ���������1ʧgК|��}����z���Ç�j�4��g}�m/V�_"�י�Y�Չf$SZ����X���)oП�2�M4`'�(\6f8LYf2����ÛF�s),E͠�w����DI��F9Zd����
���r���Bo�3וe���;d�kh��j����WQ���ܝ\�t�)��k�|
�Y:ᡇ�m,m��~�����{��p?�,����a{W�ǐ�?�W��H��"��C�z�O\DH�B�9Qt�i����Y�Kq2}|��5sR3�?��Y�U�mm=ZWK<;8�jNT�4�Hڌ�,t�~�עl�m7�*�s�,Z���耖,�1�%F��`}p��ѽ/�q���_;sp�6�o�&��;����p8���������y�m��}���s��j��'oý��O�����w�ǡ���L�|h�Ȣ��{�d-o�zhTlHy!֜u������B�y�|#�2�����[ו���9��N�0-����9j��t�Ci1�ڕc�A��$�)ɓ�Q�	ߏ2\���'U����_����0��LP����;ys�{N�zl~�l	�0uURS���z��2R�ej,������_�{C�°[��{���Cx���^܄тG�χ1!o���?�c������\*rB�9k���E)��[[�ɐ�=�h;�4��l����i_iz��[TR��N�� ����j��q��qLK�:����"�`��{��їV���}᥯\=\���K?��t�; ��'�����|�$��}�8��<t/T����rN'G9ԗ���c�2<����!�=(��#C@�-�|[�����]�=2��c	&��A�zγu��ReI��)�|�&"�[Ge��X�6�Mr�Ř 
06�	eh��:�UT��>�K&����->�?�5�
�ĺz�m|��R׿c�^W�Js��;��g�Mf�>�0�����Ԕ���K�C��}}��.�[H�oqV�嫰~���C�o��S���U��R�8��de�zu��zf��7�7�7��q�-mkf[���1�1p���)Y���#nY�֋o�bt}r'�m��]�!"�䦪B��h���n����i�r������4�����/_���g�y�_<��'O?���}�U���08�;��G��dI_y�۰���&��d�7��_|��?�{��Vi�[P#�&��������Q�܅�~�:,�a8LCZ#!���u��9СT�ID�Ȃ�
r�'9^8�$,iD�!C��F5�q%{��Y�Xq����ax�o��ȚjJ)��O��N��ŚH�*�N}
�B��F�����Fc�*�G�]l���K''�|��q_ ��ݯ�Ï���o��?�y�3��"�)��'���{��p8�=��V�M�"8f�m	��p8�9�	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8���o��<"�*}    IEND�B`�PK
     Ps�[d��   �   /   images/d3b73945-fe79-451b-b309-b64aab767520.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     Ps�[Vm�80 80 /   images/9ce856c6-be81-4769-87b3-53be9928d02a.png�PNG

   IHDR  �  A   s���   	pHYs  A  Ak!T�   tEXtSoftware www.inkscape.org��<  ��IDATx���	|e��_vs���@iI�3��5�X����(�"ʩ�R��'(�x������(7価 ��(Vc��&)G�+M�l��/ݩ�4��f�wf���3��M�����;�3�;�[:00 DDDDDDDT\�BDDDDDDDEǀNDDDDDDd t"""""""0���������� �DDDDDDD`@'""""""2 :��)+S�L�v����/))���X,[�-��?'DDDDDd���QW_��r<\��UX��eq__�;�l�͢��
:k�ĉc***����Xf`�K���8��8��o;k"""""2ˆu�����tuu�ٶ݊��[��簞��^�`/�w�I���8��e����}���������1䀏a}�x˲�a�������sZZZڅ򂡋ֳm;�՗���e��l�p~8և����!���>�������ΕB9ÀN���d2y.��0 DDDDDD�@8��+**~�,q+�/�F���F�ݧ�Kjjj����z�8Qt��3�>ݶ퇓��O�īBYc@�!<_�,���Q������FF{�j���5�CP?A���1��H8�200�Gl~^������rK���
����9���g���N�Z����l^�e��O�oVTT|ɲ�����Bia@�8۶w��N,"""""��	���܈L�5k֜�t��B�ŀ�a�e���/ج"""""��8nԨQ�'����ׅ�Ā�A'NSQQ�W�����������G>yɶ��b�+�6��c��p�����I�������Q���,�@H?g``�_�C�=���v2v�Ǳ9E�������s�[�Ue��q��B�1�{D8nĎ�6'
�َ��Ȕ)S�X�hQ�� t@8���al�""""""w�Too�3���D"�����|*��}�pNDDDTp�@@���&�u�mo�x�O��D�k2�|��������U�s�.
�l���|k!"""��C��RRR��ߕN�O�B�p?K���ƿosx�6c�����q���O|�ݥηE8����P�����?�V6���{}�qoo�`e���ȱv�Z���Q�FIii������"� rq�����P˲���|�?`t�N[���nl� Di��y���M��p���������n�s2�ާ�l�u�e8FVc{%֫�W��{�߮�z��,���}�7��J��ƿ�q�;v�{���F����ܛ�sGṣ���K��c�g+����;��ߴ�1Z����x,~>F���>�R���]K������e4O�y���|�5�6��#��� �Z_qi��D۶`}���a�����
"�H6!3�@���e�);�2���ë�/�;t�>��l'��Xn���?_VVV������e�|s�}��H��oTUU�G�_ZZ�->������zBj{[���mɺYLʄ�ȴ�����=z��t�6S�_�j�ōP��ڲ����ć�]&;�y�qZ���\�ز��������i����,hӅ��Dj�m�mQ��P�oO$��>ǟ~~KS˰P~�L�4i��k�v|���5,,��B�YK-�m�(ϴ�r���RVV��t*87��2�۷۶�[,{_|��E�kPѸ	����T�F��VsJS;��X���.���kjjښ���
D�~��Բ`��W__��5kj�&!�O��&�"��}����
Q�.�AI/���lM�B�@8w�����~���]�*����v��K�"FTH��t�m�~��wP�� �|1��Ŝ�}����c����uuu[���=6�l��z{T�S���i@_�j�`��ޟN�/
�P�n��)ؼ^|��%����$&>ÐN�����ؒΏ􊌆�P!x����o�B�N*БO���%�|��ɓ�C9����Xvďv���I�k�hz~q�M�-u�k^���� ��秮��.
�*Q�_��!�
AOjzr#_�{��@�����X�USS�_vG��,^�xp0?,����<n��i*6?��IC�`x��NqZ��=��W�y������,�	�.��{����)_��\��s 8Oґ��-��G~娆�18C��ڧ�!���1�b�����#]j�|���@����4�p̜����h4:O|��puuu:�����)��pR�m��0�'�y�d����z![ũ�P�l�J����ik;�����`h���S���X'� r:sQ�|T�	����������8ysD��t�N��z�Ԁm�n�2������|�DFK��?�ZM�2e�o3�/�~�;��B��LǦ��q�ʄ3ی��iYց�x�)�8t��`4�
}C:��Os��(_�w6��x�4N��	�G,Z���'R� ���7��}�4`ߟ��GiK��oؚN�к�ޞ�7(�:�s�b
��tʔ�R8#��K�X�����X,��_�J�{���"'NS^^>��~x�)Y��^)�Nk:�c���k8O9���=�����a膪������!�ҥ�����jn�B�\���g[[[[��>���s%VsS�L�:���>�о7��B��\L��t��B��y8���|�c@7T2�<Ax�C:m�r���	���D�4���b�"��u^���_��Zj��4l� Y��>Fȕ6��MG{'b8_�P(N$Q�(ts�$��t����L�R�}��)�����I�m!��J�2/���������sO�����w~�����f���Ӛ�������C8fb}�x��,��;�t��9]�9�(�^N�VlzU�5,O"<Y]]�,�;#*��1���~���^VV�G а�K��+hǹ7���Uw�a8�(��Ot*$�<Oὲ�s�13������I�ӧE;ʭGQ~=���	��Nd��=��w�4iR��Cp�~�Jk4=�ioA���z�0�i�p8<=��b@7N��e�!ݿ8}Z�i+�+������D"�`�>�k�c�J�P(T�s��@���nI�uڢ���q:6o�E8�A�>��s˟���p��ߠ�u1�S��$�qL�BYcH���T7���� �sR�@��%��X=�Zt&��([�q~(�wl���DÕvyשش�Cޓm8�@��AhO��f ��G�NZo�[���?+ŀn�`0��� �F�!��j^�by����]�t�
!"O�D"���B۶���(*��?��m!dWNk:�c�l¹~��Q��b�}��^��ߧ�������p8\���t��/�����F9�J���#`1�{�O�/|��8f����D"����u�&����b�c5[����-Q�jH�"ʅC�Ӹ��*��M�:��ݲ	�#�]���t]��Ч��U<�� ��X��)��z��W�6�7�j��+x�ޣ����V�`�/h���~r*����(,[��h�v�q�n���ekl��u�m��e@9���5����o�+v7�5���'4M�{X��ywj�=��{xK��.�ﵷ�������XݮK]]�(����wp>�c�m'T4z�ZϏZ�ak�;e��{���r1�֑u����:��|Z�)��������`�I(vZ��*��`�M.0�{��n��k�EX��ػ+�����&��q��#�9��Tʺ�=�	^�M7\hy��u�\]W��qއ�m�^����w�bݒZ���Z��[�D��z����h��ǹ�e��W�9)�g*0���̙��)r�Lù����A����.
�b@7�'� �c$W�������0��Ő�nz�FO\n�?�PQ,�᳼��5!J�^\�m�����L��j��t�v�7
�[k���^˃0�5֓������@�k��5�o��obY����߱X���cV��-����������3p*�<�M8׋0��)�!]_�%ӻM�2'u��3��m7Wj4Xk8��� �]m����OX�ߗ3��2, t�ikk{�+�������	�pUa����*���Zk��	��n8�r�K����*�����>��������㳝��q��k��2��(�]���7�s������x�t�8ӱi�'��è8���ܹg<��w�{s�9�Ǐa�P<�G�Ap��^\J���2�;r��FOVZ2��O+����s��l�_�C�������f^������W竮�qR�uH[�u�e0�c����y�����F[��4�>5u��Cp}�_���Xkh݋�=�7=�Kmm���G�o=	�^�O�y�G5l�5�<N�4S�P��+W��a?�A�)�v�_����w�g�U+�S j�Cf��iYӦ�gp,ތ
�=�-�r��S���X�B�`��w:Y�S����T;��oWѺ����v����w׏�������g0��D�-����f邿��I��8,�WNK(�c3��E�i|�p^���SJ߫�R�S��R/.T��h-����Uk�S02��E�^<1�d` ���Hohiiir5˲G�����+/Zy�ܲ�.�����b���x��}/VVV��JO�X,֌���~
�>��x2��/	�X�ݧV�^��5��'�p�
=���>��d(?\�y(��I�����e��B�ۤ'=��
C�Y�� i��'����S���C��!��:������Z��7�'��,//��#�ʭ�u�8q�9�����Щx���|���UgB�Ǝ|2FCI8׋���Μi�M��Ὅ�a@7D8���u��BB�\ޓ̐n��H�4,z6ʋ�%�w�<��-eee�`��$цth���b?�F��UTN���^YY���[�;;;�f�u�.�X��u�O?k�G�Z�j�ᣐ�8����sG.�;ϔ�s�:��a@7�1n��Y��'=�68�
�ӧ�mN�7c}u<_ �i���^��;?L��6���Xסּe�j�7�y!�����7u���/_~����� a�zN�X/Z�� ��a��%X��H���4|.�����kA׮�.,�՝�i�eH/�hW;ڬ��܀��� K���iK":e�r��t�����.\�'�;t�m[�R:����PN8�霎-8�m~�se@����s��L1Z��yA�!�0�B�^E��iC�
�|NI$/�Ҹq����z�����
F�AX���}%B��8�>��1�����+�V�e˖���l<��Јq:���e8/V�w��t��.��V�<���0�痶��j�<Z��j��yo9i�!����<G�rC>��.�[�Ձ���9�� ����V�9���	�o`9A��9O#�LǦu�b���5�n9/FO[}�.���i	Љ6�{l5� *�O���B�#��6�}�F���M���X-��a]R#�WWW?���d�ȝ�X�_X���~��T�,,uBYs�c���8[��ѭ]�}�B6�i�m�]������6��{�6I�܉�h4�/!���<t��I��K�K׏��ѡ����
M$Q1X���2��kjj���-<��pP��i�7،���g�G_��#�>�W1�S֊�奐��!}d�Ĥ��,�?�ȫ����f7vJ�����v�?T�a}��k]��	S�_O�BzR�����~�����D��5�ӱ�/ߍ���7��LݖL���P�)kz���M��Czv�K�8�V��^������٦Vl�L(_o�qt��k�$*��X�@X?����Oc�|?{(b�H$�&VgTWW���Wo�e[��9ӱi]ȍSJ!zj��ߣ������ߢ���9����}N�-9��dC�B��BcHO��GZ����#X.��b�
Q��h������Ac;���D[صu]��nb}���4�,Y���B�Х����<�"���c+d��-
y;������bI���ѣ���D�ǀ�szp����n6�J���)=��u@3�O����.K��è����&!��`q�d�uA��C������!���;;;W�!��j�����/555_@�G��K(#έkZ�tl�z��B����;p���%}���h8���S������r�`�4\i(ӂ�\���bH�4-ȝ���i��o8~����*D9�c�>����"����X}U�����p8�2�_h�>�� ��t�����M���ʥM�}Nk���~�M��:>���s�5��E�������Ӗt=��`�4�k���[��J�v�1�;C����|�r,7������%B�c�X�۲����=E�ܣ�����u��ض�ol?��L�
�D�����|���r�p���8��ڋR��ck���\�4gB�^z�$W�׹ؐ�p���y��i�[�3	�z ��*�ô�Y��u8}��c���������UB�G��܊��)B�^����,�z��am]G(x��ehj>��jjj~�c�G�>NXGN��4��-�;�;�:���K6�p��@����
,�9>�!Ε�LC�3G�Cz����!�ӧI'��a��2uO#Q�E�ѧj�	����r"�'���u#�?����z/�zg��T[[�[X�TWWw!�q:���)چ�qk�י�7�Ы߁.�],��̹Mթ��3��yv��#���i�uW��g�h�~�>o5�ptIii�5�*�
M�#�ߎ��\!�ђ�s��p8���9�SܓH$b�xC�qD��c�2s�������!8��h���tl&��i=M��k]ܙs\��t��z>ourD��<k�I��gҝ�6z�N��dspj�����k�SH�6����ZA��,�X���f,��e��[��m��Q���{R������[UUU�B�滺-lQ�,g:6mI�z����7���b�td�yn0��feҕsOG�t��l�뻆q�>���s�Tz�[W>q���q\���l� �[�
�#�,��T!�>�44�nD�������I�V0�n��B��������X8�f8�4{�5�M�X��K8�ވ1�Ӱ���ٴ�j��{=p�Bz�6nNW|��t�o3ȓ��\��Dƞ�QQ������e�(?/"���囨3|Ӳ�V�kX�F��(P%en�3kjj.�?�uSʱ.=g*0�ic�[1���<�X�PZ�.�#��A<��鸼ҝy0���>m%�?����zѢE]b�I�&U��s	N��ض==5�0�r�-� ���o�"���I�EYxo!�z[[[�3Q��Σ�5��l��,�aݍӱ1�O{�j8��a@��iHׂՇ-�is{H��i����y�����x<��
�^)*��`��X�L������ݛ��|98�i��s����
���z<
���B������ά���#��(��$�[8!]ot���i8מ��[�8B�N�dH�[C�3MJ>G�4�����<�%�`�px?T<�,��xZ{{��0�.��r�0�m�6��������H��X�rz��K����G8����LnMg8�^ha8�tʘS����5#n�>�>m ����F�����؜)�L��-?�m�vu�����;Q�\!���hc�sP�x<���O#�%�.�� �Nk����Ŵ���p><��2j'4�tʊN��!]�+�MsCH׫��H�>�
���!�?'�;�Ptvu�#��퇱�%!���0�=��{t;��:��EX��>�iM���Iӱ1�O[�+*��K�m�)kΈ��C39��l��(����M���^���'l~2������h7wt�����8���Y�P��@ �l��8���tl�tl��Ӌ)�yǀN#�!�iI��<�iѐ���I]���6υ>�rIii�---F_IB0��_c9]��ξ9���/اAeRg`��h�x$yS�H$Vcu�eYע����;ʼ~�E�L�V��t���9cP�1�ӈ9]]ؒ>4';��IP�'L�68 >����;�`����B�����K������p8|�����BD�11Xj��o���!�^8��8��ν�@��|xl9/,t�	�%��Њҵ%�'�=��;�X�Yg��Ζe��{��%�uvv� �_	y*��cŀN$�ǃ1��7'�H������eԛ.�v��z�W�Z5XW*�tlzA�u���`n�8~��N9�iee�`A���V������j����Pщ�o=+�?(��B��@@��ޓ�ӳ����gWw�þ�$*��Cd��������{�ԩS����:K��7�i_�=�ӵ���p^�S:]�Ή�oh��dS��B~h5�Ae�����ϟ�p~��ج�ӯ�3��������m:U8����5�����u$�+&M�tg__߯P7�1�)� Z_�u�W�z:6���ic�3 4:��[l��`�ǖ�M����~i5דǘ1c��1��Ϸ���b ۶CX]�p^���weWwHusg@'_sK������.�ꫡP�O8G\��݅i=�@.Wu&���1�:�Ӫɐ>�|�t�⬭�^����1v�؍Oc�������b���Ʋ���s�y��B�^����F��<+�?gYV����Iӫ�D"�x���d/��X�?/4H�L�tl#iMg8��X(���44~��7���eH��X[���Uzk�s=y�流A��i8��fC~}9����Lf���%�w�D@���w�ȟ�O�0�e�=���=y���p>��O�,���"��u�l�f8�<�c��v�:商t������J.B�3
��/����|�Ǿ���ojjz[�(5܅X�'ŝ�v��w��Lȳ��ݎc����)/���x���N������3�w���{��@��|��si��t�;=蝖t��MIH���|/ғŖ[n�����X�Ķ�ϧ�!�� p��EMM̓mmmo	yR4���N��"�A�	�0���o�Ͳ�s������{�ʕi�+�p�yl97:C��2�z��.�^�<���.N�r�����ܹsڭ{���ۭ]�V[�O�T��7|����N���n����x����Iݦt�m�wa���Gr�j:6���c87:�ҵ+��G�V:!]��;�y�^7n\�'��+V��CR �e��[[ͷ3��x6��d2y�t�w���"�X,�����t�z������ش5}��͜��hӜz�ގJfa@��ڰ%�!}�4��紩.��Z�'����IB�Mj�t�`qy赵�����u���7x�G"��B���0ض�#�O"�@����P"�x����9DO"7�x��#����N}i��o�ַ���pn&t*
-�>��H8���t�O��'T��<'T��e�]&.X��S� �_��P��B�aTX�ы	��x�[,�B��誥�eVg��������B�u%m ��Ou��4�ex� :�sϋ^�dH�4'���`/_��U��F�����w�c:u�y��N�l����	y���P!���5�����s�s�H�����]:::t&D.���<&��p+Cq�@f87:�Ӓ�W<飜ڽzX��y�b�U�a@שӂ���^�!ŝ:mD�/]��F�mB���/ض=�3�����b1�`�i�.���0�׋;/ S��>�LMG�ÀNE��z(��M�b8�@���G2�{>9}�����{e�/�p�7��u�.���
�,��"������ۇ�����eY���ϰ��$K���s�p��d�t�ЮU�j^��Dj�������v!��㡗FR�B8>.��&�)���s���.vs'�{T�#RS�]���(γ7b{!_Ӗs�{�{0��14�khs�#o)P��Ǝkll<���)�IP`��{�6�ŃP��r���O/^��C�3ZZZZm�~U�ŕ��9��WhH�x|�T���tޛ�SN�vrt2��ҽ��9�Ǐ�B�ݷ��z����9�'8����Z�����8��y
���q�1����{{��t۶���4!��9��݉���!][ҝQ����C��X,vgCC���^耮���V@�ßE8���k�������h4z��g�{���/"�b@� ��o����f͚�d��g�tJ�a8w7t2����!]Gx'�z�W��xBTTT����{%6�*���tcc㔦��EC�T\�ľv6O�ݻ;00�׺�����%@e�ٶ�7���yϚd2���477k�ǏP6�+�.ZLȓtz��NH9ƀN��F1���N{�#�?l0�/�Ѝ�|;6�^�����d,n�����x�:��-�T�v�Zmm=[�K�t�g�D���:�X�������E�3�<E��ݏ���!�iI��\��2��Cރ��z|�����c�9�gw�yg��)S�����T|�j�1|/g���ۢ��sB��J&�?"�a��jnn^����Ok/*)|�6��s�`@'��}4:�{ww�����ɕ�ƍ����O�$oll,F�[kѢEa��>�m���^sKHPI����n���vY�H$�eYo���|B���=G����P�@ 0?-�Z��N��v��n���OƉ��t�?�x����O������珲��;}��k׮=���B���I^�H�XʙD"�y� ˲���ګ�ӱ��s�����+++C:������X��p�n���+������fA/����~�|w��IB��J�y�P�T�^������!��K�sEmm���d�Vlo/�
��ĀN�[�W���0E�ݠ�C���@p�x���khhxa�KR +W��}���|X��@�j|7{��r�x<����w���y �&�<�D"�'N�؀Ч��� d4���P����\GC:[ҋ��[X���l_C��*����_���d�ڵBi�
��������X�"�[��?�W˳��ΕXʹ,�q�����B�a8�6tr%�%�!���	���XlD�L�<��ŋ�$�S�龱b�
�Y�w������#��b!W�wy7�t�'8�e�����8�O&�w��B������I��o�\�iI���ay���o �_�����o��$�P���˗KOO�P�*�9^�pw� .W�F�M�m녖�B�n��^`�H��(?��,�**�vXù������������(/���h��7r�������$�-{9��|͚5����r�P(4뛄��,�"����^�R=�eYVS������p�������\�	�ڒ�`�[������t���~��^{�����yl�;���F^朆/�P!�}UU�c���B����n|���Z�_�F�	�����7�B�y�s��éBÖs�a@'Op
/mAՁ�h����'�K��K��w7�����;إ��{^�/++��p4_WK$/[��fX�\(�L�{�P��m�����¹����F(���:y�b��qk#������������  ^��-�y~j�4�A�_Ǉ��;����B����R}��Rr�������~*ʔ��'����I��/��)NaƐ��G���p�~!~قV566���e�<����tM��|w�	���V*�d2� *y��FK��+BFAP������<��)�щ�ܟ��sҳ�MЗ"����mA?4�|�GxH;�s����5�W�Xת��~���c6�"�9�a��`�@�h�9�-����ގ���cul%]�?1��'9���9��k%*?_E8�S�_��+������6?�����\�5�q�(α,��B��@���Դ6?�������s�-Y�d)�\���K<��Ј83��:y�3p�ڵk�6i����U�7��p=NF���z�eٲe�Q\|G�4�	����b@'7Y[VV����P�hK�y�m�t��`�ʘ��V�sb@'���/���-����c�XA�7�T�f���.�e���]��;utt|�˄�H�҂��~r��[ZZ�	���Z��&�JY+�6�s�O��Z����N�E�f���sRW��^�hhhx'�Ý���ڥ]�72�O������*�*z1ζ����� �	���2�[�^]]=����.aY��s�:�FEE�`K�ϻ�w�pj4�C���3е��|0��8[���և���p���L���������}�������际��$�!����s�1���hww�ç��K��pn�t5cƌyhŊK�����圌�9˲����rT���)oQ 7X�H$�r���f�h�l��?���0s|�9��Nyy���g!���������"b�����@ �noo/�Su����+�����������
������!�K͗Щ�8�c
�9m:���t���'Sv����3���s�
������$�U}}}���B������;W�x��GD���jjj�
���a��\YY��m�DCa@'��Ry<��1�rco���z����+�ntvjn��\C�CǊ�L�����B������m�{`�,��Һ��nI�9��kZPjKzww�xL��oE�ѫ�Px��900p�>r#��*,�M����ǟ�,�=l�"�Ly4u3y��$Q__�5k��Ù�3�{�-�t�=�> �t���K�ψ�&N�8a6B�QBn��m����r!W�q׏��Ql� D�>z��'酗����B�P���'t*5�sJ:�x'��Rӊ�D"�
'e{ԨQ��}�&�	�.>iҤ{Z[[[�\!5�:��/<,�Y:��O����9�e�q����S�j}�h8�K�R���+�Z����t>�'�P�{��uN����ǍN��y!W(++{��Y.Df�G$�@�����e�Pw�);=?��y��[�ZI�9�D)k׮um8G�}b���_nnn6vq۶OG8��0x�!������2ޢE���}=����,���#�x�����}�ɤ��_+�t�_G�a@'���.��D"�uS����B��eXW���X__�����Ct4wt2J0���>�D�=iҤ=���5�O�� �ɮ�9�;�d]��u�D��%�X�<1�ԩS�-˺���Aǒ΍�-!�������8��?�{_2q���***���ϊ���;��|O�f��.�o���Yb(�'Z���`!?�?˲n���/	-�,�m�Ml�(D�_ȷ:;;WN�:���˗߄}��(vu��0�����k�*,_F8TUWWW��C�ݗtn���4pnt��;z�:��B��p��^�IǇB���>K<�]�is�W����k��d2yh"���*O�J?6?&�W;�r��/d�@ �8�W�A&H����&�{(�t�޳mێ`��(vu��0��o��k{;NZ�C8_ �B8����69��ϡ��3T���b�N�G�r=�r�������p�`0�8\�zEgj�t�evu��xng'J�ۺ����"�|6�7��jjj>����pN��~�[��2VKK˚�tk����8�}D4�!�}�On^HdWw���K.�ڮ�8���b(˲vA8��
QJII�W�o\�ǟ2�'��΀N��5v��g�h��m�Y75�X�vu��1��︬k��d2��D"�
lW�T���>�ƕ����655�2�cX~+DE200��&DC��bφ��Sc�l#®�1t��um��f͚#�.]�B
�v�=u���ڱ����X_&d�h4�жm�c	Q�<���hX(�����/�'����;m�{������7jԨcc���WP��/))yX�ixb��ƙ��8�O��[�}��iC�,�D�U�O��3�������|�E]���n��7�Kp(���'��hxc8`��Rӭ�"D��ȳ�H�!Ʈ��*--��:ҙ����|����x�����|�-]��>�H$3c���W���'��86k�(M0�l���O���i�"6�PA����iH����ƍ;�'������`P��zk�ZHgWwR����е�F����}{���rKT��{��e�ƙ����Ӷm�1�BT@"
�Fv�9�k�3e���ҷ�f�������Ů�ĀN�璮���b�3|�b(T�u�Q��d7!��3�\a@��z����U�`�=��u�� ���e�t�ַ��y$���;1�����k;NBW#��mr8�{Z�u'6����q�Ҁ�BT8�����A�ԃN@}c�L��Őή���o�<����xo���������X*D#�����P�@�K���>򞞞���u��f̘Q�L&���i�����Őή��ŀN�ez�v����b��ٶ}��U�r�ƙ	���8�bsg!ʿ� �-����Q���ˮUUU �����,���k!]/ZhH=z���0��'��k��s~�.���_	Q�����qg��΀Ny���!ϛ2e�8�S-������Ɩ[n���結��.���/��ɓ��~]<?��n����-�(��JyPRR�	g|/sq�K�����B������Z�b�a�`����ޭ��wwwK2��q�����B:���:y��]�u*�X,v��©������f���3*�Ϣ�ԩ�B�?-�D�5!���tvl�D�F��ƴ���筶�j0L����}�ϓή��ÀN�bx���DN3=�WUUM,--}'ح�(�t��˱���ZZZ���C�E����=dڴi[!�z�ױLs~�bŊ!{3jc��u>�|А�y����_�-��ܵ��x<~ޛ�g����2���&	Q�2w�eY�8`�9𝼈������]�D���a/�OD���Un��&�k0���-��ҝ��!]/��Ѯ�nƮ����N�ap��GF�u���\utt\�է���8`�AP�}Q[(?b�x|��+��!���g���EV�\�V���f�%��,�����-�ڒ���ή����N�`p���Ώjnn6��mȶ�bu��3���Q�����J6u��򊊊�����(&?h�I&u�Czyy�䃆tg�87�tvu�~��	�vm'�/�b17��C�өQq]0iҤ�[[[�U<��eYK�9A�r������]�����X�2jԨS��������Li�	���VC�����_#bWw�c@'�3�k������Εb8��ۅ�6Sq��q���*TTں�������jokkc���>c{zz�J&�'�8(��kx�zY����d�رy�ƭ��5�/[�̵!�]ݽ��\�Ю틂��g[[[��UWWO(--}�[
Q��2xrmm�#��|��Jusg@�\�c�L&~�ӣ�3����c�m��{�GB�u˗/��W �n�:��t�bWwo�J�f`��6��>�n�8�-˺��Bd�@2����޼G����I�����1cF��c��5��;���]�zu��א���kW�|�n�ҵ�ޭ��ݻ�ɵ�ھ'�/D"����m_���Y!2˞�7��x�PѠb</hM���P�t���煊J�G�>}�8�u�#��d�t��V��\rF�3f��èQ�/dsϼ	�^��w��0��+ص}5
�C�����pX�d����eUUU���綶GiCY�ڲ����B�ؗ������U�،3l�S�ohh8����0����5�k�O�Kχ����������U�͝]ݽ��&��a]���#c��?�l���k��\VYY�����P� P�Gt�	��^x����ƍ;��3p<��/�vk�������!Z��烶���www�����0���ֵ]o�==�<!.P[[�5V�`��M]D��Ú�����"BŲ �qB4r��X~F� f̘�I���4<���6ҁ���4����0v��d�����iO'g
vu�trӺ����$��(.������"D����BE�-���r�^�K�\Y�����q����q{&�V�߫�&�A��\�9���rKii�����~˾�2���-��U��~-�����P��X}^���+�e]��#�*����D9���y�����D<��ue��C�XC�4ҷ�z둄tm��ɛ�L���w޹~l<>��Yl�".î����N�aX������G�����vے�cٓӮ^{{{�eY�����-7n�SB9��n����O��)�*5jݬ��w�����!�C&O}��d2yݫ���tS�aѢE](�E����E���;����ބ�r�[��B�p�n���Jn�;�ᣱ�S��R�,DY�>t�{�F�c�	����ӣ�~�P�/Ľ�C��e˖vw&�/�>x���755�5�_���������.O�����+Ե������X,V��R&L�0vԨQ:(��N0DB��7����577s��G�%�42��>ӧO���S���1����:z{1iu��o"����6A��d<�Z4]h۶�y��,/�����j�#2�k��(�?�x��q�lY�u��Q�ܭ�����'TP(���G#�AEE�cB�k��F������Ѳ�&����C��{0�A���gvͼy����c��#�����"���~�d4�����{9&��G\'���,D�3&X�u#����
�E:?0Q��fϗ�5@ 8坶܎5��vm7�\Ж���{o)ʫ�[ZZ���k#��	���a�[�"���n���hum�?���8�|��	�wl����XW��	Q�p��Mh�v�y���ʎF?�.����aX����ۄ���'C�Ё�D�\�6�ߵ,��G�����{1�����~I,�%.������&lf4�)��P;Ƕ�p<�W� ��hE��U.D�iGPzV�#tz��ӧ�����!.:�
=�Z�B�@�8O|�7r��8�$��c�,3�%��ݽ��Hum�7��fz2��KC���Xl+D�S�}�b��*�����F��1!�������{X}}}'444|�|�����zz��cA�{�����H$2?W/������>�ӯ�����N���H�tm'��ʩ��eY^�"��q�����_*��΀N�b�v����7n����.��sZ��O&�Oڶ}0��+�z�h4چ����u��-�%���}��8�tmoG�~xgg�k�F8}��	��i�R,�
Gr�,,���9Fn��n��NB8�n��cHC^���k+,��n��\�t�ׯ�5O��]⒋-���>�dC�����8*�H��%B������"�� QP��GBD��Q��Cٲh�����,8Fo��N���8����O�q��x��Z�74N���Z����_�sq�-����.���(&tmǉ��(|_����q���;'?����n�ŭ��Q���.>�L���P.���s�L�V-CNH���/��E�Z�B�����`Ww�`@'cҵ��h4���p��*C��RO���Q�:�;��M�҄��[�x�_�q����XiW��x>6��Z/3qZ�iH,�!]/O�8񄊊
e�� ���:����O�i�veY�P1���K(7~�J�=MMMk��&�L����҃s�l�c�9&��ں�N���G���.�ھ)9�:NQ]]�a}}}��%�簫�;��!#е=��8���7᧋��I}GG�)X_#�7�������+S:�5y�x���}�W�y
���'\2�Z&r�[ZZZ-��JII����\Ů��sŎD�f@��nT(�Z�d�Rq����2�s��o���E�P�D"��>���
�о+��&ڜg�4�������V�Xq�ۧG˖���`HG��\<��xCx���z��~�{qvu7:�	]�Q���
�k�"����`��QM0<�˅�i�0��0p>�I\N|�Qر9�6~me���>wM���q����۶w�����n6~+TT��ڮW;����"�p�|f�"���G����477/�(n!ZwYY��Ņ�M��U 8u����*>���U�V���<�#���c@C�'����\�T4tm&��@\���nN�׋�s�����>�_�Gr��ܳhѢ.q	���������?)~?-4hŊn�V-ҵ��������B�З��ι>VǮ��b@��(v�v��������4(��w��ȭ��Z��Cp|�;a?-]�t�PΡ�\�V��to�u�]C8��lhh8!�����������Ȗ�m��L,{e�/�H$���'����$��\��n&~TE��ޏ����%�"8y��ٞBD�2~ԨQz/��B9�xu�g9��e�����+ƍw86OB9��&-_�\|x�o��Գ�GHc�/�F�,��n��]��ÀNg@����\���4>�������'N�x��M+�S��hh���#����'#��i�6K{6����Om��ɚ��O����5�K$?DHo��~b8vu7:�@�Gm��U-l���ڥ}���?�p�E��'�S(��g�
m�l1�{�e���d�D�	�Eoc��ꪔuӐ�Մ`0��]�E"��#y!�`5y��c֮]�*ֈ����,����ܵ=�E�r��'�\�X�����������P诜=�P�'D��F<_P�7�ӣ�3P���[��RZ��y��g5���cg�"J&�skjj�kkk���/^�a۶�O�Y����T0E�ھ�񨴿/.�p�X!D��*T�O��
��a:E�]�~��3�pn?���}L�8	�z����]�`�����������a������������>���b� ���?ñ��9Щ ��~.���"(�wxE���bu5*V��8�؂NCX�}��B�Bgz4s���H,eB����` �5o޼�6����?`�T�a�}}}���Q�N<��eY�`�@1�����>D���߅��Jq�=Q�5<ae���X_+�(C�QQ�
>犦��D>(�/�6mZ=B�	�"����G�k��ѣo{���?2e8>�~�ЦhC��&L��H���[+Q~���ױl+�cW��c@��+r��8�3�e�yi�ܝ����=T.�sӘ.��H!!���������Q+V�8���`�@����ʿ9�d�����r�0�~���6g�ѣG?RUUup{{��l_$�%�O��Cb�����^|�WE�ڮ�G�5��P��3��Fb˲>���B�����ɱ8�?����05�hO�mؒ��$�\O� k֬�o��Η���Nߺ��f�sݻ��������577g]�E}��̏ή���O���]���s���ඊ9��ǜ+�䪋��_8�_;����iӶ
���u,ӄҥ=o�����k��֚�B������Bi�>��io��h�B-�ש��:���cOl�)�cW��a@���n���ڎ���сo��u��BD�p *����kB�����чpw�H_D�{{a}b0���J�th+����-]x��J��P&�D=�6�_�Gޟ�455������L&u~t��gW��a@��ЃZ���2=я�
g1ض}>���BD9�J�v%<Q(
2��h4ږ��w�u�Pii�L�s��k2�GKۛX�B������Et`8���ƗүҞ�� �D"�Q�;�7���ս8�iS^�k;
ͳ[ZZZ�Ejkk�y] D�kǆB�'��Ј��Zή��������9S�N-���8X[�Q��p�:hz��݁��&���G�b�=൮�3p^Y��O�}�X,v����/�cW��c�H9W̮�8�\�B�6q����-����=s.W��+�Rq�Ј�r��4C�)������vhll�8V��5�T�'
�kpz4ԧnY�`A֣�o���K{� 4"(�G�~7��!��@��,|�{a��i�ս��)��ܵ�������A�{�ꅈ�崺���ZZZ�V8y�tvE&��p����>cQ�?*�L���� �t-�2[��?�s�⩁h��	|���#mCH�3��㜴,
}-<.�O�Ʈ��O�r��]ۓ((���ٹR\$���BD�4��c��V~���-�ԍ�ມ�Q�GC�8��x<�.�i���5Wgp;v���Ν��.��n~��5F(W��nB]nY4}<�H$O��W�{���]���r��]��2�ω�TUUM,--��Q���>"lA'�-�h4����k����/c��?,;qI��\�z�/��RG��eY�aB�����
�>���j6/PQQq����YƮ�ÀN9Q��o�w��N�%8Y���	p8��F����L&W�������Kj�>}��'t�#�c��G+J�dz�l466��;�R(_��;}���vo�=�'777����x����]���.�D����s���-�m�l|^�
*?ڊ�U��p�8�{����a�g�x�J�|,7������/�_�_����}�;
�S��ǫ���\�d��L��`�o���K�p���4b��ڎ��"������|"^*DTP:��eY�߸�.����@@ȟ����>��A��̹S{���+��M �}�!���(#SJKKﮯ�����g�d��~�S�as_1���:�H���ϟ8q����v3C8��`+��
m4�N��[���c�O酙��ʩB�I�^�4>����������~Cx?W!��*�}���o�g~\��0�'�O�s��������?U�"vm_���MMMk�E:;;/�j�QQ���:*?:�qR(#+�RF��p.�Y	,7���_~��1�m�3Q�}F���
�t�3}n<�O8����p��?�5���k;
���:�"�e�B�BD�4�V��>&��������?Z�=��Ƽb�.���>rӔ)S���;�� (���r���qs�}	�3}n,�=��%l�!cW��a@��8e���H$�(.
�*Q�ծ�A!�b��0�g���m*��e��%>��f>�-,7&���^}�Ռ+ �p�P����(3�ҟ��y�c���x
��ׄ]�}��&e��]�{Q`}M/q�g=Qn/DTt(?���������)�6�-���^lV���Z��u���755=/���:�g�(>��n���c��3yb"�x��6#�cW��c@���k;�_��k��x�g��N���'��j0��_��g��s˂V�L�:����.��������{477/���x�2�������`��{蔑"wm�ז[ni����2e�8���'J"��,ӑr/(RW �Q��	�����P;��y��-�����V��� ؗ>�f���K�P��7
����nt�eW���H)b�v��~�{�Ez{{��*,Dd�l����҆��1�CEE��*��ط�bߞ��{�6C�eZ=V�	��H˲.��g�<)�H��/���s1���oJ^�"����x<���
�#�:Q��T�	zFP�Z-�>�������c\7����������-�>�S|Go�>;'�'i�Ѯ�����=#��=w�)-��ڎ�����{��Huu���W�̅������oG"��҂2m�
�����ţt����y��=��\l�>ʁB&��(���Y����V�O�ޣ�p���~��o�dW���Gi)b�v���uvv�A�f�d2�ӯl'Dd��(׎��*��hw!�3f�x�|,7��|�/��x�eY��.r���`pN(��H$���F��m�Zl�.�cW��c@�a�k;��ǟ��D"O`�Smmm����>�x!"�������4m9/++�X��p'��7o�k�Q�@�w������(�n�J��������j1���:mV�Gm_ .���W��O�:�{|����{N�gz$~�����x�Ͳ�]����t���<�z��d��c{6����7���O	ǻq������{f���E�u���6oñ����S��*b�v�s^kk������R[[�u2�<�g`i"*6��\�a� q�ݳ\�z��r��[��+�,������s���ӫjjj�er?z,�!]{e~AǮ��c@�!�k{
�Y�A���o����I�umU?�W'*{3�s��J��������p�s���8��cǎ��ܹs�Vi)�������[m�@��u޴o���?���>_Ʈ��c@�M*r���@ ��U���!����.���8�_��9,A!�B����y��m��^��x��Fn�k׮�~����Czk��
��N�/��;�>���-���b<�Wb8vu�?-ڤbvm��R�n�F���]&M�T��߯]nu�	��;=�Ї�
![�=���+p��g���+O���8,�m�:|������7�}��ŞM�9[m��o��������]�3ǀNQ̮�(�:���.K�w�.�Q��^���LD.wX(�6�H�+4$���J���z>�ݬ���[.\�)W�Ų��� �B^�r�ĉwNwZ������~��]�3ǀNR��zu�---˄�z�9eʔ������$|G{�Zy �9ѯ[н����۱��h�655�Kh=۶w��GB^SWQQ�]ֿ������eݏr�p1��g��}H�Gm�g,�M�#tj���r;&�I�֤�7o+D�+'�p�=����ۓ�<������堍�]�Ȯæ��hD�϶�.�L�O��A���4�y�]��ǀN�y�v������gX�H�M�Ϋ�����e�tm�	�Y!�T�vB�-vC@Ū�Ŵ��z�r+B�_^}�ՈАP>���ӳz�vu�[UU������yꄋ-˺e�b8vuO:2�k�5�h�I(m---k��U���3��u� D���X82�8͚��=�X]N��q��Y>o޼�xq~x555���y�䲲����~�O@���8�N�z����N��O�y���8�\$��x<��Ϋ���iww�������@a�:Q�N@%�G8~�B���3KyGFn�`�qο��_~O(-����ݘ)'�m���t{s�������]��9P���ݵ]/\����.4b����*1G�P(�����{Չ2BEx_�Ӟ��O؂��z^�Jr��w�njjzU(c(���Q�/4�]��f�t/#�ߍ��	<�3b8�����/44t�ӃD�d��UUUʹD"�U�(��&q�5o��0���k�x��l����͛�Z(+�Ph7��ٵ�f pk#���}B0�v2�\ .�w쉵y���_�l9O�.Gjͯ!Z�O�2^�hS�����f�ءp�5o�������mXn�����	|\e���ߜ�I�=EZ�fδi�V:���_��z�媨W���uAq��(^pd�ʾ��M�a�m�Y�$�t�6s��{�IIK����d�9������3əI��9�����@�����X�'3��*��Gŝ5���nݺ-���$¶m_��O\����tS"��UP1C��z?=�;_ۧ�����f����U���1�������d�Ymƌ׮^�z�?���t:}�n^&�C�����o�|7@�3�E@�dI;����(-3��n.5����H˲>��k���A@�2��	��Ƅ�.g&�+Q����boڴ�KPRzm>V�N����s?�p������g�����h4z���$p-:&��8.H�RO
&��6��%K�|��������^^*���q�.=&fm޼�[0�ۻ�	����|�{ˣ�Wccc���ͽ�L����8��vYL��fV��~.���G�D@�d��(�*� r�^.\�`������T��5������[��4A�6�L�^3f�(����zp��)S����v	�*�N�FWx��H���qf����==Ws�r):&��XV�z��XeJ4]��ͧ�L*��ƍ�N�@���T(������ޮ��5�L�7�ׯ�$���~H7�@?�3g��m۶��Y*�����/�������{���񸙅�[���?0��}E!�?���y|��s�����=w����f�7�V_����/���.���ox�yuuuf��o峳��Ķ�k����QQz�8-�O�P=4����,�r�6 �;�s��O�RPw�2�t:mf�=W0���B555�eI-Wd2��mذ�UPq�X,���˵:K��}EC��Ds>;�~��o���W!����J�Ry�?����ֶN7�,^�������k���{��]f�;�9t�>}�H_��rC6���%KnY�re^P�<:;;�WX�c3�����?
xη��]KI�n@e�Q1�@�[�`}T�زeK�nΌ�b�ttt�'7���x˫l�^�o���]fʔ)���q�7"�k׮��`�E�ѷ��k��.<�����|v�k�?�v����.A@GEhx�?�_'�m��f�)���_�}�p~�W��3+O렻��q?��Z�֯6��z��k=eT��ŋӿ�%jȓ�������ܤ���}O�}O�jX�
4�Qz2����r��OZ�h��3��)Z7�^ w��Ї��]dʔ)[-�2�|^�iӦ=�����jhh��n�	��Wڶm�G�2��̈́��H�B}�}V�
tT�]�dr��7Z[[[t�K��ooo�'d��=[ wza4�i#g���������^��SO̫���og���(��o~�lٲ���B(�Q&���V�
�e�������ܼS7��b��ttt�[�&��� �c���}@w'k�M�����T=�Ϋ���XC�(����n�#��$����[m���V�)�zt��-�x|���r��_c�6J^���/jy�>
��~���Su�����Aw}��O&�W�Rcc�"�q�$\11�]�d�%�7o��g�P(tF:���VT5:�)kY�i���f&(�϶���Z>%�B������F��%>��/�I�0龜�R�,��M���/Z=T��9����T�~7��[ZZvD��s��xAU#�����M<O"���n�4���B!���)s�Rڨ6���:�=�UO�W����kUJ�#�տ�Q������D~�T�����{nmm헅������{�1��[�n��鍍�g��i3[��O��T�w�b���n��+zu����T%۶�2��ẗ3Z��|v�����F��6��U�����e2��$@�ZZZzus�^h��`��wX�e��[!@�xAgg�1��M|�uЫ��}��si���h8�n���>���L��Z>;��֞�����^��E@G98�`�O�P��}�7���P��Z��:�(>�Bz���dg]]ݙ����se��� �g�W�S����lV��@�z����*�Qrf򓶶����܄rǙ��8�Y�ZX�	��=˖-�l�k�z�JY����Җ�"����V���L4lD�kg�R�'��?����oz�g�%��O�QRC3����(m�����m� �7�������^t�A�Z�ĥ��bfl�k��B�+��5����l�f���yZ�����Qj71s;�%�J��͉.<\����?�udQy~�Nz�f�_ՒT�@ `E"������j�>#�H�#��kjj~����E����QR����r�P��A����w�1=ꨔ��q���+^<cƌ��޽[PU��L&W������ͻ�+�5�?��ι^�_j�4AU!����J�R�P!���I�h�,ݞ��f�'ܣ�����6���*��׾vJ��zl���c�� �Wu1��Z���s�n� @����H$���t���j�.�t�ҏ��x�I7�נ�L� ���ʲ�����!}8c�s�X�:�&�fA����u�hBL=]~���䳳�?����zn���j�Q*�A~� �hXP_��@z� e� 3��g�4���x��p8|����[�+	�Uo[MM�OUc���qs�p�&�	��m�G���q�s���9�����Z�����1�Z�e��)@i�a����q13�Պ+ެ��5� 4�\C��i�RAU���k�zs�Vk�\s~��;��9�4�_�����*�Q
Mzl�uFcT�T*�J�rm8�O�?�/-�Dr��]�_��WG���/_���}��U�Q=�](�
�H��7ku� ��x۶�-�H�=��3�����0��*�1a�`�Y�V�T�yM,���������`��}��e˖��a�K�.��5kֻ�z����8Kjp,�����L:�/�}�.�P]N���|vL�ROF�ћ���W�;ʋ���j����R�*�v�Z�,�אrUOO�i��ڟa�W�cǎ�t{�T���:�p˲N�p�I}x��Z&��_�����kU�s�T�����[wj�}Q�ޢ���x��|v��ӂ�^蘨���0ܭ��y�n�n���uk֩}� E�ƹ�^u=��Ҡ�aޟ�r���6�;�N��^�{��`�͛7on8�C�Q�T�^�c�����@�>�u�IE@�D������Pni�w444�S��&�/�@ڐ9�onn���m�S4�Y[[��@���آ'�s~�J��I�׍C5�߭�Pݎ����u�׎3�Mt�`R�Q4m^��ֶ] ���˖-��������GZf�����3���J�P/�s�i�U�}��i�*�=��Ϻ���L�H$�=�Vi�e��Yi������~��ǟ��K����be�Q�+< w�ƹ,�.�N�T0r���е���1z�5C�џ9�������d������z=�̄p��=�η�L����Z��L:����5mmm[����6ݼM��I����`��n�@:�~���	�0����}pC2�t�~^�;&�=�1\F�!���=���8�E�e��iM:���9x�6�/[�x��g�Ï
0�Y������D_�h�| 'h�>|��zơ��}�u��Y�dɬ\8_!��9�H$�m�<8޾�Tj��{�>竂IA@G1����a[�l���I�X��[�70:�荍��r���l6�F�r]��}q�6������~�9\O�/ߐ}תq9�s^0��V����!�bp�9|�L"�!j���3�᧵Х���[?��05�f�ht����~X�+�טm��ߩ£�s&��p�*����,���M��hn��m���W�Gi�Q�muuu�GZZZv��H$r�6������P}�^F�ǯ���n``����9I�MB��ׅ*}�A6��jGG�A�����B8�w���M��ֽs��>)h � z`��Yd�W�d����/�jC�]�4d�z�m�G�y�c��}�p� ��[�9| >	.\8�q3[;�^��h4��x<�y������Q�G*���B�����c[�nݦ�r3��F����?�=��9s�L������G>���p
g��_T\.���s�9���w���䳳^�����E��"�#oz��5�H$��L�[�u�>\.�H�mۗhc�L���4(�^o���!��ŋ���N��\ ������Z�#mӧ���*��LXr���(į�~�T�ImH�:�|W��l�>����� }u��Ԝ.�����y�tz�V_&��՚�-t���v�ߣa��Z���b���cz�� �����h4z���E,* P�on޼�[P1Q˲�����@ p������ݶ7&�q~����Ul*����h��U�u��Q���{�,Y������� 
�`*��LP1����4|�m��Ǵ`0�ݞ6ގf��m��j��	*���|�����L�W x$1�4���F  ?��/�ax�444�8�s� ��h{勍���䖒��$��^!t��L����^�q}n4�_�Wk}� ��~�H$T�mۯ�pn&��+�?�J��f6�3��q֬?www�B8^*���qiȸP $��]�t�}}}�1t� �(��K��F�j�h9T �JCC�y�Tj�X;555��UJ��A��1�'��� knnީ���E�d��R�`�@`���"������5������w}�Vg���e}R��QƤ���q��������^�.�~8`b���.\�63�}� ��X��+m�^m��Tj�������wl��u`ȩ�X�wk׮k����-�H�.=���c��� �0���kll���isL/ 0�7Y����+���7[[[�
&L����B�8����eV��r�5�_�z�q�¨������ ?f�E���+��{�~�%( �|f�G3��{5X�(�L�L��AQ�w�yݜ+�F��oj���F͆B����i3qt��l���������F7j�
��@ `dӴ��D>���D��7%�Y��{eCCÛu{�X;�����1�R�'ʆ��Ѵ����- �"�߮�#-�2B�� ��0��i��w555�ټys�`L��
����Z�� �2f����/��^���ˈ����w�G �M*�J,]��������8�I �3��|N��D"_L&��(���wt��c>" ��۶_�H$�1�Nz�yP�{R�/�#2] �]sss�n>������{��X4�8��k���5��a���khh����vP3��k���x;j[�2��eA@�HN�RO
���>}����nڱc�d2�`l�@>Q�Gk =Y��7
d��������y� (�;����~c���t�#a�۲ �c$,�T��ŋo۲eK�C�������_ `�,˺޶�������յ[|*�.�pq�V_. ��s�t���vJ$)=���[%G@��������V�\���b������eϞ=� ��rrmm�.�X[[�}�3��><�m0Q�,Y��'�MF.�㎀^t@�[Y���L��`0�-s�����z��s�N�t yX�8�=�m�8�L��/����U��Yˡ�f|Z�?k'm�\oY��3]PRt����$ٰaCs,3�_G��uuu��]̐w�K�s?��#���/^��-[�t������@ `F�M %��f��lٲ󚚚F��.�J�m���!AI�1\�^�n �F/�������a9�C�L700  ��c�|�v���w��s�� �֠��8w��\iY����D"�# &M:��FC��Z�9�5���t3ܽ��C@^"�x^m������ϲ�WF���5��X���������:w̞=������*(:���R L�M�6��b�X���ߛ9s��}�w��t �0�4оv�ܹu�,�B�m�J���r{�o�����v0C�u��j����!�cȿ���j0�,˺�q�O����S�{7C�u�<���������w�����͛7oZ$�*��/ *B����=�ϕ�@��^Bt��/z����{����bOh��#}���۷3y�|�<�N?b�������E/^|���n�jL T�[�2�mmm���C*�Z�Dڵ�@Ptr�P5��%�l��Ѿofw�/���O  f)�ۣ��g���%��o]b����RPi�_����%m���V�((	:�m�T�U��^���t:m&Au�b3yܬY��I߻w� @j�A}�6�O&�ߪ���#�ȫ��Z�# &�G��Y�_��瑫�X%��o��C=���n��	c�ǯ̘1cp�8ӛ y:U��?����+Uƶ�����
�N �iJ04=�?m���$�Ո`��`x;P��qzq6�=A�0eʔ����q 
pB:��u�ҥ'477W�'|�͐�s�X`�i[俗-[v���}��g���^��Lfx����L�>��]�vm���|�g�8 Excoo�����{{GGG�d�C*����o�j��������|�4�_��0��>��_�T�իW�W�Xq�����3y�^�������~�<,��ڶ��D"����,]������R�~@ T�fɵQ���*�<��&���s��^ T-�q.֋b��0�����ˮ]����G  ���MC�[5����?X�!��N�]G�����h4zt<_3����o����	!����P(�Z T�u��=�bŊ����B�gB�̙3�K7A �`�1������T*��?pѢE��1b�D T5m��^�5c|�Z�����j����r���!S�N\����N�q�猻���q�x|m9���z~�Q�o�	 78A��%zn�<�7��qGoo���!(�Ǵ�~� �z}}}W��ՙ���|}����� O��F���!=���ܬ�<M ��YY��Z�2�7������q��?�/(ݿ��p�����Դ;��Y�/�5��@�LH�c�ǵ���+�k8���_i5( \E���;w�����v���uZ�@@������3��0w˲>>��`�w ����l�>&�H<:��-��}�|_ �լ����t�������m��șE��So�e�����b�'e�)��{�nٻw� �8ղ�����T��b_d޼y�4��%��- \�q��k{��&�ikk�n���ZeU�"�}J�����u��z��d��cB��3{ԙ�@�X�u����iH���h4� �e]c����R=�Y�w�������^$�?=�H$���d2�KC���D�m�����- 0���/n�m�چx6�'����͍Z��34�AF�7k���(t�f��
 �ٸqc*�ݮշ��5��@^��憆�cR�Ը��h8�n��2S x�;-Z�����r�7��?��o��BA��>�����+����l��14û	��tZ `��,�
=�O�E�.	���/��,i	 /�2��gu������,�A�����8�}��zzzn���ۦ�9�|]Ӌ>{�������`�D"f��5��Q����V?' ��S���;���c��3��Ћ@@��{�D� p������˗_��௔�����&��ܹ�|  0�������x��C_�3g��fH{IG� �Z�����t{������K�׫�:AA����v��4H�a�%�CfΜ9����# 0=�����d2y�����άs� �s;����U�m�oZ}�� t�q�6�j�<�H����	+��3�O�.�P������П�n�����Kz� Wx�Y�!�H<z�7���*���D@�=@ZS��S����w�n��3���2l��`f��˴�����-�9=�?:���J�/(�G����v�;���gZ������H}}=˰-p�?�\��d~�����X;�R�M�H���z�G��,���k�v�b�k���r�,�a ��z5K\�m��ZZZZ�y��Հ~w �� ot�p��W x���E���`6  |���-g%��T�O�v�]�!����zplL$� �X�~���˗o��J�<s?��nBz__߈�d�Y�~3  \o���C��O[ZZ:�}}����+�'ǹG x�:����L�W�g��=k�,�V����/��  �����זe���ֶ}�/f��۶ݢ�FA^���Z xN(�(�N���`�~f.������w��Q  �]B����~A*��[��^��ӂ���!S[[�F x�C=���b�������~衇&�m��_�b����	  �cn��e(�}KKKo9~��=����D���o޼�[ x�Y]/|����~������������  �b��~�J���m��?H��=������퀇���������3vh���z���� p�@ p&�9S������[�l�m�Y�K�"���=�������/_~�^t?_ɟk>׋��  T3G�-Z~���>��l6{��S�y �{_����>�uh�X@7˩�ܹ�T�  ��dƕ_��d~�����d�C,�Z�m�O�E@��۶m�% <mݺu��b�Z=�?o���º�  T�=Z��8��R�TB���A䅀�} ��X*����e��R��  &h��_k�U2�|F�H"�h�m{�V��D@��@ � �����+4<��պr��]�� @i�rn��0/����O0&��e2z��x���]�b���l���{��ah;  �ah��?��g3̝�>���W�}' *�q���@Yz&��  `�L�Ri��m�5�e	�F@�0s�
 _Y�~��˗/�k5Z��6C����  ���J������#�B���"��n�N����a��0���N,�T��+�����J__�  ��2��"m��<�J��Ŵ���m{�V��`Ttt��2��E�`�;Z-�82m01  �ե�Z�K$ϊw<,�1н�w֬Y��lذ�5�ݣ�7���̒j&� ��۬�Z��`�#��f	��нk}SSS� �%� ���&�M0g�s  ��,�|v2�4��x�S�p8�������]k�o��������|_?��ٽ{7� P-��u�������F"��@ p�`Dt��}� �x�'�]�����n39  ()3�˕�^����g4��Y�����Q�`����^ /֋���s  Jj���-�:���m��}to��ǟ ���#�<��6i���>����e�  (�u�l��T*�'�r����1
�7m��`�Kͽm�>��� �����nq�\��1�������v �,˺,���T���>���  (�������`Έ�$��gl�Nh�<݃� �������,_��&=/�G�ϡ� ��qya�-x��=��g&��M^��s  �����a��_^ �]m��ō���==�d�	��ŋ߶e˖����ݻW  ���/�`����I0"���'���p+W���b�˵�?c�gzΙ� �Quk�4
�����UP4�,#"�{O� �A2����`�[Zu��={�  x�Z~�8��T��f%�L&7G"3��t����f 8Ȇ�W�X�F�o���t��s  �3��d2�LZ�i{ım�t,�Zp ��Ѓ`D��\���:�� 0;�Zy�^3��<!(�=o��7� t�ѓ	�����5�p�\���u=oHoo�  �cf���:yYKK��`��нeg{{����ٶ�^�,��Z-S�=6������@`��K6������su�i��9�����R��ڣe��T����}��ߥ_K{����_ۡ_�{<��e0ܡ�&k�����ݖe9����P(��w��ئM���b��Z���p��_ �g��]w���=�L>(�4n��[�����M��m���X/=��}9���l��Z!��F��֡����6��>̗wiIۚ�/̢�{������[}�W�g��kݺ�m�~m�� �ɘ�{����� JE�S��쀀���#  ��V-���_oݺu�`R���?�"�{K�����2#��}�7����v(�m��M���� vju{�<;��=��o�3��.a���ӕJ��%�0?���X�	���<֋��q  x����׶չ�>��e�'_GGG��o����н%�a"Sn43W���{��z���gz����x�^����ڵ��d2�`0ؚH$:�l�_0�����LSgr8 �ǙQ��k�U[[C����]��6����=DC�y�J��qCr��&���ۏD"ZR�=3�A����۴����Z[[�
<C������;�6=�  x��c���̥Z� �?+�J�wzR7�a�200�t���q��^��֔�����d���?�+O�O�ן���y��N�硇��b�������p  ��6ʍ�]�*O	@@����[��V#C�Q(3�>�+����=�Ng4����ǵ�ӯ?���gI~UM0����   ���5�o]�H$����8O�6%�C@���{��W7��@�Z���C��E"��կ�C��^��.�J=Ƅ,գ��3�g(  \"�������Eǀ;i8Rp �w�;����1��V����No�s��ެ_[g�������<����'��)  ����_7��Ommm���L&�hѴk������%�c2�	�ϕ������޽�7��Z�nJ"�(佌"h�&��	  �C�Jm;�>�J�xF6�5�K������ޑW�6�-m��	��T-�ɕ/�/�I�[ߧ��	۬Ujz������%����< �z9�xP��i{�r��Q�wޢgz�;���i�������ғ���=67i����LBgz�ԋ��z��~�	����C �Fz�2˽^��d.iooox���[��="�Ճ�����1)}Y�|҄v�]Z�_O�k��}�Db��G=�H$� �ztk��q�˘��L@���9to����֑ώ�P�&�&����jy����c��8�D�эZ�������ݻy��n��ض�:�=�  &W��;��t��?3�ݿ�￙���7���Ic���A��x�n_g���>7�<���ӯ��d2�lݺu��,�wA �$2���1�N��k3�`0� ��н!��sB�P�̞x�Y�}p�x�'����o���k��L<��������>�)  T�Y�����w�^�0L&�٢����A�'�I/���t�t���\\�M{R�k��Y���~�x.�����
  �g&x5����H$�+	�dno�D"]�&;L@@�y�`0f	0(��Cz<|�|h��N��k��{��� �|C��+4���`���tC@�'҃��d�AF`>�5ˏi��\�V���=�{a������ %d&v[�ז��Zys*�ʻM
����^��;����@>��`0x�=���[�J\���a���  &ƬY}�� ����֮���L��pd��>tH��yt�q�A���v���LE�wk^F�X0|��[k ����r�^�̈�[�0g*O�(�At�K���o�wgzЁ�1a�d3K�n���8f���}}}�V[��^��$  �/�e��Uz][5u��5���}�WJ0���~)mx���Y�C�G�����:J��������Z��F�5n�ϟ���k�L򿑀 IF�_��:v���X��ѱG��"���]NO��k��3IPvf��X��������h��������U�3gΜuuuG	  ���߯ץ��]xW<V��E@�!��_A�k�!���7]��cu{��3���[[[�M����o��� �?��k�F�ͨ.��h"����$�ɎH$��}��F@w9=�v����C���n��L���˾	��2e�����O��� ���<������@{{��z}�P��{T�C�Z] >G@w9=�v��eYAzЁ�b�U�����z{{��j���6w$���g� �E{�z�A��LyMMͽ[�l)�mT3̝�.p�B{�e_ P��jy��o14�wi��o��ܤۛ4�t��>'�D� �ۙ^�'���ֲ���L��\�xޓU��ք��zzR.�SRݟ���\3^s��h`� ��Fu�C �6f~3��:=��g9�����Z�܊K@w�`0X��R���2�0;��{���x�-�J�~�6�s���7<���M�����m�t	�n�'񂆸g�� �u�3�k9�m̙���~���8����~MSSS��� PM�}0�J�K <# ��\v֬Y�
|C��z�)ʿ��ݽ7�>��� �,-Z6�yy��w\�Z�802=N�1�5��5=d�<�R��_��[{ P~f>�f��3���ǅ�q� �L�_fD���ݭ��s���   ���-m�.>VSS�����' ���h	���s�    �/
�kkk�" ʁ�.t��Q�s7  p 39գZ�b&�ܤ���Tj� ��)S�l����#��[1=���  �2s��S��+N�8P�m"�m����1��Й$  ���m�{���X0|<�?�uG T+3̝�w�L1C��>  ^��r�ƛ�iںuk����U��v=v���.fYֳ�>�q   ����~b۶m���iV��qL@w����=�  �c���L�ۣ����N�ߎK@w7:  �=m�/:�z���]�q��"��  ��h�~� p=z�	讦o�=E<'�ew  �!ڶ�# \�t�����q2��  �Ĳ�C��iNٕ�n�o�E<'#   B:�z,��#���eYE�,C� ��Ѓx =�tW�70C� ��5T��F:��Uv�=��]lڴiq ��i$��֚5�%
��[rp�)��H�Hoo/��Bߗ����+>G@w�LSSS�Ob�; `<&�O�6M�N�:G}ʔ)�eƌ���#{��1� T�!��	j����������ݽ
�=7� �	�ӧO�b��9��&��ܹs�G���E�f�v� p�l6�'>G@w)}��� �	�3g��^�ך5k����Ȯ]�������!��F@'��Y��q ����~0P���I7a���s�A��: 3=�$qp�b�@7� 8��9/u8bz�����'('m؏?i���׋���B����R�����!� ���,����}�}}}���eD:�r�p�I��T�,�q gf^��K��3�0�e��-K ���A�#��WQ�!� �!��RC	��1��MO:Pھ�w��&���>����^E]�� R��a> ������^��~;ݥ��l���  3��\Í����K&�����]�؞p�xe�>l ����4��M���= \���^�~J\���  o��el��%��� p9˲|�]j���~:  @5c�8 ^@@w�b�A��� ��&k>��o��!���{Ճ�2z� fN_�\x�ԩS#�i ��cǎl�W�6t�*j1sm�L��@ ��a�7�ٕ�8t�g��m��M ��Hj.���m۶mo$  z{{M�����E�F�{����Օ+W2L�k�]*�͆�|�c�v�VY� |n�޽tx�	�}AKK�����J��@@w�b{�s�Dqt �9s?xOO�L�2��?kϞ=����f�:�ZӦM�})N�K�h";3Q\�  |o׮]R[[[�{�M07(�@`��<�[�t�盛�������Ԅ�E��{M� ���ֺ�����~x�)��o߾}Җu�?���~֬Yf�����B��9�{M�%�Z ����o��)yH
�mG�4�s'�.��r��?�%��=� ��1!��g���3gJ)��{M�'��������y��6l�! \E�5ϾC@w��ރ �L�6=�ӦM�ݽ��t��a�773�g֎
9��.
�W�	 W�c�!�W�F�D޼�� FdB��ݻ���ݔ|z3����`�I1�$��)t�uL@�2�.5�5q�A ��q���pSL@���ܚ^u���M1C�M8g(;&��"i�MGqD�ƍS�5�ZRS�UE܀��R�@�6��Ӄ ���z�@��Ao�B�����qj����5U���lqc@�A  �aFq�����N@\D�a�A���D꤈�p}���r   ���;wʮ]�oŨ�����:��9�U�z��~����+hF�^��>݈��b��a�t}��   1�f�BSL`7A=�9o޼����� Uϲ�Y&��[����~�d
  x�	���px�m��~�6�olkk[' ����st�NQ���iG�!�  ��r�Mq���[�~��o�?��֮];  �B �]�Z��b��C   ��Q�-��bgg��h�.�7���^�y��n0i�A'���D:C�  �m����������������T*� ez�I��Vz�(�&:  �󄴍�:ݾβ���m�q�ߨ�������,��f�����]L���󼚚���tZ   0��Mq监H$��L2w}0�[KKK� (���stw+*�+�A  ȟ>��f?�N�{�Ѩ�Q_��dnhooB �
=�7�]̓Z[[wF"G��j
  ��M�p~�n��gض�E��Ds555wһL=��
Et��8z1yF�s   �X�ɖe�<�w]���T�IP����;���   �R�߻�������S������' ���9��M$�w	   �i�zoo��h4����2��u���m`����:�L�#��[QC��8t��  @�Lv�YƭI���n��������_ 8�|B@w��{���O:  ��Yf���N����]_eY֪x<��u��C��n��mB��>  @U�߻�8�D"�.��M6wk*�J�}t!����X,^�v�@�O4C�   �h���N�퉖ee�px}|g �s```MGG�<F��s�@$������efbo/���  ���)���v{�n����7ɾ��͐���D� �G��]OO�󥈀^�s   0�L�}�)ο���ԩSװ�\��.t��d2�y^0L��i  ���{{{�h`�_���~��ٳ�2C<�@߯�ŝ��z�&.*����vF"�^��	   �b��7E�twwh`T����
��kkk�.@��\�@@@w������;�d���   ^��z�M/eFۀO����9x��{R�T\���  ����T����ɘ�  �A-��N6C�5��S?���Z�5k�F��cЃ.t/(j����>�}   ���\��y���m&�{Zr���`p]<<�@(�$�H$2��G� ��\�C�s�e8   f2��^v�qD��6����i�dY�F�-�v����L�cP@@w;='�UB ��S�ȺGYO��� @a�hyG�H.����^W�2ou�Qۦ��.��{ t�a��={��|o�0��|ֳ��"�������
 �J����{�eYw�����oض�	�,  &f�^k^�[S$��ڛ��Oh�l��O���=����%p���F��S}��#fi�ٷN�!Շo_��Y��п��~dD0���~5��6CBڥ@�P�I�B<c�6����*����@�~�a�� P!��T���vS����x�~�Y���݄���8�ZO��;�2�������h�����i�ޟ����`p��j����w^�[��v�~}�n���}�^k^���_�f�W��L�C@��L&�H��---z�4�`� nc>]3C
M/������m�ڵ�<Q��Z/��  �e�ߊ\�C�N�H$b&�����Vm׭	�;�Vﯛ��s��=�����kU��d�kx���נ�z=�L�������3;�5��/Ǆg���c�ƽ	�3rAz0t��fj1����w8��~0���C�{��=>��X��kS!��s�W�C@� =1Eu�@�OR�k@�3��l�b֬�����m۶�*�R��S� zT��  ���&f-�ֆ�Ǒ��i�����Л�	�Nn�Ѳs������'Z_/����;�L��}a�yL�~��L/�Tٷ�t�o
�C��m!=���v+(�믮Q0���zp.�����At�:��o�c�v�pݝH$�-���]��K@ x�P@>d�ojKr����OtE@�!�{����Z�hp�?���'�J-?�}��   J��^$�h��耮m�'���T[��2�����֮��ݕ���7۶�Z�o  ���I&�[��Y�#Sts�`�&�7Ё�z�,���ǹC/`������B=� @)=n���wg3�u0$��н�耞J��mo��|P��Q��m��fΜ�����mZ�#   %P����>��ϛ7onGGGW1O�f����.P*f��[��nzѹ���m�T�����h4z��;�,   �Q��L���G��־H7Et˲у��L��Zn���x<~�%W�L&�{�7� @Ih�B�w��[n�C@�=���"��� (�^-wk�Q�͉D"%.�J���m�Aa�E  P�`pc!�����ޱ��'�A�p:�6�}|t�mp�u�qn�:u����}��:  ��m���[|���="�;��綴��m�Y�E��Qf2�5�@��7&�ɧŃ;찫;;;�ը   I3I���V$)��ы��1�p}����X�mz�����,�83�|4��^T�  �"ijS!�k�c�����#�{��'P��v�|�j-���6�s�noJ�RO�8r��������}W��  �8t�/���S,X�m��'��ՙLF ����4�ߨ�Z�]/Ķm�vٶ}�V�.   E��U�C�_�e��н�Q/*����q��V_,�7�h�Kˍ�p��-[�t
�8�y�e}I�a  (L�ܹs�*�	��!�{H04}U���9H�1����.s?y�_���vF�J��m_�Տ  @�����צ��1�� t��l��_��gp�v-��d2�&��r�F,������T   O����C@?�C4\O(����{��0�Í���K&��s{{��~��T����m�J�~X   �W�q��8D7s �{��'�䎎�.=Ṕu� ��̷p�eY�������0RJ?���  �W��/�v��@4���>�����h�!��Zm��g}��YC�ZAY$�ڶ}�V?)   ��j�~��'��Wп�|t��s/:��۴|[����z�+�q����LW+   ckmkk�^�s^!x���a���D"�@$yV��0y�	�&�״��ߪ�<-��T*�m�B�~N   ƶ��'h��!�{�D'�33^G�ѻt{� �գ�ߛ2��gϞ}{SSS�`R����\�	�N  ��е��D"/<�{&�sn�B@G%���6�q�h�y<�T�{�۶}�VO  �QX�UP@����l6;S�<t��7��t�Y�9ޚN�Yn��������%[�l�T��M/��W	  �4;l(dm[p��(��S�F_��Ǌ}����}�z�%@����Ӳ�?9�si2�,hL�D"��D��ի  ���R�Կ
|������A�Lf�L ����է�N}?]6o޼�֮]; p�d2�Ҷ��j��  p��'�fp݃��	�M�5L@���SE�?O��|}]�H$����M��O��|P   r��@@/!�����!ȶmo��b�ӯ��3������w�^���9ac4�P���  @N��566�cTt����B];Z_�}�/0�f-H��mݺu�������ާ�  �X_��ڞX!LF=*�7M�F�/��܇N@�H��h��	���Tj5�����7�V   ���A���W	FE@��RL�L&�D"3#��K�����<.����ƺt:m�C��   <�����+�"�{T�&��D�ћu�1���{�U�S��B�oii�!���4^%L�  ��@�P�1�=���\����_i8?'�J��|`#�H$r����hu�   ��ܵmќ�@0*�G��rD)&���������[��~a�'��q��j0@�;K�,�����;=�|P `��4%z> ��� β�S����]�l�>B��;ٯ���/�^��I���*�|;�?"�%=o��[���˟ (	�9�M��-[�t������az �V&�s�s�n�f��������a�/�{ �D�$pgk	  ��*�9�>��i�z�nΛ��v�awvvv>#�}�9�`�]����ŋ�p~�V�"   �)����NK�1�����kK�:k׮�m�:�~R��,��mmm�	|-��{6�5�|�   䯠􆆆��Z����mQ3SbRM�4�]�8���ƾ�J���e�_[�timoo��Z=U�%   ����yB 8Z0.���^��}�x<~�f�.���ѳZ�
�B綴��
|Ͷ�1sK)   ��Ph�2�;�I#�G@�8˲�}��f�h4j�����M���N����$�C�{�ߣ����  @q
� N����"�{\n&�R���q#��ǟ5�����U�{�!�gi��  01����ظH7�`\t�;���aj*��;�J&��F"�v�.T�����������!�f$�  0A�`��B�O�ӯ䅀�}akf��]}�l6�hC�/Z����!�g̚5�MMM��`8�n� iP^wky� �����֖B�`��3?q~���&)A@7ǹڲ,zuq�\100�����.dp(Y]:�>S��̴�}g*�z�m�gk�+���8/��s}3�牀��@�M�z����"�H�V
��#z��b2�,�D	��c�Ezܛ!� (#�=?`&�����4����	 /�{!;��n^*��^5gΜ۶m�5�2kgk��/z��`2m�r��_�[�ы���i��� (��P(���VsMl#�b�Owvv�%Y�& ��Ў!�Yh	�B@��Д)S�l�%�4L�f6w��07�\�N���u��m�h0����|J ��z5�����P׮];����`0x�Y�X x���bm!O�s�1��?�O�a>�*I@O&��D"��Z]"�������x<�F�a�1�b˲�giP	Y��W"�qg�r��N�}�Շ� /y���yg!O�s�1�����d���!l�m_���*�G�Yuuu?�b� ������t���f<�r����3o���}�0* ����ϵ�Ҡ�	�F@����.]:��O�F
�.I�ӧi��*�u��������*�0��`2��k8?;�}S�TB��jՄ������lA#9��q˫���������ͥx1��k.�,�Pz"������5����%�e���2�
�k��z]�\!�I$��h�x}�Y'��>�˅B�{���.(�G�'XR����G!������q�S�Կ8�6tO�p~�0K;�ʺcʔ)3˩��x<�H��[�a� p���C�d����_�Z���������\�N�B�6^�[2�p}o����c�~C��@e��B'Ld�d2y�m�Ҫ� ntO!;/\��e�i���//^�hQc�|���Ϯ��L��1���ޯ�b�zx������v�V�, PY����>�N��ĵ�h��l�7��
��8�"�}FӋ��R�����tC@/�fm�|:�L�`ژ=:
�%�� T�?��������ڶ=O��	 W�QP@������h|��0�k��#�thu��i-��vGG�F��ؓu�+-a��ڤר�kԳ�~�D"�}m;L_ n�����t�;k���FA���s�ҥKkK�����^d��ٯ
�����>e&�`s�Ν^WW���_ ���,�η���R�S��P��O
���m�{����f&��*(������V�%R���x%��o@�9�f�:����_�444�����/zL�L ������o�)�1}m�b��L��( �]����.(
݇�h���,����&��n��+�y ��|����	F�F�mY�%�j &�=}}}�L$�+��̒m˖-�Hww�Y�m�j��������;���:��d&!a�@�,aHc��*d �.�Z�u�B�.ݴ�Z�U���Vk�u���jkբuw+ն
�X���Y0�%,If2yO��E	0�ܹs��������Lf�=�<�<��0@w'����	�ߋ��ζb�a,��?kǒ;찄ڕBDT�������|����B3�|>�i��)�x����E[��l\]]�������t@(��ܼڪ'D�~_"��������Ec�M!څ`0X����|\��
����Ocƌ9���!Q�׏��[kkkO@;�y�����L�"��T�F\p\n��iG�\*�L/�g��DSSS��g��M���_��~��҉v���8Et}s.�FD��u����u�H���ժU�6�7�X4�5�v?!"c�ގ�s�� 0@w������� =�����t{��������ի��hp�����o���jDT�����C���[�P6~
�G19^��h�f���Ս��P�~c��R������;�V='.�G�ɤ��:J�G��]˱�'Zq��G�*DD�����Bp���h,��ت��
mS$y5�o۶혒��AB�� ݽ%	M?y��'lnn�@��g^$����sЦX.D����C�=��K�Q��I�R����eb(�����8����?�I��c�; ������4w���ߋ{tM�)�5�l���7�fc)DD��RII�L�k�p�����N�x<:��P!�By!���Օ��q�p�c��b��>=q��AV�Z�"i�aX������D�h7��ͯ���<BDTwTVV^���x�%��'�}?�ٮ���l�m۶�p����V���~��Z�������Y���r��T*�-]F�v���j(�w��4!"*�Nl߈F�w��b�����Ѷ�+l���m�w_���h��"4`,�\.��ni�^^^~WW�Oq8D��Q�|	���	��|�@YY��8�"�a;��bq�H$����2�໅�HDvz:���q}zq�� 4`��d\P����ˆ����iR<����pݺu�B��@���3�c���0�O&����eRb�ؽ([���/��l��l����h���c��C0=�X��was|������W#��cB���	*�[q�""�%Qw� ��Tl�~F��_�������QޥR��t�7���"�I/�Ybq�����@ ��'��\6�oyG�� �K)����B���5�߅�T��3��S�T,�9�:	յBD���[,�ǟ(d	�NC��+������q�M�.D`~�e��Q���p�PA18'�қ�^��������E���P��o��Q^���z��`08���%�����0�a��l���ݝH$��Cq��=�Y---MB�\;���!""�����\���^q�X,v���(/"�\.˫�B�a�N�pj���zSSS[ еKO�%�݀
��b�G��A���""��N:O��ի�Ņ�����u}t-"�֖��ҿe�@�C\���,� �z�⚉�b�I+�7�&���ҽ�K�(K����s��dpDd��خ�F���щ\J�v��/�&Dd�g���;�y`:�'d�1������V>i<n\̼p�b�����24r�
Q��pY[[��p�+DD�[���8yS�J�_�����yBDVx<���;���	�:����hz��������.��Y�i����(cƌV^^��Z��l��~bw��{��'�_���P��y!������l�^��˫Y�:���g���E	�������sR�������5B��`0X��\�($DD��F��{��F��v�s:����:�"ꯆl��Ώ�n����ӎ�Y�v��Zګ�ǣ�@@��/��ci���b��a.� ���-�C!"��+�.Bc��=� =���ڪ��sMf���%��6��� ����bq��~��q2@_���h4��� ��\l#���kPo~'���ʹ�,����Y���c��r��xd�P(T���$!�1@�:���f�����V>)O���ֈ��a�늊�+V�\�)D9:�m²���х��\^�nݺv�~����)�=��BDيF"��l�L&�îR�rlt���R����a����������_/����c����Q�+���-DD6@}uOYY����WX4����N�x<O��#����М�v�(��i'�4wKt��z�L&���a���3���_@C�U�r��܋��v~E��l��w�sk���uuu'vtt<��	�ɼl4a��!$y� �v� ���`�6����y5X�q���4��JNG���\9��?��B����2M�+�/�Go
���ʕ+7�B�c������w�ѮD����l��P;���ps%�ԗTbga��O\Rr;�;_���g 8U�r�k�WTT<�ã�h(�d�ȑ�J�d˖-���!Dyp�.��%@���ܼA��*�'}��NP��˶s;G(o�Ӯ����V�BG��g�~�J։��M$���n�i�Vyy��8�'	�TTTh�f�VYY)C�e�N�P�bv����A��ҟƏS��ާ��;���`0�7�>&�7�iWj�������'Հ�{b�Sn�v��B�h��O��X}ӈ�Đ!C��siiio�>|�pٺu�l۶��w��畔���!Z��AzMMͱ�^��e�׬Y�(��x��P^1@���%�,���?������|���<grR�/4�>���s8'D}(//����=�Æ��5H׭��[�������By��������ե=�8�h�ٺ�Ҟ4q��A�}N(���.�B�� ���D뭷��98<��oۯǎ{yCCCB�����z�����vk���{|�����:����'�'�,�z�Z�j#��cp�>�"�7�mذᤒ��}��:���T*u&����s�V����k�/�~���"8���hp����gK'����=�^u��S�N��������~� �X�D�$��+�����P�1@�=9O��� X$�1`---=�k��@ 8?��L�������^��u���4Pg�:eipOO����&�W�WUUUVV�8~<B�\m�?e�8���x<G�tړt��H$���'F��;4B���C��n��b?�f|Ѯ�r���E'�[�vC�ֳIoφ�����g�u�U��A]�i��m�����՝�ks~<L�ܥ3�J=���^��(��By� �����[�����F�����.�8����[ZZ�!D��\�I�F
�h����[I{�u��n�d�7X����=&��z��7)�/ʻ�+Wn��},��G�}J��c~,{gO�uQ����(d蔍3F�}ٺu�ڭ|RT������+���(�R�/!8�c�A�;�T���$+�(D���I�O$�����Y����e�.�E<�
�NL&���qB�hݙ��|>���Uق:ecXEE�.���E�4F��z/��)3�)��h�)�4`�1�:���9eeРA���v)++��4XGpЉ@�%ݳ��-�Vg�Q|��B�hnn��ç����Ə�	Qq����d�@�ǣ��B�`�N����!@_�fMK О������qb���B4@8�>��\�R�K��d������8W H��W_��V����D���|��X쫄ܤ��S����mt�V\o�����/Q�����,�n\��H!�0@�l�k�p�g]rM�G4��KːP��a�c�9!eM'��	�lЂ ��T*� ��4(��t�i��7�������}(�q�x(�������t�rR���cO:���d2���e��N�N�B�� ������Y�#���Y�h���Dz)]Jm�� ����Kш�Q4�]�t�k�>AKKKv�ݣ?����\>��<=�;�AB��`081�����,���\]]�;۶m��Tl������'j��E![1@�\�
�.�z�tz�s��-��F�r���[��o������~hٲe+�|���������ehp}��$�����9�ǯb�M!��<8��~�k�{[�l�"�L�R���7n���![1@�\J&��P�����jLii�Nx2A�rd��p:���h��Gy�����׊M�i�7]!Co:x�~-�Ͼ��?�X�̦7��0�9(۾�MoY�����aÆ}O����[��QA�x8�G�|8o +f��������/ITH�PhdYY�S8�_��aȐ!��շ ?�KC&�'�H�W�X���G{�������*�JUc?�3{]NG{Mt��ªD�v��a�V�3�|����C��7n"��9��|��8�
َ:�j�ڵkO��A!2*�!�Dt)�IB��s�=�9б�p��:t��.\��I�h�3x�Q(�@����`�i�>�G�
�)))�3��z�@R��h��%�ȡ��D"�<���<��:�5�,�:A'0A���Q?e�{��sQ�_
��64v��������D��A�`p
�K�l� ��n��-//����K6lؠ�!!r�?��q�@���)B� �r��~���X,���E/*��px��.�V�^����&��y���j\�y\��fu�5�����V}}�B�9G��eee�A�������<����l�s�B�9eB� ����K��.P��(������)D�3�����ǵ!>W�CCÜN���fM�%[}�����h`�*]-�����2jԨ� ���[�L�r��ltH�W�
�:�.���|����� ���;O��z�ip8�����+Vt	��s���op*�:�_	ٮ���d2�KS����]�A���'�;���(�=��c�¶�P�0@��*�x<:�J!�Y ����h�h�|��>�Ùpr� � p�~��y��oѢE�����{_֖f�h���M����C�u}6Jg'^$TP�i �V[[{�U��J�Ap�wv)D@�s+�����l�M������|8_*��� ]�p������-[�Ye�(cI,{2��|�9}>&TP�i Ftvv~������I����6��-����zk�����A����1@/����'***��ᨾ���a�z����v.�F�����nD_!Tp�i@JJJ.�ÿI��K�7�@`�l�`�EV�g�ڵ��r� ��>
�&L����&d+��m]���]=&3�$�J'C<�����u)G�f�4P~4pO��~!���n>���&�FII��B9C��a�B�H$���O�
Ao����Z�޹��krx,{�� ��e� ��d����p�=�`j�Y�H$�B�?��Nw�F��e��K��P__áw��e���{�ޞ��..A�C��X,{9������"��:Y�����@!�P�,4z�����!:^�,�s�6�~�t��^p5�w��>����:8�S�p�^���j��ȑ#{'���qd3_�����+d�d	TBWc� �,3q��A���$!���#F<,�/�كn�,�z�����rɂ���L�K���X,�j6���SVVv��1��%PQ�������h�t�@ �{)DֻG'{�YMM�^�q�������Y�fM����,Y�,��Ïf�;:y���oذ���)�t��{�t	�񃅌� �,��x���	B4@~��fT��Ky�����~�g��vsxA�:ͺ!N��4��s��������4HO&�B�'wD�ѕ�<0=��kBFa�NV:�������e��S0�@��G�O_�fͿ�����f9o�ĉ70#�~�gv*��!s�c���:y����u�V!�X{YYY�7����/�n/!�0@'K���\��,!�@ p*v��<Au�P�!(��f�iӦ�
WR��+�������������{{�u\:�)�
Υ755�e�ت���8/2t�
�����\��r���݃�#D��e�<�~����w�=`�C�D�W��***zǥ�RlLy'�Q�2�#8ײ�s��:Y͓^���)k�Ph|ww�.�6T���x<Μҁa�n�C����H$�D�V�T����3@{Zt��=�B�_h7�:.�{�-!#1@�|�| �>�	*�����F$������<Bc�.�~�5�����B&���l��ظnʔ)�!0:v ϣ/VVV�l�\����5��f�`�Zf�2t�/���}E�v#�m۶m'��j@�e�P����T�B�8O�0aَ=%Ki�����Rl�����-D�B;��(�Z�/�{~����S�|���݌��h֮]�+T*��<��p������*O&��b������B�s-��Y�M{�;;;�(OD"�g�}�A���:���c�N���x<�`�����_���ko��<��h�N�5�ͅ����p�憆���m�/_�eʔ)��Ϊ�D�IF�)۶m�]�����nt�R�K�}p(������0�S>}����'---����DC?�u:��ڼ�+Wr`� q�5�U������\!�i��ez���k�:gy���E.٪���:��Z�h�)�<�T�:�O�4�m������&(��$4`\b�|([u�$�6õ�$v�`�������y�fٺ��P���󮭼���l?f̘ax�B�c�N�v*�����ǇP�,��!�GK<A�
�
��0��P,{U�6:����^'<=?ϯCK��ۛ�cә�BiW�Z�jc�Fp�m���� ����?^����(촗�����lg��]K��˴H�x<����l�rfv�􌊊�ޥ�6l� ��p��sYV���탲�!G`�Nv8�����^r�Y�fy���+--�;�L��}z�`κC���|v�!�(���F�q!�,[�������q8>����iʻNǔw�J�n�fO�^��j<|��#0@'[� �vG
�����wvv����N޴i�NpC�B$Y%4`(�k�V�e��t���	�F�%�sp��2�WS����{'�K��$�2w�nk���>�/���B�� ����`0x
����R8��Ϡ���>��ڠ׉mt�"����p֙ �8��^UU�����-B�I���6	�����>�~���D"r�M��������P�
!�`�N�A�u3*�g9�xL�6-���}���n?���ʔ��ٲ��C*�-۶m���%pm3@w�Qhğ���B�ill\�W�p�]��ȍ5j�������ϱ*f�onnn����@�N8'��0@';����ƞ�Z6u�ԏ��>3�S^�����	l4���p~�Y�n]��U�;��K���7����~|�7����ǎ����>����>�<]�����w���1�`�ItN���I?��/���VZ����q�l�:�[SS�!8����|{�4zg�%*��[����������	!� �sz��'U���ի�ⵏ��~~��+T4���.�����4��v3�v�����hg��n>��s�7	��ZZZ�I�Dz"�����NV�~�zNZC����^�� ��ߝ.�� �F���-���/㳷��3ӦMۻ���_�G=�'���B��\�q¹pkI_)���9������S!\��ޝh@�#d�ɓ'�FA�iM_/++;�4�?ϣi�ڃNT(ڃ��)�-S]]�Ǯ\�qp���@Է˅�4[�O3�@�T��? �{q���TTT܊u|�����6��.��p��Bl~�JsЩoЩFz<M���PAM�:uB*�:�3�LGcn@������%D����!ˠl`z��]���B��90�mev�.^���Uz����CxOwIC��H7�^��9�O�8qP�Aȉ��Ӯ1@��@E��@ ��h4���m4Uu��ɓ��>����O�Y��[�n�݈
liKK��B�A�1�		ΥA�k"��![466������36���|�ѢE��QS�5������9!'iI�R7���6m�&vC����N���egЩP2w�XQ�ٌ3*�l�r�������d!�.��\�;'*4Mo�ʎ	c�=+�u���W
�&�&���'�L������a��#P���m8�[�x��.�ebe|�{�w�+�*--ej{�S���n�F������G!h>��	(�O�?��k��:c;R8��YJ{Ѕ��k�P�����\^�&�)++�;�v�K�i���"P�;a�F�#=	,��H$�h.����Z�F���������dz@�~��U���Y�h���5�,���cʏ�V��^/=�tR��d���h\�jНo��+��f���[���|�a�KO�:u�G_y�]�ijjj��$���	��<�ħ~�ZZZza.����>��x�C��S�i����Q��m۶�AD�r.���L+�T*u<O�I���YZ�|Ҟs.�A�`z{��
9��o�B�_677w�"��nw���R4��{{z\,��������G�8C�8o��kuu.��v�fN�:1a�4����ȷf$�.����$�H�)�n�����ڞ͚5����t5(��T�
�^8c;f[yyyN���g�G�^QQ���㡮�L&���B��g��V����k���e���5kZ��#�ӥ�~�m�P��k̘1������.�{�H�����,̝1@w�����S�J���p���K�v2}������Gy<�����[���Y�eb����xtժU�,U^^�����mԷ��bL��544$���\^`�KO�4i��ؿ�̓Ӂ�����z����BI��8_ϝlA�U���Z���w7䒓���K��bX�ua �+��KH�M��w*�:���4
�a��a�^�M�6	�I4�T�r� ������u�Ї��e����;kj}Vzƚ5k��k~:Α����q�m��.�=����mذ�r|o����Im�a�N��Tf��R��\�9��ĥ�����OԠ�'���S3/tR8"�l�k����������m�.]������8o�K�>cƌK.\��D1h���o
O`���l�Ͼ����D��f��hO��k� d�E�	�Ju?2���N����@���)��35�G��Π���GV�Xa���b��6T���b3���h������p8��l�1b�ћ6m�N����˚�
�A;�Z�x96�P^y<�o�������tb8���ˊNL������^<[�lS��UUU�s����)�0��L�>ɛ_@ӏ4��3���� �+��lك^��Ǎ�MR�Խ��Е��ޯ ]�g�����f����CBy�vֳ�h��\~�ˡ(�g��4K����S�w� ��t=B�R݃eee����CQ��CP��Ù(HOľRf������)D�PYY��P��*F��i�]cc�h�;��u��8���@�d�󴴴���8���7=:�N�(�_�w�������͖����-������]�^���b�qYMM�}�^��<y�h���iM_Ǐ��g�}Ie���ٺu�������r���P�қ�'�E'���ͯ9���T��=8�'�F�:��U(A�p�?"d	|�?������w�=|��0�w���1@w���R��.����������:��AW�ԩS'�R)m���x<���K0�HpR82���'
�A0X�XÑH�A��߀�c��j����X,�(���v�p�w+�m�[r�\���]'�۳Mm�]c��2}��+��4H7%����@ ��-��{�L�<y��������hF�N
Gd0���Q2�
5�]W���P(�"l�����|]�U>�K�.^����3�F����$���8�&���C]�r�ʜ��Mm7n�d&���c��2�
Е���$`������������3f̨زeˡ�S^__����z�05G�&��N�CY�(���� ��w��-�F��	�A{�mСu�i��n��y�foz���������S�;Y�%լ� �e�4CfVwC�ν=ύ���o��kРAG�39��I��R�8c;9�Lo�#�9yO�өt���	��s���~)����ny��2���`�q����l��s�\~a�����J���NG�`��2��AW���:1�!�������/����'O��gq�P��*sKCUo�����Ƒ#G>+�7hlzz8yO��w|����Hd�P^���K���gpx�������I�&�_�l��|���?h'M���������u�|V������w�H\�WS�u�9Y���dd�E���������+
MJ�Ǚ7S�N�h*��J���M\�"�t�=Љ�	�������<��u������m��eKKKu�����"����c������~�P_��D"��:�#v�a�3k��F����̞z�3�]�2y�D"��|��'�5k������~'[���+.�7dt�9Jr�c���{������u�'���G�یm�ͯ�i�y�3���(�g���s��ϰ�؄���r�|���@@�(7=��Lm�t�^lz�m۶ML���*N�:�����wvv���xTV:�|��{��18'�H�LxJ(�j��kJӒOʫ����S�Ly����u'.Y�Ė�����玚����މ�B��\�ǣ��ڿ��8S~ii)S��:�^x���%�������$Y��EP9�N)�4!�����un���DYx���e�P�L�8Q'�#��g�����b�W���~)̐�3�}��DY݄s�H�[��ǟ�͙�y����>�}���PcEj{��;c��2�^z�mݺՔT�����.���==Ay������\ߥ͛7KggNKp�k���ٻ�;���2o�]tFw�����Ѯ3lذg������,>��g�;����(�zw�?�Y�ʹ7���>hK)�Y�|W���`1�f�Z5y�>���c�B����ݔTw����z��5k�����������)��+�A����sR8r\׏���r�����h���Y�parʔ)��^�{ү�p8����S
`����(����|gc�c����.�9�_$N��i�V��38�tڣ��D"���|)�z����#3g���'y���T1p�	�����9��V
���qB��Ʋ��&�W���m��;=Y\A���k4vτ	�F;D3"ϖ�|�ر?��Ə��Gb�Lǝ��� ���SV�b�1ʆ����~����|?W
�L�Gw�����6� ��;�?4�D�ʛ%K��\__ߌÐ�/=+_��|>VCNS�����✻M�wՈ����J.���5	:Vݸ��:����T�5;c�NY�L���M�e˖i�~�^�V�pN
GN�J��� ��8r/4�o���L[�y���)S���j�_z|����	1@,{���nbGG����؊m�[[ZZ����/�yq�F�i5��j,fv� �����A������o��b���#Gr�y��s3�;$��k֬Y,d�Aw�z�߯C��"�7�T�>�a��3i�F�j�ʕ:��b�������I�>"�A�c�4{uuu��?�d�_�������ЋS�]3!�]�L��nȐ!B���ˠ	��r�eS?l�S�����+t*t1[�t��/��6���'N�bŊ�b�x<�>]��R�x��D���$�b�X֍�tj�����b�|��g08�t����<x�13�������#��pR8r:�_�{��í���r�s��IOgw�>m�d�z�FI��)>��E{���zG4ͩ��Y�MLm�v6��ڋQ��Xq�*��b���t�5Jh�4�a���I�5O������]�����|�����"�H������b���t��qzF$Y��o:�����،�Uލ�m۶};�_�������v���N���:���M�Tw&Ӟ�͛7˰a�MvYh��,B���o�}**�z!r�5�#�w(3J�(v��Ĵk#q>�گ�ū������;>�#l~�c<��1˗/_+�JORxG0\�����d1_���׭[מ�/���?�p�FS��~Щ�2��&�������0�r:���N��xtѢEm�:�����-B��މD��fR�~µ�U�#�E��	��llv�h'|���p�Hdv� �����78#��}�K���N'��h�Z�f�~�]��`ZǳkO�	��Y�5�݅������	���;::��q�Tf����"�K�Rn�d29Z��?|�lG
�E"����ԯ��I�4��� =#����|4�?�-�TTT�ڎ�g:��+�0����0������^�����AS݇w�0�~k�6����C��m�;}�@`�NR"D�a��-zzz����d0<1�<&d��^{m}}}�Ө�O���?>iҤ�˖-[-����q������'f����K�e���jhYY�ݲ�&�14V�+���3�������BЋؤTw�iP�Z��Bsn*���v��	&��n�8{�����@���0�� ������F R����i�v�%^��t썛�lO����PhR2��
?�V��ΝxOO���5k�Ncgj;뚾1@���i3e}mMu�{ｋa�L�$o�斖��eѢEY(��Fġ_���?���t�Kmgg���� d�#F<��޾��6����;.@W����]�,�{�?Y��G;�\~!�w_�hj���9���O����n&���b7n��#G:���Vl�kO9>�ǖ-[�!�'@p�c��l�(�������F�������Z�fͿ�,�p�p8�(ϱ��?���XCC�c'�F�+�n:��󝍽���^������kh���>��ؙڞ���o��2&��wuu���:T`>3M���iӦg�>���"!*.�m�1��^��64�g���em5|������+�,�;�`���	&<�H$n�&��+�>����z��#��D�#m�۝}Z��>1@'��E�K�i`l�Y���]z�	�ls�.]���@������ЖX,��:{1@��9�����%d����皚��p8���<�ߵ�-Rh������ߤi������ ��u��k��!��d�ڍ���� �e�}!d�e��BӿUS�u<�w��[��� �J=���Ҁ#��s?��!BT\��Z.��w1�g��sK(z����U�2s�����s��L���ɓ?��ߥH�b���'!��?~K��y�A}nKK��lm�#�V�ZS���_�v� �,���Eױ���K��q��vϹҫ��?�A�����5�x�t��N�2A�����W��e�D"�k��.d�t���C���^4�����y������>��sIm7n����R��ߨ%Ք�
�ك�7�d�̝8SR�;::zoh���Ea���y�����˗o��"8��W���� �~ÄhP�����A�|!�466.���_��Z�_z�ĉ/^�bE�S -�@�5��G{����G2��h[^����%�VtR�j1�-Dj;����R�U{{{o������O�R����O�Y���9��u%A�4===K��6B����x��Xkk�Z!K�dg�pX{Z�g�K�]^^~�l������&
�K&�7K�'����Һu�ڳ��@ p)^��5��H;�t�s2t���MIu�Mu5j�Ui<o`�^�K�.�g!f�Ep�/����x�X�!���)++Ӊ�N�R!�L�{Q��y�A��4�~��y�\~��TK/d�x��T�nif)ǀ��:�I��z�` �ѻ�-�6���>�x���I�3fXyy��.*n�	S�)����h��B�hhh�O8n��d�_���'[�b�f)r8_��������K��ز�%�?h���5t_��6H�Y���Zh��7�.c��`Z���G�4�!C���|���3���ytѢEmb������>"D��_B�����|G��d���|�����U��� }Hyy����'.��А��`08m������<\W��m�<����0��9S��� �e
�ʢ��Φ��	2����A�A!�>���4�.2*���g	Q�c�n�m۶c�#�C%����v�Y"�Jݏ��&��oMswE���DtR�c}>�	���c���+�>'��:1t�B-�F�c��2��7u�˖-[�IeɌG׻���c8�?t�п-\���5�Q�O����� ��6+++�Á���H��!��0]�5���v���d9���ǚ�5h]�����Ů���G=�37G�UVVf=���q&�w���̄�v�=�.S� 93S����@{�7lذ�˖-s�,ѡP�
��\�e*z"��<�![�R������M>��Y:�������Ci"�8�ߊ�Z�j#v�<�m��p|�/d�B����Ch�ރC�&3��� �e
���c��gƔ�T@uo����84>@��V���爁kh���+Wn�t�h � �]WW7�o�Ѐtww���	v�4wW��x|���jii�*�+
U�;ӎ�Qbm������1}bE�2���p0)����wE,�+�{��Ä�%��^�������ɝ��:�R�Y�lنp8�$O��u�2mڴ��ŋ���p.��IK�}|2�ԛ)�b �b5�l�'}c�N�2-�]z�R�]555�����NO��b!r\�F^��8��C`s	ꮿE"�ǄJ��mС��b���&
_��+b Mm�,V���O��vZH��D"!��J�	�BS���7�A|>߇�`�]�\���l�t�H	�wjz0��5B�6|������:.����E|�0@�Jz�_��LMm��c�N���:ݠ;gux?� �L:���F�=���8!D.���� � ��d���2��lԫG�R�:�;�ᰶ�h�K�?y������ �M�~��}M�s�tuV�TzGO�^ۺu������׈���i_!r!�+�l�@��c�BG�^�R�; �&g���b^W'�c���@`0��y8#*--��L���>���QQˌ�1(�]+���~�k�XlN���Â`0x
/}/�E'7���ںV�vڃ�Y	��u�_����ꗆ�������P[Wr�ww&��LH	��N`���]8�"�^s�V5o���˘����Cǣ�RƔ������D���
�f"���x/��p����P.��YL�5�3�ɨW�ʙ��pXW��{�Xߔ)St�����؝!�2u�����>1@w�^��+Ku��	&Lkjjj+��A��_�`�b:���wY���匧�:Y�۟pn���y����m_���i��w�6�1�� ���T�S�i���������P���3��hnn.��p:�1c>QQQ��	BT�8��@<'�|9���]����r�dɒW��޼�un�9f���}s�ʕ�B:)�~('ġW�YΘ��:A{�KuW�=݃��s&��_�v�f��S�~����EBT���Z�����a'�ί!�Y�ǟ�>��q}����k�ȑ�c��5������~�.y����YP�� ��a`�{�cȯ��:1@z��o�=5� �U��K4@o
D7x�$���/N���K�R���;@W���� =
U��ϠN5hРެTr>�.crψ*����i\�����h��b�X,�����f�ީ���,TΓB�GrƦ�G?
{�o9X�t�S�Li����u�z'���ʆ����B�����t1�Sfm��fl���˘���cѓ�do��A�C�S{��,��F�O�|��t+��v\g�S��&G�N����j66[t��㓰�G\m-=W�Ce&\��� �eLox�8��a�UK�������Y��E��Ǐ?����Q1t-N��*�������#��#BYC���n����gsw]��s�h�~W����� ����C-lLKu״<��'u]r��r]�z�[�P��d2��W���%����B�w�Q	��?  ���UBYihhxkʔ)�gw��/}��<vѢE_~�.87���b�L���t2�6��k�?v����&,������l���/�x#6v��#�1�Z�`P��zz��N���ۂ���i+W��$�-Ms�;@��]6�_���S��cvk֩��NŇ��8�᥅Ζ-[L|χ��_;�͘u��K�ݔ���n"���k�7J�R�.�C�گ���O8�N����ݡ,x��y��C��3Ms/� =
U!8�{��tR8I*N�]�I/}�Z������k>��m~]���⽽�B[ǥ��A؃^Xh�'���NF����(�G�-�T__��I�����4iRݲe�VJ�=z����kp>AVZZ�;����\�����.-|4�=�H�iP1^WE"���a���2����}k�n�l�D���xV�s�&� �@�z���-�-ʆ�����M�ӱ�^�P8.�������d1��T�K	3��� ������G7����-hP�E��^1L$YSUU����2}o��tww�*�mBT4�g�WK���nmڴ�����8i�Kk�{���y ��v���jGŒ������0@'�e�^۶��v���w�|�����sb����-x����
��d���D���5��D{4���{�އkkk��Z�j��.�\������!\�_�����Ó���w+ʿs�pŒڞ� �o���@�M{�4�������3\�*�IOdwu0\�K�'�#sŅ

elG15�ȑ>��Օ�4�"�>��Е��M������/�e:��	o����8�NUfVwC'0�B���wx<��(�<�����=��:^�̳F����ڶ���;	��5��Ph��-[����^ol�l~�3f͚u�9s�Z������M� �[@���>1@'G��i�֭b����)4*��ok��盂~~�!Dfa�^`�c�p8H�
�Z���G�ѿ�I��p8� ����njj:���`8����O،Э�M�IJ��o����ʠA����KU����	&�ʫM����{<����?^$D�@c��tmK�Th�U�ǚ�������.ԧT*u���)Dz���;6@��|���á�cz2��{0@'����2w�޺D"�t(�Dss�1!���@ ��߈*(*~h,�%d�GQ�G]�Pmm�TN׷��Ɔp8�?b�K�VWW���N�����F�:*�C<K8V�U��#��L&���|�O��qc�h4��������y(��
Qa��F.�A��o"��u�ɜ4�o�\�����YYY�i�	��Y�;v/O�/�5�٣�.�]�X&cp@������@8�lCCCB��������l�S܍� ������S?���v���>�����ͪi�	����\z�{��Z�Lmw'�ʤo�L�E�A��w��Rd4@�����L������?�s���}�:�](:�����YBT �F��n �W[{8�.��{�W���+�>����N���O��V���~���h#�����qI�����tCl޼9���۶m��jZ�"C��3/�!Sx��k�;3$u�R��󚛛;���~�Q0�)���A7 ʩv!2����jjj^oiiyC�f��zʋS��[6nܸ�^��iֈC�%���c��� ��pb�wp3�oZ�|�����.�F��)5��.�L�Og��s����.|���|�$��n
��ơ��"{��]�v��	�=��tҸUUU����zO"������V��m�v����-�B�k���Rs��8Df�����/����<��SV?��}���۲�^{���gㅠ��09�=�<T���ÿ�H$�K�{��g'
Q�Ņ��=�%�� s�p�����('� �/˗/_�u�3�۔{p��ɓ��ˀ
�B#Q�=���Aܐ�N�� �@J��~�<��_���N\�O2��ս���"��Y�/��b���3�|�w�s�%D�e\�έP=����s������q�E��������� �3���D��d2��A��������1@/�Se��y�	�ǎ+��#�Iu����f0�D"����)ǟ:�
�K�|b�n��==L;$���1�M��F�7	�*++{A��p8�����1zmmm%>s>E�M���k�� � ҽ����z����6��g��1XG�����f:|�����X,v�8������� ~�"�1@7D*��\R�wr�Q7�7�8f��|Z�hѦp8� �3m~�ӦM�w������༫�K{��0o�ܘ�κ�o�c��<Y��g�b����	w�P(]� �uĺ�h �����b�,D�k��t!r��u#H?u�!�����k���]'���|����Lm�az���a�dp��9�]�߂��^�=�;�,����9���F�~�8 �g������<@��tC�t6��A�|}���O�����'��f�(;_��YR� m�h��p��KKK{7�g�%%�Iߓ��@�������?�1m����}>��6���~kx��BN��D"!�m4,��x����ӳ�^��B'���'���� �\�����<ZUUuxkk�q�+Vt���px��/��ɓ'�l~�L������L�ю��o��U)��uS����v��S�fЗ"�����8vě�F�����x��	��0@7{�ɉp�N.++���YN�G�H����3k������셶���āt���æpJ�^T-�=��B�A��ڸ8_{�QP���E,{�y
����1B�Oh`q�!P�l"g�����-]����zM�����h�>k֬oϙ3�ێכ0a�X�:��Q�gh��2[)wN	�m����cѕSݕ���=���{2:z������4޷�����f9����F�s7�ȡ�Y_�r(�����i�����������bƽ�曟����~���Ǐ���~��2V;�܎�Z}sJ���D�pS�K?'�����ƅ��Y����;S0�7��q�e�P#�������(b���R��g�Z�})�t�{^�����׫�Q+�C1Y�Ү0@w!���+�;u�
]z�I��jkk+����|zR6G�D"���<����!��:!ctuu��E�p:Q�`0x0�U�BK�,Y�_�{���:m����x饗����>�6�sbs����Y�i��rv0@����It]I-u�9�9����I�'#H�$�f͚TЇ����GM{w�� �����nݺ�@ ��;IN��;����N_�j�Fq'Ms�����H$>��_�~⚚���M�i���P�6)��8%@�t��0�FCMu��af H��gt��8Dz��U�`�%�Ql^���et��Dq����>���5ẻ��� (��S�����x�3�� =�N:[����-aj�{z8�ON	�كn!7^��8�n�*����}>�1�x<*�)�x�i�;λ�QИc�n��� ���g�~�mRD��f�W^i
�Ë������:nҤI#�-[fɊ��>��|����:::zۤLq�N?��;q��ẻ����;w{���N��~�������ѱX�� zS��x�����	gy��9&;�E�Q�8/�7��T�G�D�5@�
��b���>Q 8U'��a�Ly�K ��H҅��.8��(��z]���|1hjQ2�tb���� �����w�8H:��Z���o��X!Jc�����"�z�{oE����"�T���~&���u6���`�B�~%Exc_�t����렳�oN	���mn�X��x\��N��ٮ����y؝/6�d��fuwh�0�tOA���8��g����w������=�Tlz�_C��u�K�����L���<����x�t���W_���������D����+7�=��� ��g��@��ʒ�gk��i4�t�ˌG��4��c��ΊF���� ����Δwb���S1�����t� �)nk�����y.�������w�9��3@�3��P�ϐ;Ү�^c��� �Tw�J��yүB�~�8Lz6�kQ	��)�8'�Z�̓kt}	g��7��'���imm]+.P^^�A�%w��/�i�Y�uuu�h�܋�g�����t����z�D��	yo�����6l���i/z*���J[�7!��ǯ�y�?$�=�F�A���ŏG�Rgg't�x<��l4Q��zg��盁�ӑ˻����G��)S���������u?�dɒ����u����..�� ��L���/d��ŏ���*++�7���v��A�N��d%%%�!H�S���h��ϤS�u�wN��.=mmm���<Lq�b7m��Q�������i��i�&���{����C�=�m?q17��A���ɸ'�8|ۘ|��СC�{��I�˙��������IyOb�)�r���Y��,Щ�i*���o��R��j��KZ�m��)�	�Q�O��1�c[�I4H�6��:�=��� ��pR6!8Ԃ�lZ��#F��ݨo�ھu��b*�x</���t4}S�{��ѣ'WTT�*.� �8�����@nq�MT?��HkhhHL�2�/h��]�~h������Ɔ�|�����v��7Zggg��-A:�z���\� }jyy���d�b+���u50煽kE�ghϳ.�v|<oZ�n�.�x>*�g��]l��O�c�n �$N����`0�D�"����蚭�i����y_��Nr˕\��A��Qu(&�t��BA�w5/����4P�v�2M��Tm]JM/�=�w���t�"�3��Z�pώF��C��%
�3�L�?~Z�(�:d�n ��N.��9?���=�H�Z�dɋ����q8��>}֬YW̙3�;���������x@�av��t��E���͍.�����M�����&��X�������h4]��LW=�*6L�6P2�\_V�%��4������C֬Y�"E�h�9�W��������=zt�%���ㄲR���==�+�]ȭ����*�Q����8ûJϮ������R��q<U�h��\'d����-�@����*$ڵq^��q�7�����0�(@�.�D����ߊן,����tr���%d���0a�)MMMm�Ph,�����>����� �Ě�8��P�4��B�.M�R��B�����;��466.��+p8Ѯ��T�7��2Ž)����b��Щ��s��;8$�H4��a[&�^���555��{ӧ9'#3�s�n���:�A\���-*�����#;^K�_�6m�}Y�a���]�M��&�˅3��  /�IDAT_'��gF"����ZZZ^Gc����Y`���;��B���r-�1'���9�)E��h]/y��ݵe˖ލ��A�~��b/�.�I�4�]�sz�a(�
ߍ�b7�8��E�7�&�-Ob��7ݑ�=n2ꊷ{xs���"�1�h4z��W^y�)/����x~-76l��^�/Y+�H���ޓ��e����.�̘sꓮ����7�����+WnC��5TT���s��-�F9	{i��b�я��`[$�[��Φny��������)�!ݽ���v�����	�r��{� P?9��G,=���Ǐ��J�~��g
9�/��
e�Z��DR����o!HZ�D"�x����ba,���oܸ��/�8=ݝ�ɮ1@7���`���ly<�z�Y��|A08�هq�,F��4<�[�z�[����|'�����BF4hǠ
�к�p�2�+�n�D<o�"�|������5~�ϧc�7o�,d/MwW�^T� ������s4(�\h����<X�&nlTq�y��@���@ ps,�:��hh@ͯ��{���C'�����3V2�d���F=���x<O���x4])E �N7� ]ۮ�k��慣��vLi@Ł��C��~��ٹ�@�KG���ȑ#]u����1��wt�������=kժU���c�/��|�C#�g8���i:���k(���d4�'�������:~���;���_ݯjp��慗ikO�S:�X����t#v߱�y��|�w���R�.Ŏ�������|���洖��7�����bw�����2*g��,�J�-)a�;�Ԗ��=�:�H�/�N�[�hѦp8�+�����j�����A�A�=���� ����.1@/��I���]M�>dȐ��{1�έ�ss4���E�h�.)hH=��Ȥ��6My��H��¹� �`Lq'ڥ�=��)�444�l�t6��t�on6m�d}N��Û;�� � ��	aw���K]���y��#�D�>��������)��/Ǎ7���L��M���G�p�P�b6v�صmmmڂb7�Ύ���G���[�>���]���q�Ro��d�$�?�Iw>腡W����$�^L���4ʻ�&�ɩ�gF��7�H���[�3�����#P��ߔ�7%�^\�`zC׾�D)�
��:g��~-�.�Z�paG}}��%%%g��q�+�iӦ�V���tb1Hw&�6C���9����|� ��)%�kEA�9[#!��b�9RDғ�\���7�6���
{�m�Ϝ=���k�:Ѯ}#D�fq��l�}�Liw.��� �~G`"6һ�:��.æ�<)CflMǭ�m8Λ�9����+V�z*1��3��Կ�m�P^�:f�n8���i_!���	��w�:o˰aÞmooכqcv�w�tX�3bJ�s���-�k���@���A�NI����cg�6��Jl�~��z)���p��1�F�**�kjj>����$E&��	�\U��O/:$dA�tUu��!�dXd�Ȱ��0#�D�����8e��������HDǀ04饖�N!		����y��{2E����u��.��y��[�tuݺ���=�w��I��9s�|����L���eD�P����x������ �|,�H"��3�-[��?��h~վ�`���D����l��F����>cĸ��~��k͹��X.�{!���N��1�������[�}��S��pǅ��pEн��Bb�0��$�*�L���<���y�7oVJ{���Hg$��Fu?��_�*R��ߜ-�sO��c��1�n�]�n��&����������K����f���F�Bmm�����r���	1f&��z����t��#���g���̦M����L(�m���uo���o�k�I�s�
�y�/444�MSS�i�Lf�	(�:L[|$����|���u�%����^�B�T<7��={�!��'`?}����(c&�H���tE�]�/�Ĺoh���}*�]�N�����	�d2������|c�֭���-��5�h�2�"H(�]�q1B�<?Gx��9s挺�:���г
�H���t�o��@��_i��@h+5�����h4z(�NU�@��ں	������T<W_��c�;�X��r���4����(�"D1���u���.Λ�������Өj�Hg���j��[
�GRt���ȹ�9��K��Z@n{�״D"ј�f�@�l�#FEt�w!���c�7���=��`�j�߹Mn+ZkD(�6��LwP�~芠�����@0�� ��?��R��&$��������u���b��2ڧü�����U��D"��*%Ĩ�0�=���R?�9��b��p�	��,�O�e�>�x?�\�^�zA�"�A���G455���d7!����9�����t#����l6+��q���߈F��eb;Я/��r��R)�Wl��Z�g�b4���dB��N;�4(i�3�S-�>�zA�"�A8�05�<����y,���k׮� �d2o��CZss�\8s'cP:�e�	9���Jq�8,���Y0�!��Ox6.�0_f|��Y���8�͏��P[[;(�1�l{m	�G����}�+�&]�0~芠�;*�"q
N���7p�τC�	)���������x�`�u��6ل�3f�n�Ƨ�5�B����N�����XSa~V]]'��[����Gͷ�"�_����pMz%E�R���>�:�m�����o��>���0蜍�8N��I�����_��޾Մg_�gh��|��q���	M��+V���f��k�/I��w�l%�����N46!������}Q�x'�?�SI�>�zA��^�l�׳�r}�"��}OVW�=g-^y $�C	g�.�f�'�q8Ύ/��I*�z��h�x|�ϓ(�q<�E��C�"���|7�eR�G�W4 �dB�hQ�H/L�#�b8��pT��� �Y�p����~�zO��x-�]�<��aq�X,�o[�n�lݺu��h+�d���h����:)�,.�h���s� �.��2���~�����hfB�Hk�ǊDza�Hg��Z��4���;��*�fS�L1^�Ѷ=�U�>����s�x�\��ǌ�Fgg��8�SMM��p��8����4A�	��z��(��#�Ar�෌Op*����FQ���g�&�t8V�O�4I��
#�^�q�#��FLO�3�^@�\� Ӻ�"�����s�����Y��+ȳp�r"����⛨�P]��^����5�G@�؉��7!�b��m���R�u��l6k���uQ�{�@������d4� �S��a�5}�����T����b!?^��⬽>������CF����ZZZb�<����$��T���O�}'�.�
���1�^����n|D,��Õ7�n�껄��SP�-��ͽ�%҇�t��#�^%�����f�8��n�~v^���X5f�$�cbE:��#�7��x<�kp~WWW�#���ʈ��D"� ����WN�5\`��m��O�s�-�L�Aa���d2Y�½n�1�k�o��eB}%���#!�^�t^7E��NF��8"�h4���58�Q����s���򾦒H���������;,a!�� ��x<�(�J݈{V��(8Յ�Q���9ډ��xW���g@����(r�Ƙr9ƖV�3���v��x�_4!���y%&
%��_�]���E��8�cq,���(�=k��p>$켸�۽��ya8��/����ȟs�`�R&���>���䫙L��F�G�F�'�^Z��x"�?m�U<�]#|Akk�&�Q,���G�b���c�*�3�u�����}ߍ`��(w�|$�Q��5�q4�פK��	t���7GQ�5�]
��,��M�Gȣ���Z<��$��]�"rc������E)p"��Z�s�����m���'zLk�Q&�2���o�R��1>�)�#42!��Q󑰑t���P������H���J<煱i�c��c��a^�x�=8B��t:}��z��p"�Ki��.r��s����>X�?It�Bq�o$Ѕ_����d26>dΜ9S{{{��s���BS��=�X��`�D���q#�]U�#�B��@H��q��֦ocW��h4�w�S��KFM~5x�?577���k�)��П!��#����P�?�>�t:���!Lg�w�כ*g:U�jG�G¦��x�aAJMwW��0�!����ya�y�G���e`�VA�9�<D�b��P_oĸ���|ڢٳg'po}��I�+6C��@E����Z^���QWf2��Oinn�q�����x/�Q"��t���X�N���i1(�^	t�煱p7:#v��]錨��_L��<�:�%�8�aQ�^�7�p]�pM���?	�pBq(��#�w#�ǰ�ߘ���S ̧C�]��?¼�Rˈ���þϮI��H�}8�5�״R?S���bD�"腑@%c�~��7�y>�m�k�s�՝�1����/H&��e�+�R��R�Nq�}�)2Ǫ�J�����|��r�����4`^�>�wۥY��c��4���nB�W��#a}9�E��NO��?�x�;H1�6>?ݽ�H���(	>�!/^6*n���;�I�&)�>ćq?>!���󻺺:�p�uF��:v�v��0ŧ�+��/��.� ��܅���40>�������	vk`�	9I����%�ON~�u�:~4����)Ǔ;�H���7V�+�}d�9	E���G@�_����}g�1�2�����l�ꌮjƐ
@t�~�G)l����u�d����M-�7��3!��>�_������K�ƶ�1E:��Ɉb����U	������ѱ���th��tۡ��I�E�H�8CW���h}z�hoo���Z^*�Q8?�����	t��f����Eކ�������4>&�HL����&������#��E(l��<�U��H:}N^cl��n�[���Ϳ%l誉q!q^[�O�ފ�����ۛ��.�F�W��{Ȉ��]*<�p��!�:�EG���1�+��G�Y��<C}hJ��J���M�H�իWo4>f���<?��5�L�[gN���{~���D��t���r��~N�e+�>>t�D��!�89�v5R�6��c__�	;�^����X,�$���u\?���ن�m�3f���"��0_G������5hF���ӿ�N&�����~�MMM'����1!�F�k=\����cЪ�"�g�A)"��F��G]����jE���K�\{a��G�Yz.�?��f/Q!�ʲn�:��>����/�.��s�n�d2?�r�h4zd,�>�&��}��X�뵫�g��n儾-���,����+�>vt�B
;�b�GK����s;�ɓ'+����~>	��X8Pw��\��ӳ�!vD��\���\.�]��& 477������Ia��Z�Rm�^������|F[8N"}l�*��bŹ��}�$6��냑]D�>�h:��0����o��q��B���pn��`�w���^5`���	|���<潙�
aך�qǇj�t�u��?��־�a{�._�0�!e�t�r/o%�&�h�Gv�v�tEӷ1���pk6���:B�	tQ
o�����~�*��<��y�q
`��*�??�!��+E�#�|��
t�/�k�ugA$�CJ�Ź���#ӟhv挿���4�M�q@��p��f'��m| �]���ߟ:u꿭\�2���	�G�Q<,y3���3�L �W�9s���1�^��b�5	
O[P�R�WI�_��n�`��Y	�����]s^�`�{(�&b�3��.��/�x�}-����lֈm�֍7n<B��t:}���P�(�.��Y��C�. & 455�qr)��s��2��B�V���~&?ݽ�Џ���H����z��0�XsN�Gq^l�4��7��E�&�Ѕ�"��Y��a���D�ѫ!ԯ���c\�d�0#�.v�{����c&���	���b̼�SM�Q�|��Gd����U����+st��0������x�jQ3�w	��Z+�>�=a�!�/���צR�%�"�`\��ֆ����n�m?����{�	��3���׌���%r����	�Jߪh�$��	)#���*��Q$��@������+D���hzA>�k��E�X쇸nmmmU��\?�{�-4�!�ั>�M�7��ecc���1��H�����(�H�V�&���G=��$Ι�^�CW�}/����%��<�M�!Ͱ1�^�����������{0�]=�l�=�%�L�dDSSS��b��g�t����@9E�Xwer�=Ey��R�h�演�܅B(��j���8�hm����n�5�B�V��7B�o0B
�yF���`���	�V��>�b���	yU�|5w^K�RnG��c����	ٝ�Dy�@9nD�)�X�ܰs�`�t�����ϋص��^P�<2p\����l6�0��Ǜ{zz�!���Z�֠���; �[M�@�������0�ZF5/�%ym�6q�#T*�|�ʠ'/ĸ!�	l��{UjoI�~a�&��S��2���H$��X,� ��k3��*#D�P%��C��}�ݍ����b�
on�R��͇���}��8Ux8[}\Q�����o���R�J��{uw��!�R8�ت�+�x��q,ح������X����4�_�}M*��o#D0�@&98��R�C����ں�����Gzzz�w"�1�}�mnô��Z���["��<'U�M5�XÊzHq+���O|O�:�BP�W23�/(�^܏j-�/u*�׬:eW�pܿE�;�?�A�t?���	 ---S0^}���w�FCQ���H�Of��7��b�H�����@/w1[E����lꎁcx����hk,���k׮�l�����n��4��G�/=�J��}&���l�<4Y�m�#�j�}M:�Hgv#(�2u�������[�@%Q���rt>R�H
�Wzc��/�����������w!�C ��A�)��$�������M���r|օ�����$;��r�Tb�X��T�NM�������*SY�q��R:��y����r fR(�^��f���N�I_j��8�t�Mܳ���l�W��'_
�4�L>?��H�D��d|�q����j�x�D:#��n��O��7��G]3������h��\��� ���hߊ�w��߅��Vk{���8����t:��P̖:�����p�1*��{~/¬�^
6���~�x�k�_�*�W	t������8[W�5�#���P�Wrɠ�hz��5l1��!�����5�L�4Bx���@���_�-������utt�����6���W`Ǚ��N��m���/ʈu�"��w���{�qGY����(��5���	t�P[[�ُ���7����$�݅��,T�j����3:�y�ϡ}�T*���hze� ��e
q�_F��
�?�����cM$�g@���۞F�	E����"��4ub�*&V�S�ӯ��4���m0$�=ķ��yr��ҩ�nuZ���;c�ʟ%q l1�[,*�A�d2��Q]$�݅�{��W�����p�B���-�(g�\~k(j�O蛾��;�g"��4�Q]��ŷ�(b�z�Jm��k�F�bg�Ey�u�4i�`$]�g���7�}�F����~��ӳ�Qa ��*4�	��D�_���>�jeX��P��45�?6�ޯ�cA]��3fl^�f��#��WJ���2m�ڃT���p߮M�)�^*�Q�H$�x<~?����R�?!*Ɣ���k��҆g��m�ym��ڒ�dgX����y��Mظq�\�3q�>m䣎F�U����G�r�rD���(+V���b����S_aJ���Îާ��v���h��L�{���x��!�����s�O�F�M�)(�;;;ی(�x<>��4��eg�N�����>�[�lQpc��i���h5C�1�Aѕ_|�m�11�Z
v+0���hzY����}}}���8���/�6+��5n�E�Δ�*Nrq��3�~���jW����6	n�6��4G��3b�Чa�DQ��b#��
�j���Xe|*�9�͵2�D���w�2�n+�K�{M�H�>���4���pm7@�?��槙L�i5�W����7�Pm���w7Ƃ.�Ʊ����3R�h3�u���vF����8���Z26�%'����]�.�>\�U&`�s���N�3|n���vH�ޅ�x��W4�,L�}	�����h�b��C����!J�U
B�K�)�k��߷���i'q�'O��Y�r���T\��Y�f���E���Nv1�d5֗U$}8x$�E�����W�4�Vƍ�=Ye�|��s��{E�+Bl!�υ�z�{a�i��/藙~@�߆���^����Ox�^^��}#�ӦM[+��(ʛ�����h4z^����Z��b#����`�p�{�	t�mWL@���آH�z�b2����:C�ȹ���aצk�)+\��-��e��h�T*p�(+���k�)��R�Tsk]N��[�_C��ioo�`�/�wZQ�qG�����p5�_^�o�t�mtpٕ	�"�N����u}�� `�q �L/�;�[�㿣�Q��bg5���#�һ���@�X\�����?�����bз>������D6m��8���ƿ[{Kb;x0R����}�)�Q�O��� 6;T������&�H�{q���_h�`;7���P�CGĦ�A�\ؕ��W�z	���Yggg`2{�{$��;q�ӈP��Ҳ�֭[�D����B�"��e5#��&=�~�2@$нo�@	�Jbg�%���+�+5�#��W48�WA��b��9������3h�!Dhhll�T__�i��M��M1����jf�	1�H���m�֔�vT���fC�Q0P��8��xq4]�ǟD��N;����ի7!D�H$����1h�D�±������+�O*u;b��Z� "��1���+��U]E q\��r��W�]� ���^���i�������#��%x���<�E�is��8�����lÐ��ߘ���c����b��y�cB�S��M������l�_�oq�_�r��SA��*D�hll�=����X��O��FTE�E)�Q��׸�	tR[[{n:	�1"q.M�,rl!��l<�#����^�L&Y�;�%�H4����g�)�G�/�kk%�����-��^�H�wuu=k�z����r,{�1*��D�t�S��鲟`M.�A�����x^�uttt!DYq�&ߟ���18�8�h�gP�\�'zlḀ�$�������%�G�M3��F��}kj�����@��}+�>������FQ2�{C���ah	?b���ނ�r(��Èr���PЧ-1F=�G������وaH��*����1���W#��np�u
�e���N��o!Ĩ0B�gg_4����C�G�ύ����J@����/��Y�J�V� #��Q����a�ͅF��s1vm:g����^꾎�����U���r|��f2�UF���J��x|�Cpzx4=��ny?7»���0�X%D%�O�{�"=H�Y��	8R9���	���#Q!1t���J�t_C��-����;�����7ΗC�<�ז�R����	A�Dcoo�Gp�������WV���B�E�(���	� ��?`��)�pL�F�,#7�<��`צs@R4=L�8�<M��C��<�+��
��?uww�B;g��!��͛�q�F֝�8��As���]��>F���6�W� ��}���iB�])-L��k�E��	v�)N�D�ѷ)�)���
�T*���c�>e%��p����@��̓m�i�?����P��[1���'�G�'�1ϥ��_�j���`���E&�P�O��,Q<�x�ص���K�]`��;?�:&Bo��<^{����_�y�_nmmՌ��---Sz{{�C�s�#�)��1C[L8�p�kW��bo9�})�r,��ؿ�\�.�����K�����{oQCC�)fh��P!q.܀�����"4L����H��>غuk�=�SV�?{����d2�ʀ<+1N�ϟY�n�^ds!B����r���<u�^��~j�O!���]���Ϙ� ��0���/��y�	���-��Z�j8�����̬�F� ܹ��U�ƪ���+3g�l[�b��s�{���#�HK]]�^�W>�{e��}Vo#��B�oe��KM��@�	�d�����BI��B��s!��F�{{{M�L�}�c��+k֬�po�)�~[����~�⽭��+��t������nN�����n�9ƥ�L6+�%ą��`ܽ���g�	�>����l����� �"��p�Vz��t1
,��!Ƕ	2��h4��ށ�6�v�6x���X�z�F#<��9sf�����f�Z:,�6~Lk�w9�I�!D�@��t:�؄	t�������7�fh���AqΪ�BT
�I�&F�Q�H���ս��l�ۼ� �7�^JC�u��	��9�M
��7�p�D"ѐ��f�9�����L3T���,�Fy���.���;��~!��j�>#�L>�~n�M��8Ղvm����E&C �b�>����6D<�Y������k�p������h����{c�ĉ��g�{��ٻ�Z| �^����#�����x���"|׼�k�B�
�|�R�-�>dʔ)�nܸ�`4?j���E�Q4]T	v|QǶmE��%'�x:Qy����6��F���p����m����{�����-�=�|���l#�;��d�χ`�'F�>�x���˃˱��4�g��)8��y����2ǩx��Sx4C����F�m_{�h���B��S��S&�H����+Wr��	h.�5�C��g�[��q�h9�W~�(M��J{e�ٮI~�=ɏسm�?�!2ҽ��L ��E2F�}�熿�V���o�}^�1�o���B!�	Ɔ2�̷L��@�)�T*G�(��������:iL-�)���I�b��{
F,��.B�#�BT�e'N<c �;�H��������q�����F�rEr����B!���X__Bkkk����@�9�d�O�'Bh=f��2
!�B!�_x-���ֶ�	�  ���X,�)4)ҧ!�B!��>+����M�R���>�7���x�����_��=_�B!�«�����s�1��؆z�H&�+��!�l��8��!�B!��x��4�9�z�hoo�3g�G{{{���F!�B!��U�6�N_�j텐@ �W��XSSsr4]����&!�B!���\.wj&�YnDA$�����Y7����h>���F!�B!*��$gB��iĨH��d2����q�H$r	N/3��!�B!*C�����8D�$�C@OO�555�WWWw����B!�B��/�)t�?��iE͋@=Dd2�U555�@���ӫОm�B!��=���r�@{�و��@Nj���K ���	�}�B!�B�h���W���g�7�!����!<HC�����q�#�B!�c���Q��J�^0�d$�C�#��͚5k����S�f
���!�B!F�9�=}}}�����5�5$��6���^�aQMM��MMM��xΏ��5B!�B����Lc�ΩT�Ո� �.��D��I$����G�u������M4B!�B� ��U��A,���]Q��eG]�����s� jfΜ�D"{A�Ӛ��T��G�ў�b�B!�^#�}#|�Mho�q3�o@���r���g�A��7�*H���q*�w:�#�B!��d$ЅB!�B �.�B!�Bx��7w���-�d    IEND�B`�PK
     Ps�[��C�I  I  /   images/627fe4d2-0152-4b97-938d-4b9176d7a483.png�PNG

   IHDR   d   S   i��A   	pHYs  A  Ak!T�   tEXtSoftware www.inkscape.org��<  �IDATx���U�u��0<��y#�W|E�b�M�5V��6�������Sc�hMl�1I�G���51jbk5IU���F06A"UE�	�0�83�c�a�������s�=�{��~]߷�{�9���^{=����7`��ɦ��ǿT+8Qp���
{w򅱬��1���z�B��O?$8=����8��}����8<�}�1A��'�s�ۥ��r����C���O��ÇM�~��._�
��54���u~www�D�
t����wK 8�Np�`�`���"�>����0�mۛ�~�3v�	�_���r�u��R��3\�g&�@]]������_9��Ѓf!=j|I�E�u��	6K��%��� 8Dp��$�Y��
��#86���F�7hР�8y'΁�	絋��'�U������uMxQ�Cͤ���ꊈ4��^&���1v���C[��@�[p��s�fm �s��y���f������Q;!�rK`\ ���͡C���&�ǂ�'k�ȭi���y���}������g"
� b����|Bp�I�?f�l-8��C�S���b��竂���/c�}�������L�7��O�3����\�`~����N�jC��+��rD��$��f�w�Q�gq��H�~k7v�R���XL�so0V� �]�q��e�o��]"ߗ
�zX	��~0�&}� �q��'�5�S�52+AJ
�`���r`~'E	hY�d��'�%����K��p!�"���D�(��?%�Y�q>#���%�	����-HDc��S�uttDc�Qv���� ���@2�<��Cs0$
���*��4n�\�P����N�/����
n�5c�!S� !�pH}���6?%���|�Up�_X��0�>1�eT�;�H��~�=dȐh��L@�3�>�`���zfWða�v�{�ƍ�˭Ok�1��36g� T;�T�4�*�E�{�7+��J���I?�I�����	��P�R��*���ݣG��b^-?뛛�omii�$�8/�3�˂�͏$.��#��0�,�	�A�@����1��O��q 1mY�bOVE<��t�҆�����,!�b�U���ۯ*c��D�@�Ϗ)S��-[��k��Mu���Qx��#��F��!��\Ey�T%��BL��|�c`�|�-�lr��?'��`S�=q�����8S���/�D�rW
�,�wq�)�,P�X��3���X/�{3�A��1.4�X}B�,Vtm۶M�Yp��%t�.�r"R-(��_�Q~�+x\X^��<P��`��:{`mt�n�{���}F� -��3�}�TF�Ǔn̛7���է�P7jԨ�{������v�?q0|�y�*�!��|�`��=\�x�9�����C)f0��0I��X ?�/,X������4�]xekk��q^����	FO�
A�4�� �#� �ϭ��"�������3g�M�6�nz�f��Y�S����2nܸ!��A�뽂��b�e�p���-�8DT���4�'YEWE�E�#0��&oV����� ��9�FP��E�������f":��y��k@Q��B,B|��	��o֊�F9��]$U�*���lM����O�� ��ޒRn{���Ks>|�� %Q���o�䎎�C2����P����a�cC�K�^�UAQE,�G�����8P-��a��w��%�MNb<.3|�����4����|�'�\&�xF��V�>*�*�����ͥ�^�+
��x������5/��r���2p�0�	�qG�2{�V*��	&���/��M4�ս�bM	w|9�
��]�W��`�/�ҠAtQ�a�k{<�%�@TUCo��"��]�n�{�tV�E,(O�M����E�"!J�z�!,(�����2T���@���I�,�K
����MG�	��̾��ZU�����<y���s�obz�9��2]@��Sf��?��}�m߾�O�/���Z"��j���Cc�"�M��IVWn�0�@l0VnF�=��E���Y�_"��&a�4'\&��W���{�d o�s�|��Y��_��kiiQ�L?N��FV �&V3�׋IAH�J����������H/"�;Y�F13��<���2�mӦMC���"�f�PF����i��7���755�?Q��h'�z�޿���5�d��l�^}����I�&�k�@8B^�7�����X�a!s��':�h���뎝;w*q�ٻf�?� z�5� [��o7v�J�J���_�=����4��x�c�E�Z*�#�r����666�'��Ῐ�7����`�}2�|3�:�g��S� �6���g)a12+a�?2v-39O蜥^�~UpP����o׆�5 �I�f���} �����}���YwY@	��TWI}ɵ32V5��D�"��s�<?!$@�Θ`�L:�b�]�
!��P��X�gJH�~)&�_�㵒L�
�hӀ4 ,�>�4�n^������[u�@�_�%��,j��9�L�:��͛7�Q6����e��@���u���* i�������U��"!� �K�ڵ�T 
��M�6��-�2��.�p	6:��mG�9GO0vB�O*�� *C��]xX�p�8l���w�c�-�e���r�D��1�|f��*��f�	
W]ƿ���������zIN�GB�y��+���lv�X��&�yR������$3�*��s?ق�Gj���M��a,�l;׸��N��!T6�X+���ٕ�^�QD
��B.�����^��!$����;�i!��g���A������L�X�%+����E�(�=�P�̒�r�X�&�B�u�$�����Դ_���ls샆�p�Dd|b�D1��������OV���9��e���ث�Ʀp��
ΪnY`�M`b�56-	O���'��� A����J�"	�Q-B��!q)DY#ˍe���fo�����I��!��W8C��VWlJT�t��y������-��
��Xfv'$B�c������u�<"qr�=���[$�r�b2�rc��z���"�M���2y�VT�9��6lX���w�G��39 JL3f�Y�zu���YZ]Ie�z��s��5���2�{SA;����BC�i����on�ԩSu	7�ayCB���Ŧ �HWID�rVqf}�A�ys�M^����S���	10]��1�F���PF��ɚ	Y���M-G�V$�j��B�e�Tͼ�{V%�� B�g8d;��4����J"�qH8(Z�цH�5G�� W������<�C��è�<;$�#H��ˍ=���IKͱ�]�:��fAG�śBd������@D���At��'v�9��~���o���Y��_0v� �.�"��W�c��Gc��Z�`�w��!��,��+�� ';˅,B8�M1�).)����f_ɇ����g�!i���K��'	 �r�o�W���dEh�D� Ib�ƾ�c	�{*�8��������z\�����i7��3?cB�`��=����I@�P̕����$e�j�%��"Z�LG�,.S���+zJ�b�F�Sɣ�Fp@1�m.F��9J�am1��r��$9`a@�����⸩���z^��֮]۫`@�\���lm^@��s���M�ِE�[ӀX�g�+T� g��������c�ql�z�?��=�q�6`�)�ω�`��z�^�\�5�ё��Ϧ�%����EB62�l�o�z�8����n�EI������VnWR/���*�������ȭwĈ��N��UQ�ó����*�JJ��Y͌�L����E9bx��:2��,"�p�}��� ±y�L��o��� �X��E��PS9�TM��ⴂE	5ֻٰ�.�R�ܪ�r�#����p.����~z����:t�۷o%��XeX1i&9��F�'nӏ;��	�ۄ�?[I��ِlV:.�`Q���XXQ��q�)�DIN<�%-71<?dȐ�tvv;R����V��B!���0駶8�a��O����y\�	v
<��p%�C{4_�L�Ę;wn�\FQ#F�@��r[Ȇ|�7�#577�ٳgG�ۺu���A�e�g�X������\�2~�x�6�Z)�9�\c�_�(��L��L�� ����u�dV���;�q�t�4���K����E��q�~�)�&�Q���!�3�Mr�����w�!)w�1��fp��?	@R::r����>��� b���e����(Z�9g�+���,�P�F��q��utJ��8�m���vD�s!�ľ�^*�C�Y�'Z�.ܒ9�FS�@�Q	!7A�%Rcu�礡rއ� f>J�"��H��y XE*ǲ����y�G�<�_�7�\c<x��H��F�]?hР�ك��I�
�V��0�Yed�K�"��t�*�@t�e��G��'��=R��]r�V���+����l�C�� v��p�"�\l��U������Q�w7:nY���K(�3^X��&8�w��{R��)XR�]"�Q>Sk���o ��Y�����d=�"~�w�H���/w655�����Fyk�u���!�*�`�$(���<sD��$Q�,i"xL��+��2T���J	�?K/-�1��	��lժU*�XGG�ÊA�����-_4V���`�RVO�. �"�a�g<)��G���{!
l}���M/R�3�B@�UI��u���� K�;` ����9;�0�~L��K� �〔����}��n����5����!r�r������Y͌#
�������ߩ����J��(�/1BQU�KJI*rgk��yԨ�!]]}䎞���<Y��5v��PI��`;3��2���pPduA���2����E8�pv�=GV�e��ұ�*͓�r#J�����ڶ��/��/j��o +F'N�Â��ޒ���t�ia�� 9�!�� )����刣=@y�Z��=��v3�>�_*3�N�eVF�hA5|�BHƜ1N�a�EoE8��g�k83Ɣ�7���[]��_�>X���o{^`v�t���]I�>�Cp`��Nu�ݙ��4���	�Ń߰{�nD��~%pF�7�a̱�鐾Lk����+����~B�|Ѓ�P�QP����]�CX3��y�$��ve���YQ�:�Y&P�~A��1>���K�3@��Uro�|_V�����!�Dx��%����d����55�B�ڤwM%3��B��*��]��v:��ń���th��)� 'e9�&��{D�%��,�*�G� 7�����zC�I_�]*�Dw�9|��Ƭ�x���Ms��Ɖ��W/����4
1Ȓ��݄(�<ĩB��;d9����b���d�x�4�����m۶�<s�̗:::NOz=�B���LT"�h2�<�?��pa���p���`89�>wn�K�"�-q�!�sF������b�8��C�Nj;v�g�3N�ed���a�{GD�bq�a�{��:��}R���#}J<�(y:����Mc�B���:b��$	;�#C�Pw����j��A�gI�G��&�,�mH�ަ�B
E7���I�
�����I(%X��g$��i��i@p�/�!�p�W�=���1���u�&�����m�__`9A��)�:�����jڪ���C�ꦯ~J{�E&O]de����=�S���eM�3{�}M����Ʀ���nu�(#�&����� ! i?��ܻ�y$���#t���ߥ��qqi'(�e���{�[�|��;�3G_&pyJ�ǩk�����U�Y����u ����+4
]�Hð��`q
{F9�]��}�ɞ�"�(L\�
����?g%�9�¯�K�T�Ǝ��w�� l}�t�H)���l��kG�v,i"��G؃��w8��>���$LF�~��#Jc7���r�.A�ϥ/݌���PPV���KAB=�_�%�+T����Z�n�,�rѓ���1�6�Db��2��GXRE$�e��Z��:�5��:Y�_�K�����}�Gd�b�"�������,�P٪��M Xn�C�9~A�<J���z^:���ۢ	��~�_ �p�,4eN��3�}��}ǔer��C�<A��GD��x!z�Nk��HE`��3o�8�4�M ���A��_��k�=d�8"%sB�[pT��?O�@g ��o�3���.8�b�W    IEND�B`�PK
     Ps�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     Ps�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     Ps�[y�E�wf  wf  /   images/6a97e33c-aa93-4e7b-a2bd-349ce97096b8.png�PNG

   IHDR   �  F   p���   gAMA  ���a   	pHYs  �  ��o�d  fIDATx���$Gu �Yտ��;��_��h@B^K6Z/,��5�kV�فY;���]�y��v�5�#��Y����#�3�1����ŀ�Ќf4�;����wNf���Y��u��͖�{�;�]]]u*������4M�.���»��w_y��u׽���s��������x�Ew���}���p���ַ��iz=|��݇���n j�ZI�Z��j�^Ǎ+/�:�����B;M���ןh_�|yV�i��s�#G��776k������4M��2M��w:x�6�-�;�n�^�uV�^m4f�V�U۷�����Z9t�P��g��;v,�|�觉�{���Z��j��v{f�����=�	�9�g����gT&y��?�����ŋ�k6�1�,LZ3�������0�})%Nf
��q�$��s⤟����l��R��2�	�ŕ��Oәn��DR6R){�^���5�q΅ߧ@02IE�_����~%I������Z�����S���N��7;;�N �.�ܢ��u�LT���ʝ�c-�{�6���\G�/^Z�i4�ϝ;7S�Vڽ^���v{@45$V�7�q(�D
~i/������+W���z��7�o\�|y/~^[^��l�;{�
x&���5.�@�)�]�S��
ު�ʁ6����w�Fc�Ա'����|�O��O
=�A���_��߸��V�y�ٳ�^���z`e�j��

�֫�w�u��5�i���w`��p��$�o&J�I��4�Tb��^�Սp��}T�<���p~/����P�Gq7�Q�6��Q5����40�~��4[����LOQW���� 7�� u���$< 6�!a$q	�q
�q� ���@Ը����:��o`� ᩇ�i%�['���U:�"`\Ҵ��_K��"A�&��Ե�H��Z��k�{�����0V�X(ݙ��gN�^k4g_�җ�טi|ҥ}�C�#�8ѽ�-oy�3g����v������0 {�+$*�J�Z	j%�q�#���`<�=8p0��S�<|_U���f ��	�Qǡ�!9�� �F �P���J���x�00��&a��yUZG*��`z��� ~��W�k��/��7D�pC��1I��(�
$� ��E"�W���J�d)��h�g��U"���и�\�<�++pFgcc�0��0�=���������޽{/�|��馛���w����M;Bt��{�O��<��-���Hp���`�" 0$3�b5� V��c���CM,���Us�=��z��t�?�'X]�@U��(��jH��`F��_�H	/u_M�2����F���ϧ�K�ϕ.t���;~�����{�׌=>]K�{�� �T��$IWVV�<uann�Ү��Ξ={������뮻����o��o���F���/��˿��/�H� �&@�$ = �X��T��%���@�s����5Ԩ��s0So';�c�9� �a��)�ǿf�,�Y�h�M���$5}C,���mRM��3�jbx��S�vΏ�3րs���7=��Ր��F=�z���w��y0�?���7����=�z��^��WW�>�g��'क#��~������6��w�}�;}��̀�IPTo����%Џf��P���p�JF`��p�@���5ǉh�H M($�M��(�+�i�稱��Ĺ���{-�������^�:i��El�Ζ�z��O�_j��
�0�k�_�� ?=ϝ�K�w���M��0�:�z�%�O�Y��i\e{����n����/�gQ�Dtw�u�O��t���捰"^ v`nn� � U���J�]60��K��lv�&���4���!�U� �Ԉ7}�t��4AH�:x.
�D���Zl��s�QDƮ�����=�9F:ft?)�n%��b�+.���х���O}F5��d�ÁJ5�sunmm�`�Ӿe~Ϟ+����`$ѽ�o�Y����u=���p9Z���P
��Pv�9D�K����
�EJG���>:�TH��.Q�{�	����T��Fzri���پn��YxO~��=@u �lŹ���j��ΘSW���I�"J/���*T��鈍��ƹ���[��D�����S�N�n�o�b�n$)לȊ'�%8:	��:��ʯ���)�4�Lf���	�}o���Q���G�����5}cDWe ��[R_�@��?ķ�.���q���	/��.�uUb�I����}�Itp�6�f3���	�����⌠w$��L�$1�]���ƥ�^>�p@�ޭ��;�!�h;Y�X_��zoti��g��!�j]�����b0�耫��������_��6�΋U.��hM�^�1&�.(�D���c'z�I���?Q0���ɧ'�W�����T��K�_Wd�&R���DlFF �`h�[MY]�G�?����t�����H�'���E>�!�&��@n�"=N/dr�h�DWI%I,��,Y�V��e�z�R��[��H��Pm��+�\������*��<�&�����?1@i�g9�����I{��E\z�s"tH�
 �6�
��퀚�v�k#�*�([��D733�Î@�v :DV�>��~�=(Y�����}"3n�W���Iٟl�/��B*��D��R���1̀��&��8I�j��;3,���`VMm+�ItgϞm�Z�
�1�0��e\�[�yg�u� a6���f�U_��t�\���sj��<|w���%����D�JB#H{�Z 5�J#e��3mvڵ�׮T�'�՝��?{��uʈW�L�Hp�M����b	����z�vGY��6A'1�(� �P��L�.�����|v����Xe�M��(z{��Z�}�ێ�H�K�/QDח�z�[�+bqv�t�a�@m�H1¨v��(
��5�n�n����0rˋ�T�����s��b��3O����X���1i�u��ư��u��Q#��D<�ƵJ')m��$: 4L��R�����V�e?`Z�����|i�����[�2���Ax\� 'S�+�y��F���V,XZv�Q#�!̜� �K[���Օ�����t 
}����Y�Pd��@��E��i$�onkg���D*���8����I_bD�
��H�g�QH1N��S�^ܽ�����hF��R 8=[@}���Q)=(#��СCկ}�k�ڍ٫�ȹ�Ӑ� r6�?;�n)�Ȅ�IDƣ��*��������}�O���4�Z���PMڪ��'�H�H����bd�V��Fm���F݅�_��ׁܫ�1�7�j?�z�l��6W������\/7ƞ�T"�ɞK�-�{y�{��ó��+��K��viӸL����t�$V��48�U\$o�o(�ǝ\F�FG}'�p�Z��A|θ��0�M�*:o�b�`Q8�@t=��f�^^]�E�ٲ�It�Ν��j�>^����Պ3>6�a≉�
�2�Ȃ6�;��/r��7�=B�I���aQ�r7�C7L�'��nRM�\�������j+LaNM�&Cpk\��'V��
R����2��|�ħ3G|g���q@"��0\o+�M���+�\?/��q��r���LsؖQ��,�#�ncc3K�X�J�y�v3q�|/D��Q ���T2�����5D��Р�N�g\+��Dq�6Lo�a��M�*PGHC��0N�QD�U���B #Mf�J��I<����z9���)l�(#���v��$#��F<�a�Oy�=c�H��YD�E��9�o˒�L^]��O2$[�뙯1�(���veq/�ĉ���v�nEc���m(�C�7���%1�y�s�!���x���#����b������#Lj��(�t}���L�8��"��8�$���9���ZБ����� �L�sa>k�-#8��1'(o˻&	�Ļm�cz'8������j�����<ݢ�d��O��{�[:ӤLDS���:��H��ԉ"�c��)Z���ȄO5��9��A�S���&Tv�m�!��ᰥ��N j�P21p;�ME"׌z��R�1>�����t���t��%
���TۋY��6�Ќj�`8r1Sȟ�CR";���~�[��#>�۩�)2 �N��1*im�����۾�W#CA
#�K���D�*�lh�N{�Ww�،���aR!� WR��������D�\A�{�1 #�A�v�7rtڹ.��+ZQ�ж���x�J���� e^o�j*�!.g	��l�p��g�`�C�gj�U��S���o��(�R�"��+EP�#n3Ђ6�'�F.�\Wf.S�U]]]�!����m�Ca���%�!"!s���2֬�*��Ǉ��Əb�ONJ�vXN��P��&H�ɡ�i��6~:���xFX�b�Z�u>��%���ە.CIt`<`aN]'x#mHD,C81b�>[s~Ce�D��%f'����鬈��]ũ5*���b���dVD�c��U̭J�.�9�9�t�?$>�^���mM���백$��\|I���`H�ɵ���Tf�҈X�J8R���@}t���W)�=�d�$���uӰ���u
.=f�}r��p�m	�YڪA4:ʠ�������tIj#�ȘƗ�y�ҥ&v�ƃ��J��	 Sn;K3�4U�Wd��j�G�Lٓ�w�Y�)��:j��`|HX�v��8�����,��x5w,'��b�䱦���E�2�~f�ũ��?�Q�U\5bė�C�Q\�Z�(�1���Ȍɝ����?5�PtF:�WC�^I���`M���o����M^L�h�������{�OW�2��>MH��ٜ��en1�g$�����������&V�������3C�/�A�aRO	��,9��X"<�Y�d�K�ѳ�v-�w���u��гkkk�^���Ux#��`|��N\�}�^��Hq�v��hO�V��g���Y�~G)��`$����mCl�$��ѳ�-�gY��p �_��
�T"г� �}��^¿�͍��%q���$�k�IW׷�*%�>Df-���v���^��)�|��*�� ��iG�c��_4��Ū3\��(�B�Q)��v���ȉ�U���}�� ���O�;x�`��O|;��Z�,Ҫ$a`�+������j���pSZuB�d\qόXŀ{�,pv��m�&��X�M�7�~,qS_L*�mG���B��5�Wl�l61uE�K2d��)\ǰ��hc��&ĥ��WT��D���BW��5#Ӱe��%5Fr�!"������S�����?�!lL'��j��:�������A�g����%�E��!Rk@`/$8�	*�;�V9���5w�F[��t�P�n�C!Ks���U�&+�қ��o]�|_��X7�J|��ۅ�)A��.�Eō�r�(OM���HU>7�*�-)ɺE
�r�?�^������.������)�o|v�I|����t0�N1���h��u��o�@������~�Τ`�.�m��Ս�X#r�<�r��C]�,,	e��1met��~ZӖ�mc�S����e(8,^=y$��Pg�h^�Kx�)0�6%j��.��_� T�F�4(K�����`@(Z뙟��8��͋x���Km����OG�Ex�G&�]�+�8�}L�n� ��~0�
�TI�oYdZ���D���VI���lun�'K�l�Փ�x�djBX��F?�!�\ ���d��F e��_l�$[ȭ�`�>�y��������z���؂;�Q��V�M\���RZ�����%z��y�1�W��
�=�r�2 �1Q�ִ�f72�¨i��j�{*�t�Na ���tm��={s�fI4���v������l9�G�RS�&��@n*vE� ���r�m����Bt=�jY���P�Zej$�>�];V&�� ��gb�/�|�\-����s��݅Щ��0���&�t��.�i���z����
���x4��+gd�}�4C/#��������Ms4��v�*�t.��IgwA�>��D��Wz��iu��iY�E8DF���\��J$�1H���1��%�� ����m<#)��yqY���ӵ1āш-�K��+�����Xo���U-j1�G̐�R� �V��c�Tz�$P2Z��8v�e{�b3�'2C!5�*�> Q\�������/?�чG�6��?^_^^�ln6g�T��Vgc�gx����J$����wMa�$���p�D�'Y���&6c��	������la������;#&ӌ�ȋ�����{m��.�2�0��.^���u{1 ,us�����	�����'*�	�l�R
t
�~��!)�.5���)���m�7�F�G1�"�7r�r�H�e�<�K��{�����?r�'G]�L���nw��Ɯ��D�Iu��=D��y�j�T��o�D����}�4:�Ό��|�����~����3e�0�^�U"���|��^(���ոT��ȓ67[=��P�[�waJ�$�'x��}��q*�&ոjS�����l	���9fӟ���4p��H��)����[�FX�7�ֿ
t�v�n���!�Z�^�ln*�o����>��|+\�D��-"U9���0�7w���fk��w/�Y����S�٨������ghI�d'$(��z)�=��VW�v�(�#ޘq�nuf�^�b^ ��`�=|�]=e�R����yO�Jt�u���*A�~�����D�ͥ)k��԰z����j���4f�^�_�R
W�#�D!%WC~�W�i�%n)�>b��;D�+Mp��h��#9�F�E�c\��(����(vi)_])lZ�J���OAZp̃���3g�͓�>��pv}��2��9��]��C���de�q��_��r=����EtJ-JgZ�V���设 ��Nb���$�Bj�J�u %��D�b��8/U�U��`R\N=I�E�� ?����
N	"+҉L{65�[�4q�-\}���q7�N��)�D��N��Ctڭ�,vⴹm�|a$O������D�-��Δ:r��9X�.V���z�(���Az�&�0<�^ƅ2��*0���Z}<�Dk��1Q�I�&2�
hJp9�:Fj�~Sjyύ���@).�7α"��h<i��D_^�朮l����3�&������\��ã��*�.�l�����1�y��6��xLUq��1��N*cb$�$�qo_}����+x\�u;��n9H���L�Q�m�V�Tw!+l�?WmԺe�S�FB&�u�/�IO��r[9��b?Q��1����h��L�K��{5xM�WpH���p0J�iN���I�!�0v��˨�no�;�Ra#���ի3�t�f�H��BjOl����>&��7�h(՗�pW)l��,��<q?�H�K	μ�N�z<�R�wwC�F� [$V��+R%�@�s���st��J����5ja�X��fH�b ��梓7���2#,Kx���Y�+8 P>���E�E�oX�7,�5�_*3�:�nw<�ncc�(��Nw6�{r
"�b�3�����6�Ė�^��Y���^�;	�II�tU׆E66��*]�=�Y ��A hR�hJ�%Q�9܆�R�y[�P��,^E�����Lt�=#>�AJ���v'���ƶ�5�Y�[p�3�7��J�f" ���j-QfD�E�^�q�(�,��Q��I��
�!�&<��@pY��SA^ `/��������ER��������ܮ�J�SN�	��/�)\�.��j	(�V����e��y�t�..�)6�CJa�Am%�/��9��=�Y�+8dIt��./Y+�,(�7�k�$Xp��'�w���ŋ��(q��$|�N� =��d�bh&�������\*
�}�n"��N��3�X6p=*�Ѫ�t�b@l�� �g"���Q137;N�j�ڸW �G�N�����fz�@��w��F�IJ�6e�Op!�����T�8D00I�)Y���j�ۨU����H���Ϋ�J\o<���h���j��t�T�����D�b@].���CPP:Ͳ�7��-�]+uh���K�<NH3�r����VvJ9�J%�XZ�6�I�Q'Y��N�N�	p�H����������{��kuݾ*I�lvv�E$k�j>g ف�cx����G|����T�9ʜ��xo���=�Fa�H��Z-�0�薖�jgϞU5�����
a�^��S��D��j���:AH�T���q��-�r;,��\׳����4�M�hid�NG��:��F%Ե�o�ϔb<�,�.��g��fv	����m���2Gcv�ъS�n�?c N#�;u��[��e�!���H�O�&䎢�&)���{q�A�A-+:�v�R(��p{U��t�jHM�(��	Ք�)%Ԓ"�¨DZn�|�7�����dy.�\X�,��9�qF�P~:�0vK�Qo�+�}o}u�~o<a0�n@s]�dx�ݲ"
�5�~�i�%T��;�2�x�=hٍ�؎�H$@��\o_Ҫ��Ff6���U�F��Z�@G$�<F�e<t�A��MiK*� ��i�$�2��)��JA�DJÁ?ꆩjs�͔����4�5�q����G���*��Ԍ����_���?�;���e�{X֪@�Y�JԁYO���O?��֞����
�3��xvV�il��l�d(�-��O2=Ќ���6�1g� G8�j���Y��q��F&�IY�Ҵ�%|¥%��b��ʧ�ɏe4S����2~�����3�����uWwzo���e��(B{̂+~h�cR״.M�o�,%�d�7&n!
.U�(0r��V�F�!箭�ۂC�����:���9�$��^w�|=^#2�R�$�ӣn�O���t:q�^oa'5ED�z@���	�j��1i�^j;u�'����ݮ��7�̩r�	N7 ʾ/��	n�h��QY�qH�;����r��k�������y��q8�>��@p	s��+ �I���e_B��W��=������R��ˮf��&��?5[P2<�P��F��b����5��uٱ���Ոl�PHT����Q��@4U�=Uп���cQF����M`͋�6SvV�L2� ��H�J2��"x���P�l�����lQ�&c��>4�}(�bi�^{;\���h�_9�����-�D,]+1M}9���m��^~*~.e�8C�Z��h	l�Z�2۴Qv�gx�� e�a�0z^�ʮ��Z2,2��Y�b�W�څP��7q���Z�Y1-i�����(��C@��ɠH��e2�|=��d\a���yt����T�������3qK�'h�F�Z%�a�գ�3���ܕ�HSɉ*5{`ۓEf�\��Z@x���[đ��v�;�6���t�Ό%�f����	eD��sS����P�v��μ(��k�ہ�רZ<��D%{5�Ð�F«�З�Ŵ@
�Т�zfХ��M���O��t�m����d�k��\B�
O�#mD��������Hl�4�O3&-��֣	�^��T�5a�
æ(���n��h4z�v[��|�P�ˍ ��~�F�Pb��x����a��8A�n����)$.�a"U8�=i�{IFt��ۓ�ad�!��RȾ��M�5L؃ �+��ҭع��N�e6���Y�`�O�Y��ki�ط���Ua��1L������ԎX�j���z�d���ԐH%��P��t8�u�xٌ���*���"Dp�<SJϓq�QnW��$�G0�����2n�Y����u^��W��ӟ��g���L�I��l��J�\/��Lս[�8�El^7s�"��g�pQ{5�7"Fi���9�c�&'����c�(I��641e^I�����Ws��N�E�|�[u�ѝ臙hTR�0
Te���`�D�"�ޟ��?'�!Q�+��T I;�MI�cuE3dtխ	;g�L:��S �/%�K�#MZ��پ"n�B|����G	pd�CjL�K��xZS��2��<=,�$m���L@�/1��N��*���\�>���S���Ώ�菾�/��/>>lx�]euu���M��]��vl��I�x9#��5�h��R�R�'J�twKM¡]��R��HjZ�����������Rl![��,<ÇC$��đ��D⓴8�b�>'$�)���X�q,��%E�׹�`ۉy�-2&�Sb�I0�i��Y�l�Gn�T��k�_2�q�T��2�ӕ��U���Ա�2P��b�䬛"�pH����Nol�ݝ�?�`�d������p�N���o��&|�U̳I���&��,~�}�tMIO��i�从z�H��;���P8�J�U��)�f�
�2�N���1֏��]��[��ӕ�1�z��i�7�ӫ+��OdF��S-�`VVVD��U�+�jcB'�	��ƹ�4Ħ��f���u��������'�D�L_�����<��2M��s������)�D��JZp�`S�bh1��򢊽��f�J�e���	45yvH�rq��Ez7	�Kj�J�u��D��O����%�b�')��2Du>W$Z���(�r�#677u��Z��*�4y��D�%	#so��&�b��������1
��Fy�ӡ��\��U��hg��-e��b�(+<"-sk;�$����j���~R�Ȼ�&Mr�1��{�k�j��8:���>;��C\\UI�4x���HQ�ȤD��D�b��*�v�vYh�0���"�AQ�jobe����>�[ �)Q�5T�R�L~��'�����b�Y�q@H	�Z�E�d�7�%���ЋF�Yf��vb�/*��M�$ʈS=�yeY$�����g-Sn 9 3�.b��3D�%��;�)�*m��v:m���0q�9�4-y�s�$�\1&y�W�V���#��ʕ+	�rL�T<�C���HZ�)�k]���D����|:��j�3�V�+B[[[3i뚋����Hq>�����I�N��O/
���ˈ
�.�7���.�!��3Nx�6���l��7
��[t��"��e��v"��84�(W6�Wh�D�qϞ�����+�ȅ�ǎ��*������M_��z�jgj=
��O�}�\"�T��l^;�ۻwo���^�x[���Қ��������;�<�ضI�Á�ՠ���Z�. �S�V�PY�T����v;� f"�%B�%�i�2{%VQ����l#7)��+��UX:�f\>���\�\8B�[���,u8��!s}ې_�F��x+\e�h�"���5N�u���Aq78���ӈ��m�T9��l�6�G�]m��&�V����u�	� �m@n�n����AWr���USyԳ�-ݪJ^�t(ÐP���|[H�c�,/���u�V�N+T�j�Fxs�vA�Hyb(�f:����5 (�E��̬)�4�6b�nj�'US�9��=��6�e.�t �<3��U)�M��
)��6Lϥ��Ԍ]*��uK��*d+0�?#P�`$�z-�KM����}���I(M�S�� �A��j�l-Q�0	���ڍ�W��alv��j�>�Hd�ZE=|$c3h��В��c�ڔMP�i��p�pC�2�	��J�� �D����M���s\��*Um3�&о!*�Pk0�U_�VS}����9H�FQSO�4���Ca"��F� 8Gv�?`�+E}	,Q�z7�F��p���`�^�waA��ݫ2��/�3�a�6,�I���7�e+g�;l���5gL}jI����2=��9EMLгb�ȁ`b���U�R���f���z�ffg��B�eT�Ѡ��I� "���uq��e�����S�EK�va7��d�YK̊U�+>}�;��r��)�jE���g~^m��&>/��'�A�<t�������L&��K�WD�^�|�o��O�V"4��!,������%K�0��c�h��7� :$�~G����������<���ܜX][��X��������<��z ��-�h0�Ȕ2@�<8Ǳ����k��F��9|��YXA) �\'Hlhz�CQT�cLΖ��4���ǎ/zы���\�ˤkes]���r�Y�����OZ<��Êh��-�,��rj��x\N��RPc�	����������[���^3�^�{� �+@d3������bfnF��ܯ�x��y�"��?�G񝧞�9BO���Rgl��ׯ6��W�/��[i3��h]���v%�����������Kb��>5���=��A��ϋ�{�Ңӝ�o�|�K�S�NE�<�?�Ӻ������1�'���:�P\%i�����O���]�~f�97;�&��e�X���^
�%�-Y�P��!���"ʻ�[��mo'O����:�(^Q��&��g���aϞ=�����յ���Dr��3t�<�2��¶0��l�|`O=�B��'#�5@\�*q�����aa��='z�ސ���������e���CM(��4��/���ĭ�����c�]��\�*'�*��W�:)�g��a���d$kpϝ�Av�y����:�I��jm��k���  <L�=�n}�*��^P+ R�J ��ʃj�⾌>$�..�>r���v�;Ɉ���m������c��MxƆ���1��O�`�� �6���a��.���~㚉nqqtS���_��3(F·,MeL�3a2���q|E�'�D�©�����@pJ�/_���E��ƺ�l�3�E����y ��n��x�o^ٳ0���hq���ݕ�4V�Ц0�N�Op��FFn��U���Bk�|�%�0��F���,� ���b�=���W6��&��N[KQ���P��;]��Y����֕���G>������
c��+WbIz��'P�I�(\
ʯl�XQc&0�-�������o����u\/W��J &����"�P"��C�H`��Ꜩԁ�a����,Bu�����}��h�2?�ʄ�Jand�Y�7fZ�K���>y�7���g�������O<t���;�|�ɇ�6a$с��8P�������&P��x�l��a��9����*n�� ��.�x.Mz�������}-+G�(�ʅR3���5P�7W���b6H��~����׾�1Pb�����#�F�~���`DvA�m�ml �]�<��S�?~�-7���G�L�Ay����ۤ����V
��3 ���F�+��sl2_��^���c�?�Gb����w�Z��v��Z=q$���������%�����/~ɋ�:���	_����Za$ѽ�=���� ������}���%� eD��\[]S�"�����~W5��;����|��n��[!8�ǎ=��X��Z�0�v&VP\�u\�pq�'�" 8x�S��=����ܬDC.�MN��i���#�۝�^��Rű����}��/}��t
�]��(���b�=J5gt@uX�7��IO� ���i��%���"h�(��%����V�76�L���<y�����d�x���R�;��8]��� h�+�1��ow��p���o��w�|�O��nG�q�w���,X�>y�߬����ן|�ܹs�ߣ��P*�M��@��p��r��v �� ��=U�G����A
�s �%X�_��{�V�^]Q��k�^0�C)�>�"\�t�R�J�q Z���,b��̊�U�D�P^�{Ao<77����k��E�I�����B0�j@��u�7۠�%&ԤB`&+�
�Aqx�:X����Tt�pKp��&Y�;�x2�b9��YA��Q�{~��bz��:H�lo�1��zAu+K/W��XȎ�@̧�J���ݻ
��f�� �5բ����/��x�����t�z�ω�%	`�C<�	0M�����$CG�b�K_u�c!$�{T�Հ��9�(���8��G�otu�jPu�CP�N�Rt�E/�+e�p�r�JP8Z��BP�P)<��QkjH}�[YYY?r�H�q��V���E������?2�m� (�%̿@5�����! �i����_�9˸ °�A�D^�DQ�m�G�X��s���'��\��W���`r�n�����)-������z�X8p�9���˹��ܰU�Hddm�&���3"`�0����$]����':0��>%�8�|!���@�N6��0�� ��t����TQ�GpԵ�s�䄐�7|��~����\&�bB��Y��O�&�?�=�'^/\�Pj��qA�R��$W�	�������N�O�r��0�9�0�vBڐ�OO+Y\$�HW����Ç�� p%&��Μ�7��'F`����#���x:�t0@���U�w���╾o�+I��t�4I��↪ FWH��u�ݾ�Er��jQM�7�0:��#hP��K@:'HP�C����)�A	�:���랔�
t��J�UNu>��'F��D����鈽���M,���O�Xɉ�Į/���*�k�q#���,'B��ЮG)*)�G�iNG�����s �^��,K>�c)�N�8ԃ�Y��c��	E�?�s�159�s��� +�8�9s�y�M7�I@p��n��>�6�E�IC�t�k����s�z5lx	���YÜ�KKK��I�0 Jl����J��RU�q /�ز���Dl��!�?�hN��n�����N'���c!8�� (�J�o���D�t�,G&�,m��"�x���,@�����D�����p:�K2��w�Z[�ݧc�F#�dg�HG�EW0��;d�;�����I�<ڃ���t�O�7�|��':$�6)r�p��DtewX��*7$��H�'x��';�]w]0<�~m<?���L��w����88LB���\�t)�N���/t:�a7n�E!X\\:��8r���!$g;�n)&��JW*��`�fӕ����/��� p���)�:������W#���!�$���l�������&��Qv������\�r%��+`EG�g�W���A=��g��W��  Q��+�"���`�9�K$
x�+V�s NT9r䯞z�!'�I�=ǟV�D���>����a)�ӑ��@NW�=�$�X� :]a��N�����Z[[�	��U�$���p^�4 ��y���8Μ9�v�mb0	N�ď�!8���U��ؓ���)W�|-R@�+�+���aQ�q�7-�T]�|"��U�*���N�:<�,�f�!"|��h"�g���	������FK����s��BAp��<5?��'N>|xF��vS7b���?�}�v�Ԑ�E�,F��N�$��ŋ��zBS.�A���O<��$2]{ւ��#�JE/��|� A����		E���x��Q���3���-���w��F�@p��lk%t�i]�s��ť�V6%�b�S�Np]�t=�`Ο�0<��t�B��`�O���9�b.�8 �BBäӽ���B)
/]]�z�Ҿ%
 ��j��7�}M��к.���^�TL &�=�*�fe�"`r��"i�#�Z��5l_	���XJ�B��"B��Ν{�����}����!p���@xO���x���C������>Z����a���ʼ��HW2
��z�Q������������o�P(\���n�����ѣG_	8���?��3���{�wK]@��O�~m���!X����|˟������\��X����y�-������/}�K������?�������Ba8`���)F#N�<��c}�;��A8��n��;�����߾r�=d������y�3}?;;������>������-7~0o����W���!?�
�ї,@��?v�X�yX�Cw�#�o��8�w���
������gy����|���8�����{�k^�#b�0Q�&�v�s俿�%.�$�d�[M�o�D�x/��+�� nw���)J�2��2�<=�C������a� �(�0m�g*(�Gp�)��l��0��;�}�K_z�[`��0�;�yu/�=��!�xV��9{��~�8~�[��/0��� "���2Lj$��Fၨ�#���x�sh��Y���a�I]4�a�~�/��/���~��>:.<����\�.�;BU�'�xҩ��8������{��: �|>��q�ŏF�4,�A4�v�R��ȫ��1Bt �P{!��ߠ�>��ǁ 8ȝ��k�x�=���:�w�0\�j0N|�}�hl�<.�8�<��u#�(j�_	ȅR�+7H�`ǉ�'���_�Cƨ{�DV�=��D��~��u�C�6�����_Dw>i��ʹy�&jkP�<K��|��gŘ p�������l���&�1S���y �'�Kjǉ��>�����݅q[\��oxY"���={vlet&g�(p�*nW9�ű	3	a6�4;V��ς�Dns���g������/jz._]��Z���8����QC@}-=J[B�+�ޓ�?� ���Ǐ�H ��R~�$mX����V�6��l��u���^[F����ĉ�B'���0������7;Nt ��pEvX�W`��<���|��w�c,xNX�[1�-'��&l�j���Ia��	����T+._�<��p��'��k;��_(����F��n�ZVm��D��)�}�IA�ٮ��KE\������6�|px,�{���,��:�;?��x��W���!z?Y�8�sG��+�@���&����h������"�J�Z������u4�{���':����'c�;6ҵ]�,�8���R��?Elf�ཋ~�_�3��I| ���s�;�,Wt֋@��L�A��%���zk��>�Ĺ!C��JS{�q��@�~�Dl��G�pN76.���R{��z�0D At���%o�{�%�b·
777O��8VNǛ�����5�		M��D��kaR-\�rylxb��L��29��yА�`ǉN�N���7���]����h�`�r&���!NR�Y]kU�V�w�aii�ظ�ù��cʏ�g�~O=����� :g�pe�Hx����"Cbmmm�^��t���;a~��r�r�8jo�G@�X����?��܏����N�0��ϡ�D�
΁OxR���N0�@�D�?h|�r���a�����Y���$Fտ��J�F�8/�V�V7�|�جl l'
�Gp|W��p�Eb!ئ�!��a�(&�9<(8���̻�#�%;n�m�w���XM)��.1�H��*Eq��"/^Zc�4u�1<�ϳ_|?'����ؾdqqlh���}V�����g�w�G,�S��p-��){�G���+�D�ddEW.�cD���^ �y�ѱqd��Q)pqP�w�o�_������ :V�V��<��׽�u;����
�v�0�;Ǹ�E]�W5<xp�^t����&5�G4-�Ř�?�*j7nRА��*\&�2'�s����|�wP���_ĶZ���`w��ߔ�٭�r��wqBX^^kk�Җ�J/ŭ8��.��Ǌ���u��U\_0p��~��������1��,b�X�%�q㬠��?{=�*KKKA��':99��_����A���K����]B�͍,1R��Ձ~)67�:�!�Kf����B��M��X��`�j��?^�6�q��@��X�E�"�b ��M�#��}����;J�X���SN^�!
��Pj�PD���Z��¾���?��?~B�n��T`,���	�ʟ=W�7�k9��{�'�8p�-����	gt)�L�!�+�O�����?���!�66�DJ?S�$�n0������>�J�&YسX����_?��~�k��k!<�z��(��7����5��~�����ǖ�G~D�4�8�q����H� (J�A��W���=��3֒9����݀y���'pZ
�1�du�������_�՜E�]�ۿ���� ��:�+B��<�������?��#�<�|代�YN�!�ߨ�Ф�{p9|�c_��W �{ϸq�s�,�/�1�Nc�%��~���:���+_������w�Xl�]{~^,��b��@���������~�3���"�8с��`��nuu�Mt��!�k>�8@���СC�[����/zыvdE����g�yS��z��в=i��P������0ן̇~�o�~�����3���!�뮻�7O�>=��>V(��R�3w�#<�裿��|�O��v�A����k�Z��_� ��BE�h>�Ey_������i� �U���`R�}I�(����x�N�|�+y��'������27܎nw���_;u�Tt���,Zg����oS�����^��׾�DhBt�A�'��:�y ��`���kH|�A8�C�sO�y�#?�������ȑ#�{��ǻ ���ؔ�����LO_|!\�|�s_��?�����Z��o|7��A������L@�}��M1!V�+�~x�����z'L�[A9�A|$.�%=�o���٧�j���n���K� �����"�T��/j�u�ܹ�w��]
W�'O������t;�6�Y��%�x���Ή'���g�b��sQ,`Y"��8�@�A{�¢X�Ɓ$�lΜ��x��᜵�� �V��
�2E��e�� �3���7�Ӊj�ħ�ފ�\�X�D��r�2[@hҮ=�8�3�&'��B�s�X��! 1{o�ߩ���VVV&�NW�D�,�Yt�� |em�
DW����đp䠍�r�m?���P�E,S؇�݁>z�ҥ��{�Hp��G! �%����P��^o���Rb�Zc��k��8�����ν��N��ޫWx��4X�6�柹�M�v�Y__/���Ap|C:���`� JP5�ä���D��H�dC�U`��6���!%) ΔI����A����_����xE:��\&Bt��6�	��Ժ�|vE�spN�]� GglxM)q�����]�����Aɱ>��:]�&̺��ŋF����'m��� ��bsCč��S�On�����hs^�UKp�����'�$`"D�ӹ/�~�G����.��b�ķi2o��Lf�F4�o��%�+�|:��`L��K�$�""�{Y��9;;Tl�Q\��M$6 ���bP+pq$ Oe�9�>���׿ޟ��7R��D��'��U��}���dx#â6\W�^���:�������o�}Rg2DW�Ex���
�BoS���'����,��Z����KQ(4�>� ��t�We�%8�~�!J���ѣGCo�f�~Zč�]�'p;�ҝâ��(
o�&Bt@PvB�"$ ���Ow��ŉ�
���
�=�)(GN�v���}W����lN��T�K1����	Vfh\�J@�0Պ's�F��S�Μ93�RH<	�x��E�(�<�c�&Bt���LH9�M�.���;q��m%?��p��ؠ�����%EbP�g�W )G�C�u?��Z�=��/&�]�)�'q�Z4F,D�e�Њr��� �a"D����`Zo����@�L&e�p�#'�����(�Lxv	��n���qlnnN̒���@Y���;����o߾�D�.��� ����+++c�3�$����`��B�O<\c>]I�16p3@D��ʜ��x��NW���}�U�G�5�����O;�Ŝ9�QRP�%Rp ���+&㕖��t<�G(::���u ��;^��͓8���COf�I"�:I�"���skP	��&
�ٵ~FYW�\	�W�Yw��u�vNAc���-i,�AIA]�שׂ���K�Ug-'��h�s�B�"|�'��>�"',Ln�*+�)��X��Q�:FN8`j��L����}%C���>=�+�Wr�W<݊G(8����LG�S6τ�WK0*�m��ä�Ι>84��b9������`���@���ɥ�&.�b����UV<!��|���Ͼ�d�8]�:�``��Q@�Au�,��?_�t	��π{P��oŉ@��_��L`qL���C7��e���A��)X��ZK��w��Ю�
�-ֳ.S��6':PW�+"!X\���G������U�a����r����G��v�r:�0���_	g_ �l���y�5|�X�XZZ
��ǹ�r
��H|\�\\\9�cĴO8-�<���'��t�p�h�֑�c�9O?�!�XE�/�	�	@�?���(�3U���0)NgW'r�7��zx�ܹ�:ul" w	o�S�hB�y�r:�(ܯ������w	��tV��r�;"!�+�Lx�A�^]O��>;\���N��iB�L�Ϥ�p ��@�k��I�L�H�b�KQD��_��ל�^�G����A���q��!��C���SW�#XG$�8rG�Tx~!l &-��x**�#����9����r�����<>�����L|��_dM �7��!�=�3�A�ĕ��t�`,֏��xNW�+L����v���*�+(��# �����p
����s"<s�����OG"n@�F����k��A��PD���o���K^�`8��{~18N"Z��/qCG��~�����?�p<�4�r���s�+j5mb&�"���o�����7$�z�Mh�������������'�%uL�Ҍ�d��Y�T�&!�Ud�������`ŉE�R�H_"X�����;�����"<���_�3��
��t� X.B}A�RD_9q�DP�+��J��4/!Pp��}= ��6qv�1��S�	����L�����D��Gz�UПy&�=�=7=@�q�6w����!���Eۨ��0u�8a��N�y^~{U���̠�YГ�/����� n�!u:��6��p�@���IE$���Ć��/9,��:]��r:$r5�@��6rd���
���s?�s/�{ޓ��u'��t����xܧ+�	&ʮNTni�H�}q�r�7ݦ)��5=�;���'q;v�������RDp~>,���&�eRg�-�`}Kr�9�O�n�q��p􉎷j���s��QW�^���O��]��P <s�^s�@��|<8�犅���a�^?�?��� �/���QK3��&	Ep`�=�?s˕� _}�'t���p�9�
�d��哹�����9O�������% g�5���GQ�&X�S�OgW����B�#!����i� �<z2������[�PdH`9�`Ra0�}\���r������5,
/�1�O:]pp�&Ա�tNߐ �e�8]��pz��9i��+��^����3�R���YB:�So����M�����
��o^����J����ڂ��\
4��/�W�{��z�����xE�ߑ�7$��秋�Z�V�zދ_�VfЬ�i��lq����<�9���y��w���O}*�9��|1��ؠL�sDT��%��9�ЩM~��G�U �*ܽj& �av��! �55���w�����@�K���������t��P�%!�l\_�[س�y�+_y�g>���ڙQ�"BQK39m���R��� > ����Ƙ;���J~�+|73)�C�41>�Ec
:�t%q������-��.C0��588�ӕ��%��3r���������;��;�	 Jć80q8?U,�vR&{�q:�.�W�^C����:q�6RH��s���M�����^E��0�.�&/��UH���8�RŐ�ד"�9� ��y����C�P�L0\�⟑�Qckރ� �H�6�&��%�0�s�}�BwW�uC*J��c�؂+�!4�����|:�Cp���t ��'�:��~gϞ����*֊�tN�0�����������=� ��=�p�DY�{�K��6��E�}��B��N�� �\ ���{-$�!��\��P ��JW����<�E	��!�k�!�ؠ%����R�+W�t��ַ������ J��m�q<�Va�Zu�z��#ItQ&nL��� ��!���E.袕3g�LL_�8�����Nn��I�8�}$h�8���<��3AS�`�
k$Hg"+��W,
��l\A���ĉꩧ^������V��ɓ'���	�*��3i`|��6���"g��p� ��Y��~��'��E��Ԕ�f���A�&�2�{������H�Z��~%_0��� 5 �or��a�~=����}���|�"$L*��Z��:Mߙy��ׇ޵/7s��
����KG�������!�.z��D��{�`R��S<�(�� t���+,�O���������*��Y�D� ����/1����wI��I�2qf��s�S�E��k���+�c� �~��뮻���7�����?��!e��ߓ��1]�a�=�T?��Ҿ}�����g�gr�^zE����f#$�!�N� ����|	|N���8]a0�#(:��IP��n����t�666�柹���.��%�b���O��+����;D��`��"rd�&5�����t���r[oR�(��&6� ���}��ŋ��Si���^=0�!N������ח�k��#�0��&�1I����|�W�^Z9b����9��� �)��mo{�����`��26�C�҂�8	7��N�s��F�[ZE��	B�t����?�"�\5���s�i�$8���k­�ɍ �(h�IU��U�M|���z�>�w��{�� G��IAE��� b��I��v?�����o�0��Q�����~/j��!�_	t��|���4�D��������[����4�E�G����`�.�қ8�>}:����]�1�
x'΂������Ͼ�w�w?!���E�U\�E:'��^a�}��g�m2|�С�m@�{��8O�.�?�ِ��1k��)�CE9>�]�p�w�-��I�d��i� ���M_�\��ƃ=H���رc�9s�f�����r��fo��_�{��{��ƊJ�K�F�4���Γ(���غ���%�:ȼ�b���?�y�h�p����g '*��W�|!8p`�R���+{�+�R?lS�׃��>�%�%��Z��9 ��/��/����~��E8p�2�c���"��,�|t���! D��/�wˇ���ꗿ��\��V(6�!��#޼K�W��֭��*&ot��-U�~U�
��t���]ɵ� ��A%��/}i��zk�������ѣG�K���+/�#'�om�ٳ'�_	���s$)���$l���N�裏����<�[�X���ŋ��� r���z� �s�� �"��4,
9q B��{��DH ���t����^ח7�t�t�t���x알	L���O���z{��?�p�H�Z��7����{4X�")��ө?������t~�&Z��M�0���]�%!7*�,+:~�xЌ���ć��sd�yS�yI�~?��z;M� ���ͣ�=������A��ۢp"4L���i�ԹL�gF���0���������?s�0��80v����"���4�q~:�t�2��8���3����u����Ξ=�f��(�f94����fPU�'qb
oU�P{N7]��:������G�Nb�yg�
R�s��l6����
�E@���'�_K�d��`�}�J��c�=&1H�I��&����w�A9�ߍ�! ��ɦkkkSW��p:�8Tvi"qbq����M�ڲ
���;(e�a�]�z�'C"��]�yy$�+�&�WY��t%q
OlQ.�2ġ^�O��ى�S�IQ��}j�e/{٫>��υ�[}�g�P8�Z�a&����y` MWa�����0�b�	5|�����&���$0�!^vp0�u*'�������LW���c��PmoF 
zp\S��:q5޹ɜ�95����������Px½��ɚ~,�h�5 ©+�qdU�� k�Á�z�&;i�(˄���>����^�
�yjSQJ���U�(<��B�Q�i+3��L)BD��k��_}�mB��1�F���m+E�o߾�����-.
��`?���R�0X�Q���	����7&���E��>d��� ��^}��W���`"�;�����"�(\��H?v<ty_.��HQ�빹���2�~%�L�8�o�h4Bw�D(�X�#a��s�t��G�T�\"���Z���9]:��e�BA��&8���L^�G�B�9�@��ɓ��%�8��y|L����tE$ �$m���ו`�/A�銀z%m��E��u�]g�]4J�F��Q��DSĕ���m�B¤�`UX�N����OB�sVߢ�h�7ԟN�8���t:����:�xӥ����8���IE	P|����Q�Xx~�&BA��8u�TP�����K��1,���¤*��ϊ ���s`%��}!8ܕWZ�����Z�
�t"$ ^�¸.7���1�.CBx���q��\��>WB��:��\�\~�t��#�<Zt9b�;�U����t�A���\��O"��(�<��[�`XT�FP�_*�ۄ�n
ǃ�	&U#�8O��*���zH���A���t܇XԵi���P������&��7��z���?Lf��B�iC>ǫT+�(A�/-5�D�g~aa!��x�J^G�w���L����T_WZ^^�9��v(��3�}O?(�Z�^���c��f״P|n��.N�Q�W�q8r�Hp\}=���%��� ����M&yq�q<]I�H��@Y&>\�|9�_	p�e8s\��{m�Z+��i�I?q�;���ʞ���~�Y?oWZ����N��ӕ|��pl����aCvҝG�n<s؇��q���Q������DZo8��]�޴`2���?$��NG�9���q��E�9�	��L|��&�2s�SL瀑 ��:��Gxx��]QǄ�Km^�:��B�S�x7�I�I���h2�}���ٹ��[�E@H��ƥy�&��������+��ߗ�Zr������=1�~yyYqb]��r�íN�:�9�g<1�Ju'�>!Յ��駟�~��|��<+6/�@:Wxqe�Tp�|�I�v��[HQ0�|n;v,�#�i�Nָ (UݯZ[ZZ��bk�����<���2��L����Gb�_�Z��|��������0~���":d� �aR�~��kΐ�m������t�#�t��ᢂp����o�9(��};�g�1��q߿�=��ˡaR���})��D�?��H�<5�[�� �Á"]A��y�+����w�T�+��S�i�A
2]'џ��I�[_�����:Q���`�g����9�y�t��&3�3�*��I$�!1�����Q"2�.�ߛp�O=�TPN�}��gʣ#\��H �5��s��$e��W$:�V�D7�]EA�Fč���6Y�a�����k^ПȻ&�۷o�:q�9�s��k?�t����@P��Le��U�c%З��	8X��:&o��;���t&��@֏��<+�~{��$c��Do>�A����AU��@��ǭ d7��׉(���<yrKzO�
+��w�}߱�߽���!����W�s����x<+�6��t�.��Bp�%�]�D��a��v!8��.�]�ۅ�Kt�v�n��.��Bp�%�]�D��a��v!8��.�]�ۅ�Kt�v�n��.��Bp�%�]�D��a��v!8��.�]�ۅ�Kt�v�n��.��Bp��cr�6�|    IEND�B`�PK
     Ps�[Ɛ�~<  <  /   images/e65d6d59-bd1f-4659-a32c-fe6c1b0070ef.png�PNG

   IHDR   d   �   9ty   gAMA  ���a   	pHYs  �  ��o�d  ;�IDATx��}�%eu��W�s_�m�Iw��A�h�DQ$����(1q2�,��k\fMLt�8c�%Y�NV�BL�ɬ���D�@F$0*J$#����@74�o��9U���{W�S��sOrf��p��S�����~�W�	oy�[��Ԕy�gL�&I�y�����yӹ�>��陙�V��6� M�hll��w�n�^�M:K�l��1�Ld���R�,u;�Yc'�ƢN�㌍�5S����G�v+i��)~��vb��P_/������	C�G���&��hzʹq��ܱ9K�jE62ݤ�辈^'R��բ[���Z��OiL���xk���!���R���q�Y��&&��q���╯�{��Agbbt�I�޺u+�en��U��@��G?jN;�4��/�fh������/��/�����'�V���^���U�<���W=:�>M�݇E�"YB�G�s.B��ƿ$���.�]�8ZI,(-��"Z3ס����h �$BX�-&�o_\\��<�q�o(�]����A ĤI�&"�0��!d��Cm�����Iw��vi��̷[��b\B���ݿwowjr��Vk���v~��_���^�v��{6mJ>�,���0��Ч_�ݻv����{D���>�z���O�������-s���cǎ�E����7����W��u�~m���G��J;w�&I�e����6]�ۢ��2��{�������xl��y���"dƦ�{��GT�ۏ�zJc�B������a�8�Z�f��D�?�ir������8j��O���Ng�(f�;v�|��̈́��3�3���ٳ�>?��7������p��]r��~�ۮ�A��G�e�_`~�?ty�\w�u�+_����6sss�駟6��s�y�;�y�s�=��r��]�.��׾v��%tϺ4u�$!�# ��F�ς�D�,��,/�_$޵)/����-D����'� �b>��ฑ���o�ǀ$��o���w�Aӊb��n���B-!褣G��E�<��Ni~b�޽Gv<�c�կ���N�}tz͚}t�Cc�����;�

��k�m��f�O�;�ü�5�y�ƍϿ��.�]~&Mp=�@�l���'he�ؕ�0~Ie��{�K�/�(�9P�a�<�/�Q�t�eMD�?�潆>B������s���蟰�R���Gp��f�'�ј�,,,���;�ҙ(�2I��8p��N�kɹ���o�f�j��|��_��ċ߿}��7.��)�N�����we�\�3����"2���Y���!iߚi�p��MN�tgz��g�J�1Y����寁 �;w�S� �<�N�͘Yoh4������ݩ������w�;�y�r��@k������z�9�s��U�=Da�b�+^�e��He�]�2ȜK�,�k��О�vA1���q�l����gl+6����O?k�|�ʮ�� $,�;�k���!o�(�5~�M�}J�gSMU����-�A��m�0�h@�^.�Կ�@�-ߎb�hb�6n�zvX�\�����\�=����{�ڼP�NR?����Jrْ_{!�zPp��3�0�抠})65x���G�9:��[ݣ�+�- ��0�
[�G4#�y�Q�=�	�����*��VL��g^\A~?'�r��&\c%
��mt�{�.M���?m���W�[@Y����>'\:��'5[�&�]LM�&^�۸ȋsHMƮ,K�VfY�%����3�No0�����jwoK�L��%.�і����]l��Wi�*>WT�W�OL�kWaJlC�A�[���Z�ds�UV�E�-˫��e�/T�R��"�o,�f�k�hv���:���
0Ɩ1�P�ڄX��@(
�ͭ�*���B��U��@:SE��A,&m��+�V�6+v��"̴�, 㹵�v����pYS�	�|βrVeL�@��I����ԥ�[�����^j�����?��ˎ�����+�5�m�� Z�t@�Q�G�"2H`%��+��}�)�&0�*Uw9{��v�u�k@L��jMl+!d,%]�3ݣsQwq���J��;+*o�p0�@�L^�2o- ��{9(�lj�=��UV��5��V��}i�(-�n�!G�D�6cG��AZ=�B�a������W����gU6PL�걘���f��a��Yʋ�)͚:�'�R�/4��-�k��a��R=�BD��=�1�J���@��d�W�ګm�aΙ"B^;��J��]ڟ5�E,����!Pu�E� �*qNMZ+�j?�0���m�n�:Ѱ�ؙ^����c,0��[�+iYZ%��ڨ�� Q7~u�O�u�ϽW���l�n�
	l�S��s'ܪ7��/ڰl��үY�$M���b[�Zd����~�W
u�|$�����Vk?������z�blFMi݈hd�J��姙��f��ꛐ��ԗ�|�ߣ߷	�c��Y@|Q���I'FbDx�U�Fc�a���A�:D���F�n=u�c�U|7��<e�iŭ,ě�����1m�|UP@!"\l�"�k��u9vF>aQI[������	���L���ѹBm+t�ڗ=��U
u+��&�- ����q7*A!��������Iа�<���E�M�*s8��e�w�+��<�a�M�����|�B�%n�ɱ�_]�p��W�lnh#�(N�hi�2D�)l���A@�.
�2%�1`y-311��ۅ�hc�h��k
kS�h���|l�	8d��lC��+m��a����oD!�0�$Z�k1�Sz�;%�<�0����%� �����$6�영wX�Lycd/QA.�ܞ�����ZmgT+Ңa�^�5�M��k`�XXXhD!"CH-�r�P���a 2|�eAT�����&^��J��l�!��}��.��gKT0���ex_���ʣ��[����QÁ(D���v��^�����O�<!."�������<��:�c5הG7��PMl��A�r7jZf�{�rX"d�PI��!�N��XS�������1LX�Ԯ��rw;T�ISh����j����Q闦
�������R;����6~�����!��4��nK_h׻�M��4�a���>�@U��?����$l�+iY=w�����&Ě%OQ�YW����>�����D�
(#%������n �.Bjk꓊i�s�z�$3�;<�/��:���_�LQ:��Mr�g2�"�Z��rz����b�Fky�,v�`��}�T�f��:19�{��$����a�'hYq�%6��芈ql��L��>�L���V�:j�������1s���]��B�>d�:t�{~s����8V���1�S�=9��99�C������8�˧o�'�ĺ�)����[cx�}���R�BN9���a�77w�dB�W�#Q������`<�<&��"yfoQ�;ś�fT�ϔR�S��1~��'��q~�FYz*�!8F�&�1��)���Bz
�"X�M�J�{ģ��Ě �s��D��_@�X�l���2dF�6K���U��M?�3?������ʿ-����jE��	�X@�T%�y�D�ƭ�J,K�l@���|`������@LpR�B1�~U^V�;���8ޑv�"��4�y�����B��_д)��zuA=�b�)�(M`E����E��9`C��OD׌$s:9Ū�k�`�u+��T�@����NA���P%�\Z0|�X��9?ž����}�#D-��ߕ���G�+h���#����\����t>$ؙ���G�e�W�2��=��yH
�32���ld$��byTIU}Db昤�Z��$MW��n�����bk��Q��B�D��A^o~V$�}v�����+�?U%Q<�׻̺�w�����XL�)ҥ_I��/�}@��^���h��������>��"����!�!�G~�A�5��[�c��'�F�: .w�s \G�dFbh���v��;E���
$4��%i�(Dvwf	��[����ِj�۩��� ��h 6H\p#��*�i��I�s3��dG���L47���B� ,-.F��*ͩD��r7Y���[6t�d��i�T�eF )`�	+3~�fz>���"8(
Ð��ցÇc��4�0��.:�lI%�~�i`��}4�*R���_��e�]~j����
H�aA���i8>��o���wH"��oZ��.�
��c�#��,�4n�H�>�-��� ��
>��N{�ˊ
���Ei��_V�Ϭ�!��!��Y1^7�G�J����Ĉ�4�BN>�d���N:��Փ_�O����X��`]Yv[����Y��
`+>��9���S��W}t<��P�5F�r{�u��d��T8���6������g 6�;T#E���NX���FT�W܈��F�\�\Da�ß���*����q��V��x�w�U.|�QN_A'4����|�~�T�H�"���2�2K�U�!���l��u�ȇ!���'p��!$�g�kO��.um�Y��%�P�K���J��p[\ZG�#��-к,dU��i곴���Z����2��pu���,M�rj����	����:|X��J���a��	�n[���m�~J���H�]��(n�G��VUghpp���y�r�B�[#�-�Y�?��:�	*>}k�Թ��;�%|�w�u���f�I�̰)
��q&*��?���*''�rCP_K�<�ٙ����u�Ԯ�e<x�Sȑ#G��3�F�W����E̬$��5X��D�8�,��Sri�5�g�X����*'`�#�!�����XV���u!�J��N�+~R)ԅ2�Jz��U�%>��X'#�?�P}��	+X�3�ڧev��5���ij�7Q?HU�0?���Sް&�H Ň�SG�q��8�[@��G�ʓJ{��LI *�F����+%�.eK�ɍJ7
��͜� ��eE|�J_d<M6�3�dN���Z����a�w���B�Į�t%��aOO�\�'�,�8iN��<֫�^3�\��5��"哇�,Dh"DhlɔY�:d,YD�p�����C�Ŝ��V��1K���,
!���w�*'+�BԶH&2wt�S��[�J���gFV��=�Q��{+,K������b��;I������W�vJ�S�0��E+�DB$�W�x��������rHu3+ջ��Ÿ$K���ȩU+h�jh��2H�OIYӇo���G�ۆ��V��qj�X���+�33�s�}�!�e�$h��פ+iY�$֤��WlK�򆤸���W�G�R7�����p?'��r/ϲw+�'zoj�hR��!g�,2?�m
�"®]֢��T-h?WJ����N!���- j.�T���㳬E��;�����IF� $?+q^R�.�
5&�E2?� 2�.�Wz�y�ȇ\?q<�a6�g���o<��N��?�S��ύ���~C��Φ��3F�v�~�zo�\z�)�E�!�����v/v�ݓ���6	׹zW��"[e;�t��%�M�"տ2D��3݀m��/��[��|y%��#]V��l~��fR(>��+�:/CKF'�wr��i%�����5�f�X1W���@�I�g��P�LY%�>��$fqq>t@���[Ǚ(.�X�_�x�0$����c~dL�����ٖ��,��ޕ�1{����3'qѻ�Xpg�/����˂BB�Z�#圧�_36o�H�u��WΟI[����"B����_���/�+��y	��
A�-y"��A�瓦�<� T��ש?�����W��~S�h��LcR��s�0#�&b.1�ieK��Σ	.%cUE԰	�4#�pX�J��81��B���B��c�x�I�Mćes$��j�F�k����Y!J��'W嫗xv�X���.۴S��Ƒ��E<�ԇ*�i9ȧ�?E���ʻZ	ٙ�g2U8����}f!3_*[�t�SK7��$Iy�"�֌2n^t�XU�6���m�?�Ņ��t&>~c��'_q����n��uY(*=���֤&�;���D�G��&D�=B� �Β߽�7k!�޳)G��4�z�	�I�&Ԛ�슍O�L��?���_1�Hi���;��"�HW@B&�x(a�k�F
���΢�t�Y\��EP��[%�2ݱQ�@�y��<�q��!�����M˳��E��<5���Oݎ����쉴�K�c��Q� {eɓ���pl��r�qʩ�����(�j�2�#�h��� �ܴq��q�������|�)^��=�˙��е��SS����O7�6m6�7o6�֭�Sjtzz��<���_�"��	^�ڄ.��b��;#��ʌA����"�_� @v��f�4³A���m[����5^x!z��?�;��gbr��u��1���_��ݚ �L'J�,��� �,�y�{�E�\LH�;s�Ƶi�F/���-䭷��>�G�H8HDQ�<��F����ȪK%M�}���u"��3Gf�Y�6m���6�qRW1�#G�.�yǝ�k֜d�" �B*s�-���6	5��ӫ[(6=9ٝw��������~�lܸ��0��>|8B�)6d�å�Qӄ�(��y�{�����n�=Fj�Q�B��׬?�LՍ���s���G�z�m�O%D6�� ��v�/'�8N������I�q�;9>љO�;B@�7]���[��{�؜gKxȌ/t�^�q�y�U�Y����/�������8<��qD6/�h
^u�����x��[1q���x��������f�1H��:�'��b���y��_׭��3O�^NSX�6jŇ���4����	u��-3mZ�=03fK���z�frl�F�4��k��E~�D���D���n�M�M����~��}��ѣ~��d��!���a���z��+�|�'���w|u�X@�gIն۾�Pgaa)I:����5�u��8�̳ӹ�s�o��o~�G�������O>�Y�����_��;>&�
�i��:I��iÆ��W��woڼ���u˟q@Mυ��q8��ye�y�z��!�n��?i>�ٛ��=�m�;>���,,�W�k��f��z훮������o}�\a.%�2g�&C�up�iR߹U������ҁ�n���M�L|Y�]�YR'�y�+��+f���뉔qϑC�C�y�z�`��؜����[�n��m��!�9�Q�"�}�xָk�n��;������o�4x����Z�}�kM����/��$����9r��9g�xT|P���&hkAnE^�hO�3֞ᵲ��~�9��s������d7�Z1��X��?>?����f����7_����裏�R�mo�ȳT$�����ɾxΘ�|��ꋐ?��?���?3��{��^C;�77���s^�H���Z�{~���e�_n>���ج�E�6�#��]c1 ���hҠ�V;�\XZ��ۿ~���g߁U��}�v����v�O�ƢZe�ܾ���� �_��_6u�L]��y��|�3���ױؙ�<����N��,�NLN�a`�fm0TgH�^����X v�r,7�L��'���j�����~^�kp8�)n��K��Ƶ�2�ڭ``dt���.������4(R�`�����ͳ�w���?B�E��@C�x�/�ѥ1%�C"��3��E�Y6O�k�>���B*
�{f�iA+�y��lѓ�Tǖm��D� ?� �SI:�.�Z��>�d+�Wqg�q�IH�qb���.b�|�=��� ��įF�b"�m�84�Z&6�B�	ffYR��y�k_����:ݡ-<�3�`ȟ�%���ҚF����t}�"'h������fY ��h0c%B��P h;P�%s�E�h�����g��P���"�e��NR*��!��؏_$��ty!cYa�02Iv�N�=u��hv u_�A��!�����0Ќj@J���A��� k}@=Y)3c9`�ѥ6,��sd�$B���J�s��E���&��{R�-�a���F���p�B�F�/l��K�h> 6\A!�X�z�$m	r�������D\�%%�2�=:���j#d�ڵ̑C���?C��ZyJ���7oN8�G"���z_��yU�����*6�}�9���}��b����Y��߳}�9b�v��u�o+Zm����B�cTRF�/ ��K������|=Ů,>�*L �!#H�%C��9M�q�?���s��g�u~EAM�"d����G�5M@m�������֬�|굊aa��B ����cMU�N��vpo�v��g.�+trOЈ���v��Ѓ�;h�=��,�N�Q��C�����m+���W��r�JM���);������^�B�.��C8/	�]N���w���*QcP`��J��8�g�PV�1��j#��#�����		�n]���9��ygT��?R��|����3�����'Ôd � ɦM�|�T�˂�o*Jej��A�u�ֶm�|@�ښ��w�6��K��GM�n�:t_²$�#��U~3@S�C�I�t��!ȓ�ǎ�u�^ �bZ�E A���h'���,7�F��h�P�� a���	��P �l�̎���aH;��������/�|��xGv�}�z�"�7ܐ|�C6�������y�?/P(���V{�}����n�m��f���:Sj#�c0E���UZ4���G�:��ڱc�9��sW��?��?�=�����RT��G��e��r˥��z��׽�u�2ڞz�)�k�.󒗼	/KGh~�u�\��Hy�n߾}w��]���=��Sk�j!�;�&��K@��rn����i:!�n˫^��w�|���>x�+.5_�җ̵�^;P_<���F��b"����vI�����/�����7=��E��:'h�@-�6b{o"�F�}jǜ1/ ��j˖-��C��7����y��W׋��C��n֓F�6"��0������B���i�_{�e��f�M��k������i��N�����>D�c�p-����~5Q�EW\q\(7�y��G~�GV��o��H�� Q��P{�ċ-��(���;��?r����O��ij@m�E;�4�ߦ�mց���n�����7��ڳ����{�UW]����Gc�i7���WiA.�w���ޣ �^��d��W�w�y7�u�]+΅��o��۷���{�_/� � ��E�q
m�ɺZ����	ki���m�$����+�kH��OT��J��1�]���Bȸ"��z�|�g�'���o\O�^�/���ώ��]Mm�Dr�5[�1q�%�����A-�������4��J�O�'���� �?���&j����٨x�O�L�OG�Ք���O<�#ĵ�jr��{�����Y���D��y�֯[?��ZΈ��p�4d�Q�rAH��h�����v�Z�YO��D���ӄk :#�	BRx���߿��e������ZmJ�� zs����3/"�2�� D��5R�F�	�%��wv9@��fhq����L�8�u"O)�'�w9��X�����;Us����^p��E�-o*���V�#��m��Ha2�d�������
{H��7����;�G���ƣ�Ϻp�1$6KvQYΥոۓ�m�]��s�k�rʖ��z��<N��9��TV�7��=����BxwdBA�+Ѱ��	y����c�	U�H�A3,�]ع8D�{5&�0����M򧕶H޵I+�LK�n/��|K����hZO<֔P�}� I8��S���G��;���B�Z8�J���?{B��"'���c���c#�1��5:P�e�><��EE��2H�T�H ���TDƃ"D���5��E��#1�1֪������D^�߅�Y鷜L!�œ�6�ic���~�y�[�j����a$��-g���0y�\���ڐ��S;c_/Wb�����8�Kd#���On�B.�|�y��Z�ñ�Hb,�GV����}�С3�:�ʒ�Bm��?���ה��H6$�{v%no�� ��S��'��_}xu,􅒬�kNZs�9g��j�x�d(���h���2�|Œg�,|W���a>��P/|�e�!��,M��J�Y�G4ˇ$�4�<��y����9&����c߻��~����4������	G�J���N�#�D�ޭ̞⡠.˲2�b�_�ѻLP��y�̬[���*�t<��B;j��	Ǐ-�N8�=>>��q���������(��UY�g?0-�)������u�ܹs��+��?��O���e��}(��� �N&C���t�w�
a������<{��
�:IQᘁ��(hff��~��~����WdYh������}�B'I�F�j<��������{�5y���n����]�nBX��p��W��X{��{��]"��A)��ϐṛ�Qm�����&#2 ����}�{�?������=�Ȋ}]r�w$������ٚ%	�3�1�|ٽ{�}7�|�o~�c�����}��aah�`1���2	�ߥ�_����'Z ��N�o�zʖS~���O_���裏�ڛ�1�n�H�ڙ��s`�E
����!��3O�{�-�|ta�3?��B�Ⱦ}�@��P��.}��9�L�:��~�w������2.������004B0�={� B�;��-�G�"��+	����c��Ϯ{b��E_������<��K��f��St�d9"'}��z����=���h���_�����{l���G}|s�y�����y��
���~�9����!�e˖Z� ��8�(�}���F�Ee�ȪDk�%N� ��/X�@i��9������L����W\q���p�Ї̧>����A̟��������0_Ѱԫ=�3̍7�h^�򗛺04B� O?�tQ�� 'V<]��X�CH�)>ع��LP{%���[���=�A��y��Oኝ%��C*)�pH�.��bw���sT��@ĊGaM_#���ج*��y9ؖ,�h@�!�V莩�'���ֲ�{�@#��L�H�+.T��zwh�p�G�椔y��$�U9<W;'dڛ��m��"܀��)O�M@Sg0�d��7�9�؈���8�(۵z��c8@D���Er�|֮ m0��k$)�'�:*��D�@�sD�s���F���0�}ᱦ�N�;+"��A#��~
y*�*�B��A�T5E0��>:Պ��l;*�*C~�^�T��Y��8[��a�����g���4_\l�z[�eAck%-�ك�2��f ��:)9,C��,�	�!�+��_�:��B� �H�;��Tg�a׭[W�p �ICA�l^R���l�Ӈwt\�.4β4H�8 �o��@�]"�AA�E���ڵˮ�P��t8WS(Q���B#�j� -d��1!$J��|$vmT�L]F�C��m۶�:�"��P}�L��\���:E
44Ʋt>���(
�`l�h
�Q��}u9����:QE��5��%	eF\��4Ͱ�`:e��$���h8�^K�*6 �����_u��u�3i-K�$rQ
X✊d86͜l�U���������e����q����k�F���}Q�9��ؚ�F�R�8��9���hDC�T�kRNrw�uhʣŲp46�@�}y|G�?�w���TE9�bJ�dW1؊*��2��e.��ւ ���+�O�_�x}ѯ�St=C�	h�p@_�Ž0	��J\�V���cۢ]�@C_�V-����&~$��.�\%�8�t���~���a�)$�9��*� r����3B�*]0By��iyҟ�l�&�1
�?Q=:o�T�\'\�*D����Q>�k%�Uwj��	r���@�ŸFK�5Y!L'G���r���:�^� ���Q�E쫖��c/�# D�A!#ǲ�r���T<�:ÃE��a�����h�N\'L-vrj�ԡF?f.�Yf�hW�[�X�~G���wPf����g]��lظ�V�X1eqt�m��j����b}M���5���f\'i����,>�N�Q�W��,�N|�Wϲ��=x�`l7�p�GqV�]S�
m.+5N��h�g��F"Ņ:�*����Q�zb�9Ίf�.V�����;�<�v��a�
e�s�vb�"!0r�����wV� �l�$<8Yx�X����*�P�^�l�Ey�9��lAu��x��P��J����E-A�1	9v+�l���X� ����\V�C�p�-����_И���A�U�VEә���u�¬,��K�<$�p��J�5]hEE�{k* U��X�Q[�W,��j�3�{Fee���@Fr"RC�A#͚D^�,F ���ǌ�P�Iq�X�Y�Z.Qqg������J>�L_0��h�O�1 �a���$�x ������յ�M(���d�P��H^�W<_�B�E6w!�� �Q$�����¶$�@�n�(���R	�%�#�C!��d���P`9�^�D��$9$�����)jb)`Uۿd�*k�"+�O<{�+_����۷���NJ?��+l4���BM@�jo!�Y���������Z��
�Q�Ca�2�4QH�`�j�S��HºM@#��f&l�WV���C�Â�YL]'u��C����$��r}(�ܒ�:r�M!���Oh���Ak?�H�(W+#]��d1
��xM�ãl''&�����X�L��%�&Z��c1$*�4���;Eb!:��Y���(-*K��1� $��[��ƭ�,+3F!/�R�v�@�����!����d�_�r��.P
J:ɱ�a����ζDC��be��	|td*[+�2
E�6�d:��@ �+|�1�1�a��4��$��
HA3����;#�('�z�L�!�n�b�E�-�rbb�u-�D��Ј�l���s��ִh,R�!�w�&1��^ˀǢ�ǆg��i*�6�Ȏ;6�ݰ ͑�\&�E��u�S7!
i���4�:��b��z�B�8Bo��ٱ���?uB	е��ݑ�����ϓ0?CB�B��ȹ�Yf��ڶ>��)���GNPqe��kP�!�����TQp��sU�:Иګ�D�����"�4�P?����w�7���wNG��k��_�e��t�둰�&�ɼ�B��v�����P��.:.��~��݉��]�v��C,E��>���6r���`��,?�sr���z�c9\+H����7���0LOO'��H�=MTl���:d��#n��Գ�"l196Gy�@İ�	"�T�?�a�G�-\���P<<&7rY'�����U� x�r�E�����S��d��"�����R�=���"נ�׉�kh��ve9����ϫ���F��h%� �ZGЪqfrQر>�b��{�T6�'�Z
^X���������jwZ�6@4:I9�{>D�Y>],2D�E���:F���j���kZ����t�+[W�����N?�������C�TB�mk���`��(��O�&��IB��z�>�e-�T�z{��E;4C���N4DL�)O-N��9�y@���H�g*kB��".�T!p��޽mg�Ag�K��|���u4�����٘��I�Ȩt�4�ۛI\4@-g����xV==�u��if3���d��\M����H(�)E����Ն�B��M;�N��� `d�=z����E����;�ա����iO�1T�:e<44)��QGx��} �Lq�RĚ�F�d��H�I�Ixf��"M@�'� ��K
	Pa��p�9���y� �*X�ZP�V�hY�����5Rv����M��`��D�jaY����֭�G����
%�4'7rǢy��V����-RT7�U�p�"���Y	�S)L��U��哭G�.C�����Cu)��(�U�!��Q���SO=X��Bf*�KVv�X�F*H�Z�,��YOM�	?n
���Bi Ȫ;vt�D�:m�[Q����=�H���6M��r²td���M��]���,,�:j�r�ds�z\�(X��9��;��@����ES�+���0J���Nv��yJ�G��C�f b(i�M@��� \ĥ��ۺh��( Y$x{��&*�`*�I�^DN�TL�8��'��klں�]v� �
�u�od�4d����i��h�T{���*$+Eg���/�j��ȣ�D��R�*1d٫�ÒȨ
M���U��y/-��uu�/T�সe`+��+X�M�6ن�;�b�"�$�"B]��64��N;t�L1���k��e7��^�ʁ0[7���K�ֲp$�NxQ�IHyڍ7�&X���U]n?��>P"��sQ�!�G(��ݮ(}�d����k��-�1|>id�kY�A�ʼ(��~W'F!�y�)P�J�<R���Oʴ,yR�|������e�!@H�a"�ƨ�)'Qh�E���v)�7RB]�l��Le�

��ք��x�N���Nl��ګ
$B��"髬�ۑs.jo/@�d�.�$}IF�,�$��'1 ���a#�TV\<�7�2G�BJ>�,^��W|��U��B�c�{+s$��Z�B�����O�*� �l?xp)n��6H�r1 tN�X��l����AV*��n=̫;��ȑeUs���C��AR#^^>��aYB�N����ԡO'j~�X���5B��!(�_;bȆa*�3@W� �p$�ԮJ���N� g�����Յ&-��>�)���
��(�!�i:z'��!�.���z�h���x�+����:�f�ԕ�(z�f.
h�!���1���sN\'�+���4���<�,Ͻ��������F*�p`ϧmH�eqnݞ��PEk�=�R�d��;:�6�,��,��mD������/s�+�&PvB;��PV+ǫ�j+'�Xv�F2�N[�y�����$���"<F�=[�B�:�K�O�҂81��ix�^�6��EO�\2�FeҌQ�$��4��>NWb��\ �/�����=,p;���OcW�����_�<�=��]G嶠<|�^?��eC��g36j���"I)#��k"b(ڔD#����j7�i��VK��A6�������� � ���+�@�L��@��c���ѫ'`�p!#'2bp!#'2bp!#'2bp!#'2bp!#'2bp!#'2bp!#�}�zW%`    IEND�B`�PK 
     Ps�[N�Y�R�  R�                   cirkitFile.jsonPK 
     Ps�[                        �  jsons/PK 
     Ps�[�赚#  �#               ��  jsons/user_defined.jsonPK 
     Ps�[                        r�  images/PK 
     Ps�[P��/ǽ  ǽ  /             ��  images/0b351edc-7875-4477-b820-546ce15be531.pngPK 
     Ps�[$7h�!  �!  /             �u images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.pngPK 
     Ps�[
�8b  8b  /             � images/a7e3301e-fb46-458d-916f-a05c0bde95f4.pngPK 
     Ps�['�Y��  �  /             n� images/4bf63cb1-3675-4452-8ab6-1403298522d5.pngPK 
     Ps�[9&��ސ ސ /             �� images/b01488b3-8551-4b4c-b09f-2812c4acc168.pngPK 
     Ps�[d��   �   /             �� images/d3b73945-fe79-451b-b309-b64aab767520.pngPK 
     Ps�[Vm�80 80 /             �� images/9ce856c6-be81-4769-87b3-53be9928d02a.pngPK 
     Ps�[��C�I  I  /             	� images/627fe4d2-0152-4b97-938d-4b9176d7a483.pngPK 
     Ps�[�c��f  �f  /             �� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     Ps�[��EM  M  /             �a images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK 
     Ps�[y�E�wf  wf  /             gu images/6a97e33c-aa93-4e7b-a2bd-349ce97096b8.pngPK 
     Ps�[Ɛ�~<  <  /             +� images/e65d6d59-bd1f-4659-a32c-fe6c1b0070ef.pngPK      G  �   