PK
     �a�[�łk_k  _k     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_0":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0":["pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_5","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_1"],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_1":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_1":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_2":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_2":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_3":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_3":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_4":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_4":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_5":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_5":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_6":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_6":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_7":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_7":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_8":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_8":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_9":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_9":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_10":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_10":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_11":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_11":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_12":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_12":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_13":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_13":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_14":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_14":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_15":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_15":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_16":[],"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_16":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_0":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_1":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_2":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_3":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_4":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_5":["pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0"],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_6":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_7":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_8":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_9":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_10":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_11":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_12":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_13":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_14":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_15":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_16":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_17":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_18":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_19":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_20":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_21":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_22":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_23":["pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_0"],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_24":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_25":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_26":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_27":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_28":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_29":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_30":[],"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_31":[],"pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_0":["pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_23"],"pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_1":["pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0"]},"pin_to_color":{"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_0":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_1":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_1":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_2":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_2":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_3":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_3":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_4":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_4":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_5":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_5":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_6":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_6":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_7":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_7":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_8":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_8":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_9":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_9":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_10":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_10":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_11":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_11":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_12":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_12":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_13":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_13":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_14":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_14":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_15":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_15":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_16":"#000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_16":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_0":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_1":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_2":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_3":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_4":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_5":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_6":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_7":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_8":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_9":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_10":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_11":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_12":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_13":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_14":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_15":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_16":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_17":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_18":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_19":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_20":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_21":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_22":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_23":"#ff2600","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_24":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_25":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_26":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_27":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_28":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_29":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_30":"#000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_31":"#000000","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_0":"#ff2600","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_1":"#000000"},"pin_to_state":{"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_0":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_1":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_1":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_2":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_2":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_3":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_3":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_4":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_4":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_5":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_5":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_6":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_6":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_7":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_7":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_8":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_8":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_9":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_9":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_10":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_10":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_11":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_11":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_12":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_12":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_13":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_13":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_14":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_14":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_15":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_15":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_16":"neutral","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_16":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_0":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_1":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_2":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_3":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_4":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_5":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_6":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_7":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_8":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_9":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_10":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_11":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_12":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_13":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_14":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_15":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_16":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_17":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_18":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_19":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_20":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_21":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_22":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_23":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_24":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_25":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_26":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_27":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_28":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_29":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_30":"neutral","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_31":"neutral","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_0":"neutral","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_1":"neutral"},"next_color_idx":2,"wires_placed_in_order":[["pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_5","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0"],["pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_23","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_0"],["pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_1"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_5","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0"]]],[[],[["pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_23","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_0"]]],[[],[["pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_1"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_0":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0":"0000000000000000","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_1":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_1":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_2":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_2":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_3":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_3":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_4":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_4":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_5":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_5":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_6":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_6":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_7":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_7":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_8":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_8":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_9":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_9":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_10":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_10":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_11":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_11":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_12":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_12":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_13":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_13":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_14":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_14":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_15":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_15":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_0_16":"_","pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_16":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_0":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_1":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_2":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_3":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_4":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_5":"0000000000000000","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_6":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_7":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_8":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_9":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_10":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_11":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_12":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_13":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_14":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_15":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_16":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_17":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_18":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_19":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_20":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_21":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_22":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_23":"0000000000000001","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_24":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_25":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_26":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_27":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_28":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_29":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_30":"_","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_31":"_","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_0":"0000000000000001","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_1":"0000000000000000"},"component_id_to_pins":{"5de9ca32-fe99-48fe-966f-1f075be431e1":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"556ccbbe-d96b-495f-b600-4f6b4261bcd5":["0","1"],"ce8fae60-c065-4ed8-a533-6f9fbc58749f":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0","pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_5","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_1"],"0000000000000001":["pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_23","pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_0"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1"},"all_breadboard_info_list":["d608a8ee-5e2e-42de-850b-40ffb6529dc0_17_2_False_685_265_up"],"breadboard_info_list":["d608a8ee-5e2e-42de-850b-40ffb6529dc0_17_2_False_685_265_up"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[1101.25,387.5],"typeId":"23db5403-7550-740c-a02b-8b3755757442","componentVersion":1,"instanceId":"5de9ca32-fe99-48fe-966f-1f075be431e1","orientation":"up","circleData":[[1082.5,530],[1097.5,530],[1112.5,530],[1127.5,530],[1142.5,530],[1157.5,530],[1172.5,530],[1187.5,530],[1217.5,530],[1232.5,530],[1247.5,530],[1262.5,530],[1277.5,530],[1292.5,530],[1028.5,245],[1043.5,245],[1058.5,245],[1073.5,245],[1088.5,245],[1103.5,245],[1118.5,245],[1133.5,245],[1148.5,245],[1163.5,245],[1187.5,245],[1202.5,245],[1217.5,245],[1232.5,245],[1247.5,245],[1262.5,245],[1277.5,245],[1292.5,245]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"14518dab-8e62-4186-8529-cb7b7ef7c537\",\"explorerHtmlId\":\"4b9fd0be-56ed-491b-be4a-ced622eda9f3\",\"nameHtmlId\":\"c3954c1c-d16c-4753-a909-3159667b6d4b\",\"nameInputHtmlId\":\"bab530e2-a5c4-420f-8a37-f03f3ef2fc22\",\"explorerChildHtmlId\":\"91752118-6545-4c00-942d-666d836d26a8\",\"explorerCarrotOpenHtmlId\":\"a0dfed3a-6279-4cd3-916a-9216c6615e92\",\"explorerCarrotClosedHtmlId\":\"596e02bb-3de1-4426-83f6-ac6aaf752a05\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"e39bec7b-ebba-4158-a3e9-e3977a78eae5\",\"explorerHtmlId\":\"1f9a279b-7cd7-497d-89d1-083f5cdcac5c\",\"nameHtmlId\":\"2ad16319-f0e5-4d17-a65d-2d21ad55a7a8\",\"nameInputHtmlId\":\"574637bf-6919-479a-aea8-e63d7b260c36\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"cb236ab7-e75c-4534-af63-faef9366be25\",\"explorerHtmlId\":\"59e53064-85a2-4465-8948-3c78b1d08dd9\",\"nameHtmlId\":\"2f2f9346-ffc9-424b-8683-d6ec41aaf248\",\"nameInputHtmlId\":\"861b69c2-a006-42f4-bc84-79375ed23cf2\",\"code\":\"\"},0,","codeLabelPosition":[1101.25,230],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[805.0076005,163.0704425],"typeId":"773dd385-6643-437a-99c0-a6e92849b80e","componentVersion":2,"instanceId":"556ccbbe-d96b-495f-b600-4f6b4261bcd5","orientation":"up","circleData":[[812.5,185],[798.57886,185.143103]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Buzzer:\n  - Positive (+) → Pin 8\n  - Negative (-) → GND","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[975.748392210648,157.22835000313194],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"ce8fae60-c065-4ed8-a533-6f9fbc58749f","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"82.61544","left":"632.25000","width":"700.25000","height":"472.38456","x":"632.25000","y":"82.61544"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0\",\"endPinId\":\"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_5\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0_4\",\"rawEndPinId\":\"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_275.0000000000\\\",\\\"812.5000000000_267.5000000000\\\",\\\"865.0000000000_267.5000000000\\\",\\\"865.0000000000_560.0000000000\\\",\\\"1157.5000000000_560.0000000000\\\",\\\"1157.5000000000_530.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0\",\"endPinId\":\"pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d608a8ee-5e2e-42de-850b-40ffb6529dc0_1_0_3\",\"rawEndPinId\":\"pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_275.0000000000\\\",\\\"790.0000000000_275.0000000000\\\",\\\"790.0000000000_185.1431030000\\\",\\\"798.5788600000_185.1431030000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_0\",\"endPinId\":\"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_23\",\"rawStartPinId\":\"pin-type-component_556ccbbe-d96b-495f-b600-4f6b4261bcd5_0\",\"rawEndPinId\":\"pin-type-component_5de9ca32-fe99-48fe-966f-1f075be431e1_23\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_185.0000000000\\\",\\\"812.5000000000_215.0000000000\\\",\\\"1163.5000000000_215.0000000000\\\",\\\"1163.5000000000_245.0000000000\\\"]}\"}"],"projectDescription":""}PK
     �a�[               jsons/PK
     �a�[�'���  �     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino UNO","category":["Microcontroller"],"userDefined":false,"id":"23db5403-7550-740c-a02b-8b3755757442","subtypeDescription":"","subtypePic":"0b351edc-7875-4477-b820-546ce15be531.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Buzzer","category":["User Defined"],"id":"773dd385-6643-437a-99c0-a6e92849b80e","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"f093df24-6efd-4d47-a863-17c5645b3aaa.png","iconPic":"72f663bc-d85e-4d27-9085-2f4219a623d3.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.39400","numDisplayRows":"9.39400","pins":[{"uniquePinIdString":"0","positionMil":"369.64933,323.50295","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"276.84173,322.54893","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     �a�[               images/PK
     �a�[P��/ǽ  ǽ  /   images/0b351edc-7875-4477-b820-546ce15be531.png�PNG

   IHDR  u  v   ��:   sBIT|d�    IDATx���}tSwz/��$۲0���Mblc0fB��3���@��0�b�!d�qN�bν'�tAgڣ�rf��i��Ճ���M�8�Ms�z��� N�`L�~��-�/��ClE�e[/{k���Y+kY��O��g?���S��ҡ�D�P�C���{HDDDDD�;����_��{�R�=�p����V)v9""""��Ή�:�t(I�R�)xZ�Q��5�cR�GBנP�@��x�1�cR��+o6I���t�|�&�I ����W��ǙM~��<>/(�^h�J""""
O����=�p���`T��F��:ix./M�8�IV�0<<,�0������ ~�}�M�Kb�J�/^:���Q��)��ӣ ]��+���!�L-[�,(q��~cP�Qx��+u>HT�*�GT�K�N�F#�0�����BN�T���@{��c�NQ9*���!�S�=�p�n�DDDDD��abg�{�aR祄W��="""""�G('v�~I�v|b��
[�M�6ן)�B�;JX�&"""�^�N�dRDO�f੅�`�b���y��A�����DF=T*~��"�bb�������_��g}� �L|v;>��f�@�|y`��6��~�PN�JU�Pث�B�GIDDD^B1��^Jx�PI�g9������~�1��y��\oo/���@�Z����80w��Y���G'Q�f
���c��	��0����'�C
���䎈��h�P�:�aLv��0�Ə��8��/�ҡ:m�Ҡ ^��٨���w��cqyX˸�˸�Ըb����q7��
B�b�J��X���Z���qu\e����MRʕP��{`<�}���R�a��A�<�,]�q��G��s"�������m>=?*v�~I��v\���H�����_�W�J�@�g�DDDDA
]1���1!����(F~�r;"""���N���);`W�*���	F~�r���`�#"""

�r�f��0e�tk�f����봯��f �S&&�ݮC�RA�R1.�2.�W,6����O�P ֋�y�q7��I��f��b�`xx `�Za��  � ��������"��<x��:�����e�?�S `||f�FGGKllRSS��!�2.�2��q�b��1:j���H��R*��?���\�e\�<n8`RG����`�Zq���ޅ��?�6�������9Z-���/��#�uB�)�o�<`�P�B�|ǟ_W*�P��D h��q�?>�v�Wg�˸�˸���B��J�9s�tA*\����xu1ʸ�˸��L���������z��c;Vcn������ݻ���|���>�����ݻHNLD�R	����	L���X`������͎/&&�y��]�����BZf&������(�k�Z���?}(��"<����8f}��6��1���F�oV�[���pa�P(`���q�q%�+�@.H]/D�q7�qCYd���fý{���ڊ�`�Ղ�y�H���%&c�}p���� ��#QJE,���0������F���`Q����b����ܩ����)lF��� 7&����q�q7Xq������˸��	���&A[k+�:��א9/��x���`��8J qJ%�J$ƨ`�����������'�=�RRR�z���.�Z��ƕ6c�MPR8.�ZZZ�~�ʕ�D�0c\�e\ƕ�J����;ר�fɒ<Q.D�q72ӟ�|U��Ʉ/._��cu��j��Q����qc
̍�A�J��]��f5z�菡/-EFF�#�"v4�=W#�x�I�ꛦ@�`
�����&�)�e\�e\�X,V�_���~�q7��"��d��_��G���I0wv`��W�1
t11xT���}�O���B{{��1"�ݎ�oa0�K4������:��d�o��a�ڄ�9��&��$�� �T���x�_���＃��nIbE"��� �&�D����(�0��r###�M}=p���`W�A(M�*H���D�u4��?��ݻ��$""""�DLꢘ�f���1|�7��SWWP�����k���gQ6��t��W��!Q4aR��Z[��#;I�� 't�X�ɱ1�{���ٳA������(0��R###�ZW�m"�;�2�r:j��qq���Z���m� !�r�a2�MY"��������(����B�sc����e��F��vxW~�kV눈���|��.
Y,�7��|�C==r�c�����~�vÜV(V��ЫE&uQ���Z�#���N��,N�D�݆�S��J�
�J���@DDD�b�@4��ݥؖ�,�Y��5O�C��`���54`�ܹ�Z���
�����s����{H�'��9?>T��A'Ʊ��ӽ~nll�!�q�qe������u			�˸�BqC�� �L����z����_H�X,�tu ���m0�X��!t~�%��^QJn
@7��C�^�N� @�MY!�q��Ұx�b�~gxxV��7H�q�qŌ+�����;V���Ì˸�+s�P��Q���/��T���/�P<�Q*�Q����,�PB��.N"%��@������D�/!!j��q�q7hqŒ��������{j�:�J�2.�7T1��2��혫���phn���cm]��~'�PB�B�����=��WU(��K/��^�1.�2.����Q����˸�x�P��Qftp�PȾ��LT
��^ht�Uj��h����^:��P(���u�J����.�			���^Mkf\�e\��5�X
E��!)�f*)�2.�70��2C�3�'�J���.���(xZεu��!�*]LLFGG���+�x�v;�2.�2�$qŢT*#���q�\1��211*����ƬT
�G��P���P��/^n
fܹ�*W /r�͆��Q��ĸ�˸���v�,�g\�e���5uDaJ�b&�F�t()X1���P�Jc�����E�ؘ�(�*Y��B��J���nΏ�ؔ�6G!""""q1�#
sBb7�Ǉ$��oʙ����(ېh��j4rcF���,��B�@A�Mِ��������])�x�P�æ(~�����w2�����:�<�������a1.�2.�J�A�<|�rیω���q7��"^9{)��C%1P�	��K��?��Ǽn����+z�իG��~��|y��	Q�-���	Ld/Ď��I����%9n����Ʉ�f~��@���ʡ
�BiP EQD3���,�+uQF����/>Gl|<F����G�v;�͐{aK���1P�Ѿ��'v،C�Û/x���ĩT�
����Qx`Re2�z|u�#h�ڐL���vL���Z�B=�O+�|Z�w쯼��ݎ(lm6�\����

{�(Q(P L�%"""����.�:�ڝ^<��>�R?O��&��		S�#Y����;�?P�v;,6;�=���P�i�Oʩݑ�8N��Z�>��  �ͷq����#"""�hƤ.����M��ۛ^=�؎՘+�ǳ`u�?�-�B�Z7f�#5�		r�h���4��� �Ä �m\���.�2��,��`�Z�����Iu46m�5�������CDD���A�{�i�3����*�P܌���۠��?�{(DS�4jԾ��-��.@��2��I5�v�PV���t�ㅙ�0���/+�'""���J]R'$ ��߃��fHU�6�s�h�j��B4E�~1����� ��q ���#;E���AY�竺=ې�Q��ݏQw���gBbW�gJ�����$�()�%i�����ꛤQ���#�����U4��`	�����I]�Z�y3>�������H�6F�6<U�W�y����6��Q�� P�w�3�[�� �a�ԕ�03�oECKǔ�7u����h����X��3Wd%��$�U��P���V�0[��kB��IΧ$�Ez$͉��B3�zM0�;Ө��ك�O���G�؁�Y}�rпk9�:6?�f4�t�� �9% Z:`�o�}��1���P����(�#'U��7�a8�i�n(5T� �T������R�π�]����Iա��է/OIn�vJ���Caf:*��(�L��A��I]�R'$������e$��b�����2a��j�!q�rV�$�؍ӈ��t�Q�|��4�q��}�^??ntK��J[`�1��[U;a�o��TI�03M�=��.�"�@W�F� �]��8V,q\��t�$/��b�����9�Iա�j�󮼐 U�_���-h�Daf:��lsܬ��.I�FyAJ�fKrq�� ��B3J�`ܽ	m�&�w�|��+�B�!$��bT�_����]��$�%yYh�ډE;O�d���1�p�ؚ<��_��B�]Q���B���)�����s~�m�&g���HҨQ��.˿CR�(ңzG)�zMh���o���AR%�rbR����p��e��Q��`�b�� ,6�J��/�"�����'��^�Ռ��x�I|��Ը��� ��+nt�>���:���˜�i��P�w����[��:��iҜx���L�<�ԫ��:	��s�*]����b�P߈���h�쁡����0�����fA����8Ū�+U�IS���ls\ؾ��(q�V���0l~ʭr"er'�o%�G0`�¸{�:{�>��ӗ/m~J��M8\+w�k~�><-J�$�U�W�����g����U��r$�6!�5�7:���F��)��5l~����`��*�^�S��*�����2�Z���|�#�%��(�����?�	]����ڂ�ؙ'&`��P��͎�+����^%vb��&�3�s����Gб�ȹ��5����h=�t�^��4���gO�	�J��=DI^�ǋ�����VSg���\����k�����f���:{P��%JL)�XP��Ǩh�pT�&�-h��ASg���sRu��v�y��1����vK��-I�vN��:��B3�o�qU�v�#BE�����b)��r;?��\q|��r{�����Ϸ���oEݞm0��$i����9��k
ڍ:�����^�O��o-��(�NH��?z	��7�@F��:����Yl6Xl6<��z}PbF#�+�l��TqgJ�H��wocw�_���6�fck*��=f��4���#p�J'֜T�E}��V���rR�n���z��
����sKĎ+�f/4;�r����V �zMn�[CKrR�S�����dm[E��9�q��b^��A��M0���V-��b��n������3��{1�}0[Q��ǎX{�IV}5�7b`Ă��U(������0[��TeMҨk7E�Ć&u�y�����������I_��yX���{�R��g���J��%vR����I��	�_b�K?F~َ��|���:bO���iHr�<����6���]mA��RwoBCK�V��X��<����C��R��e�����ݛд�nu�;J��ԕ�WjBr��Q�di�#����B3��ls�w���>V�_�;'ޙX�y�?0b�m�p�w0[a�Ќ�T�֯���j�5���0��PV�ܣS*7�a(+F�ي�3W��h)/�s~O�|�B\C� n�;oX	�_��I����Q	��N&�$�I�:*ۓ�/���(_����Hä� 8���j���~�0��+I�q��	&�
<��V�$$ub%���+�kb���5���Q/A�`�xu�t�l5ቶiH�;J���O�i��tęr���	�/��W����3WP^���-�><-�U��T �)�U�v$)��-q0�7��܀�*��.W-�u|�;���*li"�6�7����/4;�f��%VBYx��VT}x�ys	�d7w��\AҜx�t�����K�r�|��g�8���,�ñ�I���ZQ��<�B(܌��j'>����r \$�z�$�3��wl�j̍~�mƥ�%l-7��h���=Q�����0n�#&�Q���	�����{�3u%�=v�44#��[̔�(�FG���#K��ێ�1K��v/X���&i�h{mϔ��+�d��<%u{�9�	�֯Dݵ[nI�q�&$͉w�o�".�m���ׄ�w?F���:���H�`�-�3���>(���C��{��J�4'^�q�$'U7�1�	[P��3j��A����_�
	^�>/�r/l{!��TF,S���3.0��Y�~%��e=�� |�#4u��|6���,�+u�F���5�{��܌k�|Z�s���N�d�f�æV���ǲ?�C�Nn�>���1Y�&<�J��S\MW�4�����d`�"ZBmӐ�F0u{�9���0��n�6g�W9)Z�,�FI^�dӢB�1n����dO8Z:B�
�{������ӽ.�_�lǏ��P����*ؘԑGz=2~�:���q���	�qq�%%�n�atx��a�'<_H��혰�a�c:[|<����d�ȅ�{�T�gm�-���<�8����g�8�)��t��>ga�]�$_DDN����/����S��e�����`�b��4�S������9|s�"�{�C��F������v�Y,Ǹ��ݎ���1O��%6bޢEr�I�R����bb�������_��g}�߿/P+��C51Ԙ�΃�l���-�Y���ʊ�����$R�]7[�Nh�`Jw8��G�4$O�w0M6\�1���(Zp�exj�#���{cc�]|����LR������ہ�۝�u7O�뜺hQH�7�]˳�����s������ΰL�����q�g��{}&��[�M�x	ӳ�O��ݙ�����~��;�q=6�u]�S^���M������R�]7ݴ�$�ڹg��Y�S��q�X��|%U����g��d��w#�N�F~Fηv-f��'��z)��ԑ�ع2��$�Ŝ9j|��9ѹ�g��3l6qo8���0G��Wmw<�������fO��!n�(/ȃa�S���"6��tp�:�.@s�}��|+�!/?#�+� ���j/ݐ<f��'��z)���E����P�Th���x��=��B9?]U����F��U��u�~q��2�&���q��Ձ��w]!6/_��Wc߱��� q]ﾇ���b�'p���o�-y�q��E<��2<�jYT�'�ߋ�[ס��)��kr3 &�U�}]�3�P�w;��q3>��ɋ8x�d㐋R����j��s�O����R�".���_$�E%yYh���l�!eB8����$��q���|k'v�s��B�B��lE͹&�w� ���ηv:�h8O\���Z�G�6����gp���{�9g�'o:aL���:"�($T�=ڂ��J���|�ś�w�I|k���E�yM�7?#mJU�sּQ+I���ϭZ6��-���Lꈈ�����FU�WN��^�y�h�ϸ�$u{� ���,Gv�Źp�s�^
��q-�I4}/jvn��XVr�dSm���2}�պH��ʤ��H&����=�$�;0b	�F�MXrRuAm�ϸ���������}?**�b�êJ���-�[�,jΓh�^�۸��y���Bo�-z����A��8�uݴ�9��m�7��7T0�#�r�� !�}Ͼ�ix0<����q A��i2{�Ed\Wf�Ǥj��DW��+�����\�578��uT#��L���;�F��V-CG�P�.z��<����i��dRMì9ׄ-�\�.��A�h�V� &uDQ����T*��
T*�����װXş��so��I��TJ�`�"\��+H1�]����T	N �����T�����ͷe	y���,xU�h;O���z�v9���0+?8���2��ȩ��F�I]��Y>���Gg��y�wa�\uF]������סP��P�����4�Q��~�l�	���i��$g>z�� ��>���mbv�j�������Nː+n�JҨQ��9�:�TA�F��Mn�ih�@��Ge!�3��q��ͬ���nv�:�:(��z�D��n��d��|\����4�H�v)`RDm�Ch���;��G֜�ٟH>��l�|g@�a����<����<���;���6H Q    IDAT,$͉��}2I����-�v�LҨQ�g�c��ӗ�~f�oD[� rR�Ά*rOդ�s�l6/_��Ϡ��e5�=$����{hl������k{���W�'�v�8y���?�_ock��鏮-��w���Ps�	�cZ��#�:""��`ܽɹI���R��}Թ��� ��O!'U'�vEz����	����J�f�di6�:����N���e�;�1��j>B�>����?(y�h;O�����|4�~t���h����D��:""S��0[QQ�w$y~����(ң��G��K�f��f��0n���t���)z��F�EU$�on�4�h;O���F���PŤ��H���>}�Y6��۳%yY�>sE�΅I���n�lE��+n���"I�F�F͆)�N�bתe0����|#���������o��cDD<L�\\\�^4	�%8���&$Jm.SO�d�03]�ꜧ1L69��9&t��N�:[|?���X�F�,����jl""
&u!*F��J5}�>�(�ʐH�
EP^/Q��>}Y��j*���>�$/K�M�#���N$��ߢ��-ؼ|1��fmz����i��1Q�aR���P��������oJg6��9o|�	��A$�6��@ݵ[�*]��������T�_��<T�����&׺�a��ŲĖ�)ɇI]����\�+}��K]}���F��0�o�Z�aE��^�O_���%yY0^hv&�9)ZG�ˇ���y3�=���  K��L��A�(�tDD�I]���i�_���AsHT���j�JT�_9�c��FѧdV�����AT�a(+v�Y[�	��Fne �5���JN��An� ��\���D�]�����:"� 0[=�U�����-��ڂ�T�s���^��Id��f%��?�ڿ���IQDbRGD$���#^=/'U��i;ö����k�4F��i�(�]�����O��HCVr"���s]E�.���řIQ*/�C��%�f%\���3�  �]�"�u/l�MD��03Ezf�;g�q�zM����K��E��<wo���-0�7�M�2�ބ��[R}��w�֯DE�9��o�s�ٱF��n���S��L&��i{m��}�\5u�x]� 
G����d.'U��^���p�]�Q��w�àe{�9���^���Y{�#��uO@�Q56E'9���"=�w�:f��N9~I^e�(/ȋ��I&u��̕)�f�ø{��lC�ύS�����^�=�۳9)ZN|���P��U;QR}d�4.o�9��۟�^ۃ�^SD~�&�Z���qpL�du.���V�;�	n}�6���֮�%u}����)YbQ��+��(�;�a�a+���,��ن��+#�bǤ.J4u����T�(u|��8�K�P����O�]l
���v::�M��}�$/�Q�+�C�F�'͉w��Ä.��^���K7�.6E9��$�������M�=H�p�Pä.��8Od��<M�l��Aҟ����#�"I5��ls�l9}u�n9+ܳMY&""
Ur%Wf+�Vf��xS4I�v4 ���L�HN� ���p��Q�++FN�M�=0^hs�DQ������>IDDaN���x�U�W"'E����M�f^����K�ύ4L�DyA*����������﹖��VT��1eŨ(� �w����-�>}��<��M��.f딵tD�"��FE��y��Q
CY1�Qؓ+�2�7b`����Փ��-0��4"�8`R��֯D���S��D��QJSg��>�$�U����Q;�U�Q���)���g��0^hFaf:J�]e�VʊQw���QX�3��>s�g� 'U��usĂ�Ξo�"i���1��@��/sRu0�ބ$�zʖ�0[�1�><�ܾ�zG);V�������H�Ҡ�H���+��ك�w?���DD6�M����t�������$��?���+80��p���?,Gݞm+iު۳����LV���l��w?"ѳ�O��ݙυ{��ۯ�7w7Hꮶ��j��
^^����t&uDDv�K�b]3&i�0��03U��x̊"��Y$΂aR烵smXk��ܤ���VǨ#�N[�ɱ��mU�n�;۰{��!̝fBRRt��Q᫶;~�����f�˸20[�w:���7��]1f�U��B�_V�m�%$|Ez4�t����y��I��~�j��Z�q�Q�R���������!��KN��U�(EN����MҨ���P��Q��N����*F���>���	���䬘U���hܷ��ݛ`��r$q�W:�Y�E"&u^���~�slԺD�q����Ά&��#���%�F���Z���	8���T��圮�%��2s�����7w{�S(����|#w�L��4�;�W�zM(�(Z:D�j��yA�T�(��Qw�I���''P�~<ܲ�[�N	d��: """
?rW�\��������C��l&uDDDDDDޒ�b�:�L�V�(u&���� �oq���*fR��Q���h��A�ύ0^hƀي�w?v.Aj�ډ�"�dc�+uDQ���Hиw|�^���C�0.�$�3a C}�ǥ?���)��;J1`�F�>u��E��{C�J9���:(X�	s������&G�l�lE��Gg�� L��ԭ�X�#�R�{�`��ݮ��9K-D�o;��H���df+�O_�r�iܽ	%K��4+/�CE�%yY��ꮶ����.Ԯ�_�~�[�jO\�XW�(����(�c��U;a�oDCK�v:��=����F4u��j�JT���������nݼ���
�I����ԡ;'U���?���᪢H��<Y����b&��+��BҜx��MҨ��Q�/�0�#�R�rL�;U���h���PyA��BN�n�}d�d�P��h��m��9m#����^���i��䡩�Ǒ$�T�0�����6>O���7��{
�M�=HҨQ򰃢�di6�V��e�%u���h�5����L��MN��W,���q�¾�Ez��&��\���i�#T�f��૜T��>��(���sw��E��K��/����dUw�����H�r%(�LwV�\-�B���U���0-�P��hn�R��P��&A4��9�:�䡡�f���"�����)�7&'����4կ� o��#�g����-��܎���&7s�sv=��1�����%i��
�l���&W�;J���s��p͞��>���
�4�H�ހ�:""""��]mA�槜2O*��h�왶�2y/Z	chh�pTU&W�Z��2�q�a���,�v&�B�Vw�e��?�ꐓ�CÉOݎ��ҁ�<f�;�ϭ>s�y��wor����Kv��{�C (�<�j[�p�\�[ ϯz��O��b��Z'���t�i�m�&��ن�=�7$�OnL�"Шz4#�݇e"&V���sS��>�jb,�q������3c��$/u�nI:�
&L��vE�Y��Φ�H��؅����4n��U�
3��p��m�eCKJ�]�Uw��m
f��%�W�������2%U�|1��q8x�"���]O.��Gq��.��e�}��g�CG�Z��x>Ea�\[ߠ�1�.�L���+&uD��e�x��$���ĳ�p;� ��w^�,���EX���Ci�j\""�ʹ�+�C�^O����zf�_�ufBu��f;�֯DyA^@S���{la_�~%�֯t{��j�]�Ȧ�geM�
UɆ�gϵ7YCK��rVq��®���Qs�	 P{�j/����L�]W���;�]���'��|�Y�Z�b�W	��B�䛁W���	���(b}���˪N���A��;/��  ���������5.���K|��t�,y��r6Ez���9s�ʖ7rRuHҨ=&��L��Օ�e�-E����}����n��L7ƺ�-0l~
���0[��2��j��
�d�[;q�uj���}'�㍀`��}m��<�s��E2&uDL�krB����`$vL�HJ9)Zgh�!L1�JI^rRu�H�Mi,�4'~��,ꮶ�03I��4N�6�9���칾�%���.���S �����E8���:��ΔXI��1�#")��9�|�0M�x�ٱmA�S!gC[�	�~����f��$5m������kKա���?{��s����j�w�pt��$����*iN���n�ȑ�y����1a��H�����r !!a,!!!V��^zD?2fW���#���?|D�1�;����7��N�fK褊�Mb%EbǄ���TQ�G���0^h������C}#��7�:3�9m1'U��Ι��~_LO׈E��:��K@M;����w���vT��������E�>e�	d���������P(Rl6[�7�x�b���h4���[
 q
;  �_(�a�4h4J ��Ð���x��i�YG:Ψz�\V����N���n闟�������ݛ���g�J��B�W	S��+h�t44��9���2eSs_�����U.��l��p�d��:]zJRZ:`(+�j�_ݵ[���t
3�e�|���G�
�X[z�+�O���6��^�����INN����Wm�
7�Lꈈ�䒤Q��/+P��Ѩ���E��N�JK�3���,��r%"""��!l�0ymI��������������I:Ez��):peE��{
�f&tQ��:"""""�0�JQ��N�";Y+�0�����z�=�"l�s&uDDQ,?#�{�C'�P�������>�j>���.f��#J�|�0Fu:�l�)���f��A�j_������>cn]��#���hX�#�pm��A[�i����T�sASg�c�Ym�+��(/�s�Z����f��n���z0`����e��'i�0��mJ[w��������&��z�8+uDDU���c߱�rCTLꈢ��x5�t���/��S���0��03�~�|�𸡾�ou>nܽ	�ݛP�QO�e�o��
��Iա��� ��=� 8:�5u� 'U��M��a9J��` ��F�������Z��#"���5uD�rRu��Q���� ��\AҜxT�_��k�����U0^h���U��1�2�Q�~�W퓫�\AyA��P��i��03U�FSg ���C}#��l��A��7���A��ADDD~bRGe�֯D�F��ӗ=�|��I5�4j�z^�Zx��>�o�5�03��騻ڂ$����:�4'ާcE#&uDQ�$/f+Z:<�|�l������-(��Bݞmh��P�,'U���Y��03 �������LꈢLҜx�X|���<����F)��b���&)3%h���z�I��xEz������IDDD��Ѭ�VG�w?vLߜ��Y�~�Ǧ(��bʊ����T�3�ބ�Tݔ�~DDDD��:�(30b	h�����Q^��槜�T\;UΖ�yb(+FyA�����?"""�h'߮�D$��k���Q��77YyA�s����+1�7?r�ss;��/4;��4;�qwoB����x�c�}��hfLꈢL���0[QU����'o.4T)/���|��I��v��S�����?@��l�TaBGDDD�#N�$�2f+�><���{�6��SeŨZ�-Ω�M�=�>sŹ����9Ͳj�JT���EN�ι�x��G9咢Nv���Zd�$�m �67�c�\�e2[q��>���k_A�F���4�g̃N����A|��=9��u��:�(Tw�%�&GW���xSg��'��h�5�� m��q>����H��RYQ�G�F�8��8\�Y���~�(�g��L�ks3�� ����_��`ڟ5�v�\k'�o�z�=��*�F�|���f"+9q��)���i�2��8w��[�"�=��������BZF���'��t�,š�Өa��#��_]����4Ծ�Yɉhl�¾cgq��ޔ�w��d�bד˰c������w���[��6>o�k¾cg �6���uO  j/}�|�u���~��'/N;v�F��[��U���?�'/8��؂����®w��z�=d�hQ��)�O�Z�)X��~#b�J��V�|���������O�?��R�@���_��ɏ��DRQ��Ԕ(��3r !!�k�N�P���~�t7�r�(�}�5j�,r{lB��X�bUP)��o�u|jK+���bhb|O[>~���H��u�(��Κ��k�2���V�w�ηvJCj��\�-�\l^�X��w������5Ed�L���[׹%X�V-Á��ܞ����q����P�q�����p�'/�%э�](�����E�s���7p��E\��
�c<y��oLy|�����}�+�q{|��  ��������_!?c�Ǳ��c���n�����7��s��9��"��o���-n�TG���δ�����
���a��_���]n1�q�o~�L<;�����Y�7G��e���/)f��X�#""�'����p{,sI.�sf��x-!6�w����o&�P�%�ZŐ�6>ϭZ6�z�t5*�b�'$KxYɉxqm!^\[����8|x���ӨQ�s��=��������Q:n�L>W�s`Mn��&;y�X�1m�|k��Ǘdz��c ���X� ��؅�ɳ�G�5��Sn���k���@JB<�-��X,w^*�O��ޫ(Ê�#��>&uDD��AF|U� ������^��B��~��I�t��q��8��i���9�$�8f�d�}�<~v�o,
�ؕ0��d�����p������xs딤�d��d�N���*�k�s���8�ډA˨������?5q9���qJ�[���}�㞎8�E��V�c��}oʴda<��p�鷍�]n�����Z&�6�}J��쭎)cl�?�-��)�g'k����޹�N�tR")��lْ�P(*�@\\�)>>>I����}� �-�r�HU�W�_��?�el���}�G�M�&���%A�Pa|�
�Ō����A��>� �`��c�{�F�W���f�~�v<S����Á:F�?xl!��q�����_�!p$��/�������O��{�!��dMn&�� u�
:���B�~��wܞ�x���"I�ƪ��`�2��?:�������7���Y�����͆�w7���|k6<��F���.�?E��.}������څ�N�gh���X�$�[����;�L����:ׄ�'/:�ҝ�:}׻ﻍ���˨�|�ۿ�8�K���;�S����|�|kηv��>��-:�����_��?���������9�������}/t=C#h�@Y�b(
��@�q���.����Y�P(�34�m_�F�5�*�����q��&H)Z���t�����?����#.��Q��:�dU�W�PV��fﮞH�\gw{,1)���n�����I�Z@��a^�b�'L��;_��2�r�G��	SߤZ&���F�S�5w��HC���g̓%�7��%����۸zʚ2!i���63!�6g����MY;(�ף��5uDDRF'�KY�R��Xb����p��-$ν���ˠP�_��K~F��n�m��/6/_��?y�GN����D$�.��Wv��MGX��ӨQ{�\��ų���n��4�pg2[�$k�SovonŮ'���U� ޻�?+7'""�R�e#!1s��	 �զaђ����t\�R1���8�Ņ~b#�]O.ùW���N����{e�ٹa�'� ;E���
��N �G'u^�Cv���݀��Dh�����B���x�e��[皘 ������>���.��5���m�s���L�$
+uDD䗌��ߊo:�����FO����ڧ���V-s�W�dS����n�͋k����uʪ��[��(��ȹ���}�κ}>�nj��]�ۏPhb�����6���`6[1<t�c#r'(�=��3���O^�8],P�k�^EY�&t�����r��v�R��HCv��c2y<D����<u����'��X�#"��d-�.���u�:t����=$�H��]���e�}��kr8��J񼷗?��q�߻e�?�uk��!�{d2[q�ս5���,L�B�-�    IDAT�Q#?c�3�DM���P_�]Ҫ�������{���P޿|��9�2��^���������?CaSw6�!10�#""�`||f`�L`��M����3f(�\[(j�r���o��ý������5��آ_�2�d�J��N�.�׻��K7P����_�b�G��y�ٹ��9�f�k�2�=՞[�Ǜo#��oI��Wy�*�����\���Jvq�ܺ��s"0�#""�%$$  t:Gu�61�ί?C�|xL�l���mA����8 B���A�^���.}�S�⪣�_���/߀6>{�=�]��T�4��iԨ��.�vR�G��|{������qp�:Iײy�0�g��N�$���4����I�F������jo¼�Q�5)��a���m `��)F�)ڀ�E����ɋ�iWb����ɋ8x�"^\[��W�=�0�Į�bK�	����[��ֹ&<�j�o\�wr���B�k�,�:�b���'l*��1k'u�l���}�7<������{���%v\cG�bRGDDS(Uq��O��wU1j<�Y�{�����;�Q١��nj������lE͹&<yQ�QM�hm����k�:�?�]��nS}e2[q��E�6�Ry��c*��uO���B��X��=�6(�i�صj��sq�������w�\��qn]���f߱����t�cp$%�T,'�^{��hS�3�ܶ��vL3Y�����
g�B\�o��A�(j/}���8���#�pp�:d%'���7�wg?þ���{�*|��%""�hS�C��sal\<2�W  ���a}��v&�h�e��B��������~O!�Ǡe������V�<�����6>5;7x�$Ц(�ͭ�<r
��Q���+��y���[|�lj��pp�:���ܺ���.���oL����in窘�b���~}&�^1�x�mQ*�:�:��	�����	{���O^D͹&����7�:߇5��h|e��gϯzܯs���4 "� ��b�͏<�W����q�����ohԌ���qv��C��6%���KG�Qc�������K7������йjl�7j���Ϙ�ڊ-3>'��1B��yc}P:W��]���;~U�6/��)�a$l�1�����E�L*���+�� �۸�����"d�:��zq�I����J��0��Q���z��;��>�l������ߙ�L��G��;�T�o\�״�}��e*�l-��R�+~vv=�{� t��4�mד��n��7�]��hvٚ@.��Q���{}�?�u�(��k��Jr�E��W����bo��Ϙ�׺T]|�$�������3WP}�J���f��ɉ��I]��N��E?֥U9%z��@������ZC�1�c���~��z�=��(�!�;��.���f%'bד�^����'8���?G���x�m�+�bp������o8��:�2;E�5�����=V��Y�z�\�۱�����:""�Iv�q���ҍ�K�B����Pvx׻�!?#�{��U�ńN0h�.�q�Wn�ij���E~'ukr3�������T��P�,����uX�F�,�����޴9��m�;vv�ϡ�o�}�f&kr3Q�s��ݞ�˺T���nKͯ�&wLf+�:�aMnfT�8��#""�d�'|z���N�� �7>x�_	�p�*l�i	����>�إ4+9ѯ�ukr3q���۸�6��?���z�x5Á>c��]Z�Ө�ݢd�����^�[;��Z�S���߇�(�[;q��E�X�����v�|�_�ŵuaH��F9�2�#""r���e>%.Bӏp���S~��g�õ���k/:���[ס�r�����1<����)����^qͤi{��8����f�9���Em[�y�~����_7=Lf+�j>�ؽ����)Z�)���8���[o�|��H�����c���ɋ�u��G�SA[�c2[E�н�p{	O����q:�&蛗/�����]+�pv��gn����I���ǣ�S�����y�K��S�6Q	Or$vLꈈ��i�3n<<Y{�`Ht��Še�GNy����f��e�C>_���?g ��������>�o�t�pt��k��E��!f�)����yڭ'&��c���V-�Zw��ޔ��q:��<���1�#""zhMn�O��bP���%�2���ِض�N^����VwMf+�s��yc=�7�c���'١�Se���uAٻ�S�x������K7<V�}�Z[V��������N�&�n��`&vLꈈ�Z����}�!���'>���)�P�ꍎ�!���r3`ד���k{���#ܺ.��� BE�}����D��)��L�;e-ݠeT�
��)� ����{��&�O^Ĺ[�x~�㨯��J&I#X��:""��|�8��<�����s&�}����{>�/��8���4j�=鲒��F}s+NL�����P�N��n��7��^!��p3#+9ѧ�)e�\غιf�����7�!q#�cRGDD��/�߻�#	�}�>�qJ���n�''>�������OIK�6¨<2�<�n�1x�as\�u�&�����Og����2��Rh�:����DDD�|�=���A�׋��n�&����Lh����۞�^���֮���7�M~F��]=Ϸvz=�-;y�J���Nt��mV}��-"��lŁ��.�/���XG�醍��Wx�xs�xޜO7�K��{��a���*�>6�:"""������rm��E���7����h����ـ*%�u��V��͹W���g����+Q8���uR�671��]���﯆.^�s7��V5皰E��b�*������ۢ�5�tS��H��4��S����8�p��/o�k
�6$$=�;N�$""��)Oӹ�g�N���ߓ�/��r���ـ�]J���{l).�u5�u����Vv6�c��+)�����K٠��/�}+��@V�܈M��)�e(�I1�I|����w���x�N�ӹ����M#�2}.�W>�}W���u�����"B{���je0�����J]�ߚ���sq��]���lG�{Q�&2$�;&uDDD>2Y"sO����~U0"uj�/�G�ur�ٻ������y�X����5�b�]�I��k=}�&o�0��[�9G'i�����:"""r�Te����Q��Gܧac�P6�&�/�y)����1�#"""')׶E�Ó��5�vEl��W׻��I�X{�I�EJ���N�׏"���:"""��s��\�ʛ���ͭX�s#�����BY�GAY�8p�":�ݛ��1��S%y�[����]��8��m4�v���7�T2)���qK"""�g���������� �"l��c�_��&7��/��0�{����u�ZG�д��}o�Y''�J~F��s�Ө�����-&3���<r
�+�q>&��uR���[�0Y��o���F�] �0�#""�o��z��Г��V����Zq��zr�߿_�s���������4j|�ڞ���_�z�����WQ��󾍫a2[�*a����N���66/_�|,н���F�씩7|i��Өq�'/8�4��������E	;N�$""�o�n"m��6>5�6�M�Qc������ƛ�F�^_��y�`&;yj��E����|�V9�vs н��F)v�.X�a��/۠T�-t떩Ϙ�]����B�ǟ��Lꈈ� �6���H�Ey(�ٹA��ʵ�(�db�2��ٟ���^T�<%��C�r+'�ي}�>q{,н�<M���ٻ���;��H���e!"8�Xp�d0�f�T�2"����=A�dfrj5�����`������cMrƐ��(g-r	V0Nl.��E�`ld���ڒ��R_��;�����[?���r�~��<�H����<�'Q�wK�_P!ъ6��  �"�bf�y�g������+�,��mј�#X+y������ӽ:`Ц��X�t��e,�^D���'��x��We4��Eya���F�;9c���P�/��h�� �+����;k�~�"��Ƶz���*��灻�g*<r��:?ҭ	��P�7��;^xY�O�;��������|v��dT��<sf<{�S,����7|�p�$;�����=�Ԗh��Ǵ��c������"v�:  �8�L3O5�)+�k��BvݺV�xP^F�v�yh������*~�a=s�����zC>�Gό*���3򔌑:i*ܼ��3�źw�ۧυ����|5��=q����w�=֕�ЁǶ�ÿo�-�Wh��"
v�:  ����}�����0Wm���Ѝ��<pg�ih�Z��f�7��ĝ_��o�ᕤ'f��3 X�蝹f+/#ݐѺ���z��>l����9k=Z�{ׅWO���
��.p"M}mF3���c�C�?��zC����p�`G� ���'��ւ���I^F�<�=��N��h��%���myံ��i�?[^8`�3�����Ϳ�k̺�x��4'�>�A�g�q�'"�jj��oה��4�y��9}oe͠ue+�Nen�<�(�����k�`G� `�h@�����*��{]o���L�ڞ0&�u:���sa�9=m�C�Dx{�F�9����!��}�v����F�֕��3�6�,�軤����/��3��̙��W<#b���ٜ�	=3�0N$fO5�kK�|��P �4m�����i�� /}垘*]:��ㅗc�s]�
Â]����Q.	�f����HK���~L���-}�7�nH���_?6�㼌th�mT6���j�H��_?�����;��>o\S�[W�b�F��=�ˣQk���hb��hԡ�C�`G� `��_?���n]kȺ�D��;j�+��x��ԉ�K��r0����6W��z^�륦k�<=�n��~����������״��A��������"��W��{oW�_�3���N��hǈ�3gf��ٵ�`��޸Vo?�+������S���#�{�o��b!�5Uj��%=���k���*������I��
��l۷o��X,�jPzz�HFFFA�������1����n 9�ׯGn�|T?`�}ӵ:;�S�a1xx�Z5��ӵO���P�ק�O�j�>'���}�����7]�W?�X�/��$JMY�~��;��f�꺽o��_��l���u�Z=��u��Ks�tq����>�=��>�{n�TinV��nS}M������ڕ�.-TEQ��33��ժ���#�~^�޻I����-U�s>�=C���r0��ݖ����{'㪜�=�ԵEya���F�/�^V��3�uin�vݺV�k��۔�f׈�#�קue+t뵫����ڻs���s׆�{��ׯ/���G�W[�����>���<U�j׭kuནQ��a��H��?��:���Gkt�z �L<��Q����c�o�lІ�Fx�+��<B���:0k�ቾKz�翉�o�?���~�E~k�Jb��tOD5N~��g�[�f��Q��Wն�Ks���e������z=��=�]�.������R}MUܣ�������k�J�|T:��U��ը�jK��Q�o�>�/,WF�~	 @8�=��}ݳ(�h��H�+�9�;�z��Ԟ�V�+[���_ZU�btRl�fk��̜j�oP#좩�:�ξ~տ�ꢙh�4Li��x����%�k��:�I
{~���|X��a�%�<�_�Չ�~}m���Hm��REa��>����5e%:��v�}ӵ1]����O��;�j2����nԺ���gS�Go\���ᾘ]g_����1�~����L��ghT�>���rm��ڶQEyq<�קW;>�ۧ{U��PuiaT���������z��.�^��FO�:uqHwT�Ϩ����麇����;��y�1W���?����~,��-U����Θ2��{'����bj�/˾}��V�T5 ;;�l~~~l�u�<��N�R� &�̽���*SS�JjY�x�+MM����bL�,9#.����[I������g�rS�{�9�	�j��%m�6���;�~���Ж�r�++�-�W���y���:���^C�_EQ�*
��N�]ZS8�SQ��'�U}M՜"1�t����̙��-U�:��v�e�����W���[,��0B�<B�x��a;Z�=��_?jHI��l�Z�}_�'�}�b	,�M�g�ߊV��SϿ~,��Έ>z��o��C|$����3>v�'T���'�YXغ�Z��dF(
��x�xlFp�պ���|?�B)  \Ů��z��]��>������h��I�t�C�����z����W�-���
sD��(O��G��{�^:ܡ��ް�N��V��{o���^~�d�]8��> S�e�1��oI��� A��a�c����k�D�%�u�����1��U����J�7_רS�S
������v��ۧ�E=ʹ�0�J���1������^��{5��,d׭kC���	}󧇴��
U�{ȩg~�֢�����+[��L�N�]ҁ��3F�������P�%�P\�#�tך?�������望�R�����ŢQϤʬ�����������d��D�����=8��!��]�᪢0O��)?ӡue%q�6�f���L��<pgB�v:������#ij{�[V�PEa��T�6$��R�>V�uh'�.i�C��X����5}���=���?���z��	�0�/$��;!��`���4����nB��Z���2?}l�IW_��5.�<�H�J�sT�]���옟c�Xd�X�i��б��9���co{2�軤��^5<�m�*��pF�����vEy�(��at"%3�IS�58�rv�x�u"u*��f/��H����v�?��g��7�r��ict��H֬r���d�Ŀ����gҫ4�'�j�ߍ����?�G��0��A��x=��H�O�����jo|(�s;�]T]�+j}�A�U�QS�5���
2jo|HY�k~E]����}���˞�#) �,�H�W�#�u~�1�R%Q�.�^��v��FB���W�����bڠ|1y���)A��SL��(O��{�*
��o��>�k�����:�w)l��p�G5��U�r�������{����g���{���W,�=c���@@���# O�P��b�U@u��'�-�: 0������oPS�fu����S=3^o����,�W�Oތ9Ѕ��9tV�.�QFf��)�)�[|ۦՋI0�xl�)<���pGB�q�ݓ:��o�>2r;�X=���{Be���[j���Pn�Z��¼�7�Gb�^���7���?c�����ڦIϰ���~`O�UzF�����R�q���X���5�c��O���O�z�Ԝ��7�q��?���"�=[�O;�W���u�����KW���-�/<��EO�-ȵ�,�@�EJȲ3B �Hǹ�*���f~��Ӱ�35J�s���7�����k�[7��z��O���h�!m�Xm��3%I%�*��9tV}���▘��L\Y�d:�wI[^80���b��ׯݯ���}��}4{m�b�!���t�����Ӫ��im�*׉�KZW�bN@���\{tL�n]Z���]j�y����e�k�w�~߫�փ���K��&<����I��ǆ���#�4��{2d:����g���뫵c}�Z�ר�'o��~��j�'�%C ���,����j������%5�>���b�6�u `2-G;UW�F;�W�y�65��MՖ���~��F����yNN���^5�xኛ�;ߩ�K��h�u�<ˬ���w�Q���3��YО׏�dDg��Ѯ�U_S�=ܹ�G�9%5o_�������ۣ=ܩ�����-e+B����:�}�o����GN�jW��9Ӳ��{�Zo�
�W����5��jxxX��.�ᰫxE���	oC0�u���h�%�[7�q�F5l���x�`�t�����n'�k9 ������l��F_x�EO�mͳ[�,ғF�S"��)�\æ�?���͡���fW|�Z]�=���ߑ=-]EJw��n��bY>�)����ۧ{��;ݨ�����K��gm�����s�}G�����j=b������E0:���A�^~�d���=��yL��~x�ywG���،-&��	�{n�F\�P��ٕ�?|����Ј�3c����B�XW�B������p�{|�����*=q% �t�#������d�    IDATu�Z=���q{��/��F����v�QU>���!g�k>?ӡ�wԆ��{��A�=����O]��������Lӛ�Vk�Ƶ:r�wƿ/����S�?]o���3U�����\Ymv�9/�\��UPP���jY,���,;�W��zMh}�l͇ޟ�~�?�Pæ��3[��T�Ԛ����>�:��.�)c�V_|j�)5�|co�U��w�&��	�<jz�jy�>�>����o����%��b���Z��z䛼�1���̑�jU 0w���D�%��{U�n]�g�ݔ���>:������,#.���~L�wLMI��Ji�s�'��[�jM��W��Kou��;qy�tO��G�{B�5��XÕ����w�N��N�vb������{u�T��U�umQ��T�Y����_dL/��j�F\�}t&��	�軤k��gs�jm��SI�s���ܢue+f��RU�-/P���Ϩ$���\�ۯ�wԆ�o����ޫV+?ӡ]���V� �1����{�O�5��j{�Ka�W޲z�v��S-�`�
K箅��[������wy�Z���Ӧ���z���{~�8I�����ڱ�zN�kj;��G��23���w��uz�᫟��~�5�[{��~k{��.��� ��h=~*���k`DMmG�ކ��J]�N�I��^�vISB�=�_O����7̎��=���;�[�s�v�?���t���=�_{^?��~��?~C����]Љ�Kz����tʗ��`��/�����go71=��>o�u|��V�	��k�TQ�7��#��ծ0[\l�Z�-aF�wm\��53�`�e���0O�gmi����ue+tǬ���j]ي9[`��^�k>�aij�qKUy(�Mn�鰇�|^v������E8�7�5���]�=�Iψ�3.j�K�50r�"&�~"Ia��I
��;�ھ�B��������}��k������� ��*��UwcE����	M��e������}���'C0�m��ӄN�
�GZ�T���k�+o�|�e��#w��)Q/�Ow���=�I���1m����m�茜�ۇ��u8�����>����u|�J��3��{/���+����<a��=�Ԉ;�}f�]��.�uI���z��M�}��՞׏���j����[uy삡�-�t� ӡ��]�Ѱˣ����V�B`����eFH#�G2]���>�ᗿ!�{0� L��������Tæ�P��. ��Z��e~}�{R�%��ͻ&imX��>}nj-�+o���JwTMM�="���Q�軤{/��ӽ�v4.Z�~���#�u��aG�"�tO�����a�%�u�IZ��T������-/���u�	��[%L}���g��qy�ďߘq<�����;Bk�z�FC�ئ�������{d��C#d�}����ȭ��}8r�W�=���33�����I�軤�_?�-U塯���P��S��r�x�==��7B#fӧ�N�{�k�v�릿�g~�������N=�ũ_���/���J��^�k1���U$�?���)+w��3c�w*��ڎ��z��nP��݆O�����y�.Co��~�5�/�k�B �PS�fՖ������t��M5j�����%�~�?��m��Hekn��s�9��V��V�#[nט|^��F�~���p%�}��� ו���Iq��3�O��m�EX*�jN�]҉�K3ʾ�*�_���<:����S��{�vzi[�i�{�\hs�`_x���:τ=���^U��8�����K�;TQ�7�ks�+o��׏�9^��U�+[!I3B���9>��h��������R�=�{n��\)|�'�.����{|�s��~�O����zo�{ZJ�N��is���3���SZUPF����;��L���݄}���B�4��)���O��f셧Z�a��^S�����:B �L�7�]#�@��YW�&T9,�i9Z]�Qc�^��=!ɮ@�+�-���IҤU�u�O�ե�C������42�*#.Oد���wΝ����FL�;>�ߍh�'��.��ْ����K��>�Ν�@��(�`�q��ר��t��\Fp�ѷ���z�ڱ�Z�[7�ն�<���@��ŧ�O�m�X�����5u `"�������4�o�w=B2X,6��W���MZ��Z�y9r��]y�*i�my  fc��U~�t�����+��5֫��Sr|����l�E���;��`�Y	�׆G��x�Oޜ*f���@@?OŴ��F_x�%��)�: 0����?�@��Ȝ�d���Q��g�TKs�++�L9y�dO�Qzf�` H���1]g�ٵb�M��s]�kt�3y'���M\��i�[Ԗ����9�k�[7���!U�ݣ.�a�'��ymyiT�	�o��}�D{�/�$�nm��F6[pyp��|�E�b��]�:#�$t/�ͦ�K��
 �Q^����^���Y�Z]�^�44����S�P_��}v��gj}�����WN_'���������F��9uk�f�Z�-i~kTSu ��4��w���C�G�bY4��e�Q8s���>Y'G��d���2r�W^�_���r����'$���� �����ʟ��V����r��S�K���l�Z��R��oC��?Sæ�9A���)�~�ID�.gk��k����y�uF$���/6���>Ց��G�)�B� 蛿����v  ���Pqh��O�d���ҭ�Ϻ�d�ov�+���ۡ��٣���W��Ψ�y-��Nijf��A��'P���J���e���N�   ��o�98��')i�Y����T�a�@@B  @d�wnU�j9ک��|Ֆ�������8w1��A��P�  ,k�?yS��^h�W�7�*�P��Ў�Ւ����k��Eiܻ��_F;zH�  �Gp�dI���"�R� �l�:  "P����?}]���uu}���T燞o�nij�)x?D�����H]æ����Xܲ�Muf���uQ���f  ��L_s5}J��a�G]#j�߬���<�n �A�  ��~�g��f�~�G���
���T7�T�O��q�F�%*�Q�d�X�=$� p�奪-/���~Iu�kTY�0�`�z KK�*),���t�4  �*��r��O���Eu�����R5l�YpS\�K��g|<}ۂ��fǹ�Qm���P����������!� �G��5顏�'s4�cW��snN K9ʊ�A�F=�*��:q��y$��%Ip=]p���������M5j޹M�z��vD�;��F�Z��RÏ~1�܆M5��;�]T��筴���y�R�^k9�*�_W�F��?8����FT����q�5l�	�D�<j~�9�g���HS!)�`��H�9�ػc쟟jMu[$��6D}M� 0��֤���B[s��W�y��*�,����Ue��(-;��X,Y,}�y4t�du��e���r;�WOU�tyB��Z?�DM��U����d:���}3�Nנ3���6��-/Uˣ��dD����T�,�t��~��n����v��ᦢ6n�0��'o2�`Q���E�����: �~߄��㲧�H
�/�2����5��f��$I�w�*v���T���h���Kp���G���G���Q������7�	{�VY����|��TS��<�,�W��m��^z��p;=��<jj;���ҩ X�F�;��� ��X,z����JϋOu���O�m�(����R  ���:����х�?�u��ώԨě�uA뇟�x-P")���v$t~pM^A�C��6J�褩i�;~�3u$Zjp��� ����BO�ӧ[����f�ێs��?M�l��ϓ�  &��%�xro��bm��RB �X{�C����io|hΈMp�g�f�M��n��?}=��*�M���;rUZ�N�׮Sz����a���N��|m��=�(S��S��s��pU�n�}��|o���.OJ�,�{��
gӿނ���h���a��8F ���b�]9�ػ#U�ϳ[�b��u ��Ֆ��Yw�~�G͇ޟ�*����\���q�b�HF�r
oP~�-�)�VNA���t��*\q��ӭ��i���,���٦����p#n�Ey��F����:%��g��CA�#�j���f�����*kKַ�&}���o��a����z���"Q��~���`�kܺaF�hj;Z�4�XGA�#4:��r��׬Յ�:{����UPT�tG��v�,KB��l�������
����N�,9��^K������_v/xn��{�0��o�Y[���:���p2������V|S?��E��'o��TO�����$��~s���TY����#	�XlZY^��kV)?7Sc����Z�η��(]�� ,N���٬�zroA�������v��=�i�A���	̷n���E5�QS�f5�ܦ�㧴c}uhzf���W�f��y갼^��m��iF�R��T�Y�[7�
�DZ�$x�|�۫�v5��>:7}�n��,�G �.����p��Ou$�9�ػ�귶��$F� `Q���-/U��H��ܤzz������v�,�����^�ˋ{�H���¯��n���lAܫ���t��Ia�x�����)������0�E��~k{���k4��O�-��Ƌ�6YfD��u �ht}��9�/���xhZ�BO�����{I	
rd�PY�M���I�:/$�ىڛ�T�UGނ{�Iх���B�nm0�|����)\x�Jiz���BdS�fISm&�0��o���=�b{�7���{�ܧ�6�٭�E	�P �\���5������a"�k��~�&''599)[Z����,�P�z�vh�3.Ir�����}Ѕ�?�;�pQ�T��7]��eO/RM�N�mܺA�;���Xmy�Zp�)��+f7jܺA-��q��r�30[p�{��`�kz�Ii $�Ţ���{���ܧ�6D�������ܧ�ט�����~�t���cM ,ӫ_�X_ڬy�=���@װ�&�~]������5u���rTV�gs��|�	Ym��y'd���3��j�Hz�����t�i=~J�WBَ���/�r�S�5�o}�k>�~�Ѻa�G�o�*�����3^�0F0c1���G�Pˣ���8_�;���q��� `f���zW�]�O���@@����uM?���Z,�JTg�h����}�: X��S�ZP-�ާ��aGꂁ@���9����u����b�)7�B����h��#��s�5��Ž���Q�h��CV�`J��z_]�N5l�	��u��Z+9��p�u���h���צ���8wQ�����nPæ�ｩ�Z?�$��1 `&��Xt�d�;�1��$}˳�۷��j�J������>���o�$�\�g:9�Ju3�����Z��z���4��}5���Rmyi�}��nPS�fu�����9��>���F�mGB#s�jԼs�T��W"j��}�Jݔ�ٌc���O٫bzO�M�����^������ׄ{0�z�d�������  �+���"�|���u���`�����T��Ֆ��=Zc�Xd�Z����U��5�/�I�E7�jK��M  `&�_�"���7����6ը�T�Z�����2�n�������oPæ�?u�i�N_��kg;?�urT�Mv�-����z���eM_)Gza�kpBҙ�� �rE��E�k`$�^���?W��ݡ���~v�װ�35%�J�pS7���/Å�?�  @��Kk�R�5u   �ǚ:    01B    ��    L�P    &f/))Y��������8��=K_q�D�   ,Q��   ���    ��u    `b�:    01B    ��    L�P    &f�t����1U���^��>UϏDFFFaFff��?�����⾧;@�N�7�M    ���/�גnJuC��>���������z�����O�    0\    &fOu ,]��"��ޛ�f   ,i�: 	㷧�U�2��   XҘ~	    &F�    #�   ����   ��T��@C�o3�*=_�P�j��G�   `g?PqW����Oߑt�a���    ��q�u}��[
�.���wT8h�h#�   @�4nݠ�m��n)� ���   @�d:����*��P���Q]�]���P    �wn��e��ڎDu�RtA�;
�    H����j?��5e�-�@T��;�H�S�9�Q_�H]��Ҿ��6    fm������d����:B]n���Wz/|��v    �lL��P���5����:9�Nus    \�V��U���7n�G�'���>5�E����f����T��^��qѰ��F������댮R   ����1�S+W(=}n����ٳ�
������46��ʕE�?�T�~��ϝ�P   `	����a��:k���w���+Q��ΟTaav�����$���    ,~������y���|��~6湉t�R    ���   �T?�E����0R    &�H   �%��%τwƱ4�_��i�}���<�3�kKK�s%B   �%⓮:qp�q�զ��I�	X�t}����<ע�Ң�<s�s�    H ��:I��}�8,�w2��1?�2��zn@}���O    �����#8�'����3#�>���:    01B    ��    L�P   `Q�_q}���4~�M#��b��P   `Q*Z���nKu3�o����wk"=+��	u    ����t�   �"�T���N"�   0���
t�   �I,�`gd��$�!w   �$*Z-�6�\:�����ut�   ���^T�k$�͈Y�ؐ&�u    �������+�͈K��H��ʨc�XS   ��B�����r/B   �Eo)� ���   ���]���P   `�Zʁ.(�`G�   �(��~��]P��({l �k	u    ���T7!��Ƈc��P    &�>u    L�s7��]��d��o�n�:O�׻|j���F�   `j��4�tj����ύ8�=:{�W���S���u    � �ΟVaQ����!��w���+1��R��?!�   X"���;/��?��?��f�
�    ���    ��u    `b��   �d�����8�f�+==mI>W"�   X">麠���Zm*+-������熞�л   @�Y�7XI���S��ay��K⹳1R   ��>>}>��|RO�x�l��   ��1R    a��7�aS�
2�Q뇟���H����0R    !�wnS�����sU���ƭԼs[�[��0R   �p�5l�Q��Sj��/B�ZP�j��vD�.ς��_q�r����ܔ�[m)\ӵ��   0\ݍ���?	vy�z�Ԍ�2T�Z]�ݖ�."~�M'o�[�Y1]O�   �4]�Ψ�_��.�@'�    ,rK5��$B    Xj�Ψ@'Q(   @U�i����;.I�w/X<e�h���T��;	ik��$B   �j�����"THe>�`Wr��K���m0,�I�:    	�q��5���h�V~�Gu_���G�   `���5�1��g?Pq���M���.y���[}�!��P
    SX
�.���p�א{1R    a
2j�T��?Q��H�X㶍��^�a�G-G;���n)����/�]Y';B   ���-/U��� ӡ�Ag(Ե>��j�KC��U�QSQ޼k�b�2"�1�   @B�<z�$����?�$5nݠ��R��T������W�q��mTA�c�=�r�������b�    n��jU�����|����su7VH�������P���4���z?Z�.���w�=6ӵ�:    �N�l9�:V��P]�u����))4�W��1��c�Ih��5>�u�:    Iz�zRܒ��B)    7|�-I�,�m*�c}��?�������nX��6W�f�?޸�u�<�w?�4�g,���F�   `��h\��jz�*�th��ju������.�<@s:�re����F����=۫@�؉��z�l�:    ��8wQ-G;հ�&4'MU�j޹Mu�kTY��+CL    IDAT��������u���
��e��Q��[~�_�Y}����	�   @B4��Mu�h��j�<j=~*T8%8B7�����3�^����;/��?��?��FI�s��    $L���n*>���G�P��S)h��B�K    	S��PS�f�U���Z��j޹-��#u    ���T-�ާ��|Is�T競�T;�Wk�~皺勑:    	Ѽs�*��`��ޜ�+����vD�5��f�3�]�pi|Ɵ��IC��+1R    �ר����EP�����5nݠ��5qmL�I���88��jSYi������zNB�   `Y���B�B�.,��&Z�V�����wqX^��#g�z�l��   H����50�3>>}>��|ROo\�Y,ϝ��:    ���`���ω$ b.B    ����X_}�s��P�26�:    ��8wQ��O�q�5n�0�y���O��U$e9cM   ��h�ɛ�,�WS�f5l�Qǹ��tJ�*��T[^���|u�����6����m�ڏ~%�ߗ�'�Ǒ�K�T�t���,Y���[g��P��   �IA�C��6j�-7�Y_�50��?Q��i��	{}���%�<�l���ޘ�'�E�P   �'82'M�H��-�`o���~	    I:�]���Dz�N�|��vF:�P    
2Qo&��q���0�Z�3*�I�:    	Pwc�Z�/�k~��?5��K%��$B   ��8wQ͇ޏ���	����bmZ��Z�r>J��R    ,Fl>    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01{� s����5=�RZz��2?�_#���T�   0�q�8�У���T7e^�/_V mT"�  `	b�%�666����T7#�˗/���?��    ��:bllL�������������@��   $��SZZZ��2::��&    	G�ò�ZT�e�l�,G�N��   +B���4�ʍ��YRR�����a�   bE�    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &fOu��
3��ސ���C���ci�����|�c��n  �]y��+�R݌��,�zzc�k��
=���X
c�����f  `W��T7!*�:,�>cC���   bŚ:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� �P�f�Ck��_Ia���/v?    V�:,�t}�q�%9��   ă�    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� ���Kg\~����v/    �:,�~}�g¸�\2�^   @�~	    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���S�  rm�Zlܗ{aN��߳#��   ��n�������F\~C��?i��%�n�=����\B   B�2qflB����o֐O��   @�XS    &F�    #�   ���    ��u    `bT��i�|>��n��~�l6eff�b���Y   @R�`J>�O���
�$��+�׫��\�   ��_�nw(��|>MLL��E   @j�`J~�?��   �RE��)�l���   K�����)�u�oZZ����S�"    5(�S�X,������D��%�   ���e�X�p8":�������۸�|θ{   q`�%    �#u0����R݌�ݮ���T7   H(B1>>����T7c�ϧ���T7   H�_"n�5�I���S�    a�C\&���-(UAIy��2��_�Y��n   ��:�er�u����W5��    	��K    01B    ��    L�5u �����A����n  �p\��&D�P ��seU��  ����K    01B    ��    L�P    &F�    #�   ���    ��u    `bl> �jJ��o�ָ�:����g:�t/p%¡? X~u R*7=M5��r��c��e�m)l�yџ  ,?L�    #�   ��1�@T�\�*�՘˘�YΡl��������\.��*��D���ONhrx@���2�{%B�k\�?9��˗��Ŏ4��o[���CǼ^�F�n����}�I�Kc�C�>�x��  ư���r��VZ�����+*��\Y�7�\s��ۍz<�(���u�~-��-��<E7����ؤ���T7e�  a)��:��~(�m����T>0���n���oVVV�$���L�C.�K����$��ŋq?o��d�gFF�._��,� ��lY����<���'�===��'�a��7���v�r�-��?�3�p�*//Waa�$͘&8��������&&&��ե���9sF��c
&�%�,������ٳg�D ��-�PW\\����<��?�?�KA�$##Cw�}�n��v�|��r8��H�|>���kddD:y�~�����O?���"�'  0��`�C�xV�������l|��SFA���Mx������!MK�XȪU����k�ƍ��Ϗ;x,dhhH###�����~�;���Gt]���	  �Pg����r��p�je���z�r�\���]�����٣_�V2��4��U�V�G��͛����@ ��VNq�\�������~��_GF�Db��G}T_��Sڟǎ����z� ��Y�.Uk���Ҕ��-#u���x4::�����s��r:�S%�P��&�dggk���)	s��\.}��gr:�:x�;����
"�'  H�e�R���D���JKKKe3�˥��A�^�z��������'�۽dB]��n�����׾�5egg'tZ`��N�z{{500����/X$�A$��|�ǔ��C ��-�!���C���EVV�#u&�~�����y�������D��$�.q" ���z��'��C�f��t4)�á�������v[(��SPP ����ߖj�4�����	  �[�i�P�x,�Pi ������|G��r�|>_[�ժ��Y,]{�*++����Þ�� B�  H�%�6u��ru����K�>������h�|������)�á�7�>�����"�'� �d�,#��E@�mۦ��~ZYYY�	 A999���T~~��y�egg�=���R��O���b~��'F�'  �:B��E@�|�ISoϑ���믿^iii	"��\;  ��	���������T61p���ʕ+<���������Ą�_.� 2���ҙ3g499�={�h||<�y�Vq�?��O  9B]�|>edd��΄&''5>>����ϛ�������7U��4��]�V��������$�.�Ad``@���w�=/� BN����VSSӼ��  H���b Q�$���g�UVVV[����*++Sqq�{�y�N�����9՟��'  ��X�2�� z��'URRb�"�*,,T^^�jjj�iӦy�+..�Ĩs�{џS�YXXhH ��� �q�}���n[������L��k׮y}a���5�\#)��	  f"�����Z?�pؽǖ�ͦ��2����'�H�3�[�Y�&��	  �"�����򗿬���T7%irrrTRR���r�[���{/�����LX ��u B6nܨ��k�O��k����Z��G,�Oc�  �G�K �Ͷ$�X,Kv'�e-##C;w���MuS��f����D^�W�a�=�Oc�  ̏]��b�hrrrɭ��Z��X,���,��V�|>ߒ�����jݺu���HuSR���D������ׯ���G۟  `~��
Kr��|��n�+==]�E�@@~�?�-C��v��o߾,G����K###ڴi��=��Oc�  ,��0�����˗5>>.��#��*�����5�\�[n�e��"��n�q�q݇��bT ���>�/�$��jbq����+�����)������<]w�u*--��>����  ,�P��
r��r�\��wX\���USS�$�
�"??_N�S_��c����)��  W�O�H
��/�˥��IF����UWWS�押�<�|>�_�>���ϙ��O  pu�:$���._����ȝw޹��~Mg�ٔ���իW+;;;���ϙ��O  pu�:$] ��c:fj��v]{��Y����v��nݺ���?�������X��	  "CiB�������f3������:+oKQk"������J���Ѳ��u��]��Q_G�k ���R�gI;�ͦ�˃�nF�


�f͚e�A�|rrr$I7�pCT�џ��ڟ   2�:��R	vf�j�*
z�#--M���Q]C�/��  �aA�ǣ@ @�$#����p(///�k����ҟ   2�:,���<�iq�+--M>�/�>�?�K ��갨�\.��K"*5�/==]n�;�u`���b�O  ��aQ	r��
)�����jrrRn�{��&''�!   )E�â������NA   ,Z��~�=`�w���Y��X��
��b��D��P�EirrRiii���LuS   ����7�����w���?��X��m$�ٚF��,v%j��P*vQG�W�΋�焯jܽ�(�!,��=lv��E�[���L���oþp�C�2��]j_%G�nD'e,%��&��-r�^P3�(��ΐ�~���4���cZ���{� l&r���Ƃ�~�踽�b�
���Cz��I�;�Y�2�eɿza,\�/�ŗ� �@ۙq� �~��;&udZ�t��:"�K�����n�0��,�?�����x��/����u2��u�_���Ů����,��?h{��X��v���Q-�`�K2�Z:��j����Қ��Y}��E���Ç��Ԅ۷o��1���ʙ�z������.ڛ�����8��gB�Nf�g_�_�y�,c:-Jn�:�ű���Q_�	Hh�� S�d25q���ں�k��L�ϬVVV��imll�b��4G���ʙ�zu�DU�?w�/!��2z �^'s{��S�1�����WǦ�����PZ��Z$v\~I��N����Oj"i6B*�*yo'糰r�^��_�k�o����Bu���y�4I��dV���+3������X��EI�:6�rn�m�İ t��<L�X<G*���e�Ւ�d����d2Y��8�;+w>�ٕ����P��ש��@"��<�H��WǦ���Z �U�s�#e2�ZY�Y���8��鬭e�A��Ζ�8���ʝO""�j� ySǢՎ�r~,$�}<���2�,��èK�D�h�Is���U�۷��~I��|���$""�&YƵ��c!��/�%���x�A����_��IH���U������|����<�̧����=""��TF�:��cqY�|�<�wT�GI?��կx`�L&���|��Ge=�����|�t>��v� pr�β��Q�e�̈e���/�˩�1�#jp������e�iii	{��){�W<�|�t>����A���c�,��~I5A�$��P�VWW1==�g�y�t���.�H������/�z<�s�T4�fao���œ눛��<=��ن�_���{��|�'��}������� G��� 89��cO�  x.mm`:}ng\���h���'�կ{���:^ṕ�7�r��u���W�cj�����ف��_B|-�_\�������9������?r���7��Kptv�s�-�#s[����q�?�v�^Ͽ��焫�K�Z��M&n�<u�#��R��ւ$��K�/-J�=�8Z�c��QM��V��������6|uiccKKK���X]]-�y8�YXYY���|E�Y�o��#��@;:;��4k%�{�����\���y\җ��w����7�:}����������7��<�^��$wv��:  <{��mq\�]����9z��7կ��=�n�w���I�u�f�/>���|/����aDc	�[���-�,N�xsW��v�d���x����W����z�����\���Ww�#��� w�͒?�*�ukFF���K�:6�~�b��s���j�,�쀩�{��arr�����/���}��������|fi5��8:;��߮��;ث~R�5����]�(����w5�I�_K!89O�S�R�G���l�;��0p�&����V) `j~!{��G��;؋xr���G�_wtv�7�Z���:�[��(�����$��������]=��ȅ�#��QJy��d���ϏB[ө�x_[MZKQ��֊,c��w��D�I!�N�ʕ+��d2<x� ���wiT��jm��ZΧ�n�Fpr���7@T��k)����-����!����a���M���ݥ���~���A|-��{GIDɼr+j����|�X��7���U�>'³w�u�f[Y]{Ky�+�'gv\�,-ͭL�F��[+�(��l�JM4�� ࣏>���߰��!�"���I���裏��{�5l���|U�����^�g� �ހۛmE���g�l��M�/l�u;{05��pdnK��݅����b::;�Pc�9y����jUMY������E�Z����lC��mDc���BJ}�k]iε��M[5���TSA�:��������7�7�,��`qq�dR�$d}}?��Op��Q�g��_@pr���C!O�n��$ `oi*�9ów�*���)7��X��.�#sp;{v�KUh�f~����S���yy��L� ��f)	X�����u�N��o���5��K�b����Nv��A���BU��_����������uki5m�嗒(�E��u��3�������D"����w��d2��S5��9�����D���|j;�;��4!pr ��H�^%1+�r�U��H���7���F)��I�J���CM�����Dpr�`���F)J�{����եQi#���MG89�Vn�#sN��7<��q
een2�u[��۟K����L��N<u��%��zݴ]c����ӨKت-�N�ҥKX\\l�����
���055���/Χ�{颱��u��=�})���%�?+�U��(��q{�S/��ei��d�ꏲG�X�����rM�1�����-I���N醩�2��Z*۔�ن�<?�Gm���K������J[.�<�xr]�v�sn.��V�s�����J}�Gc	��b�[k�V�tR"Qݥ\�J�.���X,����A,3z8������O?��������|�'p�fիc��&8:;ؐ��'gԆ��	僃��������V�$N�����Z
���E��q�G�mk;O�S*j�+׷��
�:���E��|�':}b[�47�*�� ����RI+t]9˗�zݴ�:�	�R�0�p8���Y�����O>1z8��x<�믿��9j
�'Q��_��M�N�@���-gw���|M15��=�+����=Ww���J+��BG�7ԏ�t������a�Ȍ|���N����Y����t)	���+{v�G�($=}�]�J}����.1����䌚�z����n[Z��^�6�ba��AJ�2�#�mdY�ݻw��3�`qqKKKFIs.�}}}�Z��/̝�D"Q��jΧs�؞(�P���\  BIDAT�)���\z+[�x�Y�#_82���;7;��t�������#�N
5J�M�	��	��4��f*JI�vJL�%������<�_��]R�YS:izLh:�����;>�����^���|C�p9��1�끫7�<����׭�R���.��:u��!��j�j�8�r� @Ū6�H��X[[C[[[��666 I��կ���s����E��{wnWl�o����G^��ֆ��&���u��9���Kx����o�vyy�}�[XO����p>����
�����+�������������/!�+��b�`o���+�!Kd�[��|�'���qQm�����Q���P��w��_��V���,����hH���hii�7��M������0zH{�'��/����ʾ�\���ػw/�S'�f[v�[K���t�;jz����� "�mб��g��X�� �U��>��/�����X���Ckk+�}�Y�ٳ���T�'����Eww7~�ӟ��+�q>kH|-���f4��c������Sy%"jD�\z"�#o�`��L�	�9ܻw���>[�&3% �������B��7��>rP�6:5��{#b��߷��;RǢF���̸W J>��I���j��ޝ�����~�ݻ�������n��	s�\�����'�|�4	Ƚ{����Y�����i��ԛ��R��WΦS����g�N����v|���|�'tI���ID�a���JkP���q� ��rʤ�L�V*u+++��ں����yҠ������hjj������֭[�����\���nA�$�A���E,þ}�jv>�|���z��&�`Z����o����y�Spr��j�o �'������59H������}�`��{N�@��'{.���\zK�$ˈ�Dd.����[�n��T� &udb{��a�Z__������o���|��)��v��N����x���ҎVVV�L&100��,Q4�@<���g��r�O�WTEs;{�9�=�|�\1�ȱl��Ko!��B��	�G����F\�]�N�;Ҽپ}�Ͻ��V|��1�ȜD���s���cSՌ���G F�}<�:2-A I��àH��h4�'�|_��W��_��Tg���v�����~�3�/�$	w���|�(p��p���D4�P�y�7����BprF��g��?r��.�Ԁ��5t���ߏ����lI�k1&�� tX3b��n\�W#f˹q�(��J��I���je��ܽ{�(��v�Ν;����L&������׿�u|����/~a�X���ԇ����%s�{����;�״>>����%�k���*$v-��]VI���R���Licc��q7J�LX__/z]:���b�Ҩ�I�ڵ��bdd�H���UMF����tbqq����*��,���	�P6��;d\�����X����<G#��ڒ$���_K!�,��B��ē�L,��4�$v�s�^��b�;;�%1XiB0�#E���D#Hg2�WCWWW��'�����'�O>�sss�{��f1r555�駟�7��M<��Sx�����Q�8kkk��Tr>wo7�[ng����-�=}N ����b��U�D3t�6|��>�ݯ��H#������`/<}�-�5���ݲ�3x긚P&n����|ϥׁ�F�$"��Y%1�v����~XVW����7�����.�:2Q��5��$�i�^]�������������a�Z��"�U��455��p����~�iX,ܸq�n��h����q�=t�f�Z�900���fD"ܽ{�n�s��Gf�g�K�#��������	'g*��4D�S*e�/4ѽy��|C����9�Mb�Rj7N��1 ���.���b�<�݈�DT�C���3=A�W�|mgƽ� ���FC �F��2:t�m�Z�=�=A�N�M��/�� �J�����u��˶�6����������9Ċ������!<xP�f4� �w~�w��҂��%ܽ{���H&�XZZ����n��n��'�@WWzzz��ގ��ܾ}��_^^�.�����c_)x�Q���c��/����l���`�����a��=p���l%+pr���o��{�Ww���SO�f��ܫ&�J��WA�:<u��v�A�>'��?�������VFDD��2�ɐ���v���6:��k�xA�i��)X�#S1CB��<�;�{�H$tODdY����YEtuu���v� ��������b�ǿ������}�>��3]ǘ/�L"��m��!]$���OeNͧ�b���>|�>��ABWL��M�:GgGv��?e_�w��f�nU2{K��6�5�#sۖ*�A��Dc��؛mjsV	��A� �+~,��xM�� E%���D���nA@ �:.&ud
� `mm��a4����o�z26����ê!������qUc���C,..b5��M@�������AI���:�sS��Y	-����=�F82�m��lC���o���t@�b�v���Ec	u�`82��tD�`˾�z`D���jY�F>�c���<"2� �9A�s�q�77��*��dRG�cBg�ŧ~�O����֍5H��t&S�18���G��e?���~��}�6���#����@ =��.y���S��Ep>���n�[�89 [U�7���_�xo]n<GgGիb�+�|�yO߲����D��0����߈ʕ��e����VM�}?
��C"z$&ud�zI�������o=��-xʰ���_��aߖ�#��8���(V�W��많j�4��M�g!�X�����;5���bGg���������*B�x7��^Q�2K��7���@��k�臈�:2� �$���ՊL&����F����ެ��T1ng�#�Ԋc�A�z%t���-q�J��\U;���Tٿ�r�!��7�`oiR�\��S�LIGgG�^�Qg[*��Wy5�Y�L��,R��.�߉�1�.������S7�ă�3�7���s"x�8��?�M�n���FШ����\U;�����lSv刊\�X�n>����;ػm)s4�@pr�n^�"x�8<}N�g�����I���z�5��]��=��9�f���}�M������D��_|C���;7��*����	�8z�hL�j!�S4�LB��� D�c��fXͩڮ�&�LWw/Z�h��TZ���*�ĵ�x�����9���8�Z�J�����s�7< �� ³w����X��Q�2�ZO�#�\�~8Q଼hgG]$;��~�G�!�C`�Ɩ9v;{����K�#�gD!Z'�~��TϷ��"�{�������c6϶T��*�� x���:}���۾noi��ϩ���~���^�瑲�AY�`o�m���^1���`u�
�YH���F�n4�|O���A&n �S[�+7��Ύ���t(u4��c���j����_�6E��O�3{�����MGt��f\#*WFV���;eI�N�.��3�*,��=z�>�#�S:�j�;؋���}�u�x89�k�LIr<��R���7���^�c�ów�9�mń�ϩv�՛+?�����f&u�+�ł�����;GD�|�}��m#%		��<|C�e߈���[Yf���;���@��M�JN��Q�j�j��r�\,v���I�J�� �U�Bϭ����X�X�����v�Ճc��s14�.OL�4��� L�y\�������͹��_���S�!�֢���oX��k&L�Hs��$1�#"]){E
-G�7G�~#�v���P<�bdoڪ�߬q�H��L�]�]��>�z�S�u;���P�Z]Wx��w�S��$W��٥�:�+�/�SϑT~F(U�����ȏ�z�5�{ng|C���sh:���F��	&��z�;ث~ �,�MG�+66_�s3&uT1Q��(�2��4R�����r�����rtv pr����_���zc���ܛ&=؛m�A��.u9dprF�O����/�8�ju��FLGgǮޣ�R%�_���q�i����4�k)�.OTe�Bٓ:}b����t����^/��_|��
��]{�������h,ϥ��9�.�ԓ�G!��=puw��ݕ=Sts�|��[��}�m]�`�*�q^}�r[�֫F�A�$X,�AH��l�,�2$IB&���$.�� �J�����u�t��(b�?�����vS������>�]N�s`w)��6L��7�\�u���O�7<�h,���}⮴�w9 �7)1:�"prX���	RDc	]MSI빂��܎�
e?[�+�
=�*U�|��l��Ko�����<}N�g����U�yV�{T:�V��7w�`�_�QX�����2��٣V���H;��|�o�Om+Y���tz.��pd�����g;�uv�]��v�d+�U����N�����}Z��3"&��B3��ԃҡV�_֣��N�7��5?�^{��6ڛmp�oG���sh:�=Ba��g5��V&��z� �1�#"������P��ܮs�P�JwKe����U��[pr��5=.Wi6�׍��g/�S ��<e���/�Sa�� �����+��_���wt�˸�B^[:?�eRGDD5���;�޶?G��f���;؛Mb7�f�S����B|-���͓{�m�YO��3�:(���Q�J(dj~�>'��ܤ3�Q�I�R��=���O��~v�2n�Q:��/�����.O�庺T2�|$=T��?r��~� �h,��郒�j�`�[��N�S���g�s�<0Z��s�'�y��LUc���i�9�������Ҕݧ��Z��p�e�Z�k�܄`RGDD5J�\�$����W����-V��(�l7��	\�	���j�,����ϩ�M�!�@v��w�WӤ.K��YT^_4�@0�:���P?��՘�u�����S[�+���
θ�k��F�O� &uDDT������r�Զc�����vـ����-M[lG�%��^B]���+���[�##�#s������Mh�D24��x#bc�9�z��89�P?B��޻�˸�h�����J$�~Y�x���r|C�r@�w���c��!ttv`�� |��[����&s���e�o�_������j�é��TZ�m3"f���T��z\>���P�V���.O�t�q��J� &u�bRW�����(	�rV�B阨Wg7�X�l� ���%L�����|C��l��=�[��4�<@3P�*���qT�2n�)��L�t5??Q����F �22����+�eYF[[���ˤ��teo�e�gy]7j��r��;��٦&����S�SL�`����^�r��ۆ^�3.��j\-=*������?62<U��?��Ƥ���H�0.��z�J�&� �$""""�0�ƛq�lv���~IT3d�daRT���([\� ; �-�3h�DDDD��R:�I���2�ɐ���pq,^�Ұ�l�㎽�Gd� ��DDDD��R:�I�)�2�eɿza,\�cSǢ)   �vf�+��������L�LE�,��/�0���-_bt<�n�0��s�QG����O�����G_ȸ�˸��5J��3��w\����������x��AU�~�k_S�<�9u5��s�V�&���2��ɛ|ul��'*`��q�1( z<?Շ}ˋp����� �2���D�c���#�U������f��f�1��A�t�,�����u�$��x��饌�ƅ���*�r~,�rn�m��0;""""s�4����j���Ts+���ș4�)$�[�_�� d��XJBW��&���M1�#"""2-:�I��$�3���CF����2�H[$���|�WǦ���Z �U��DDDD��V	� Iݣ��E�~{�Y9?j?{�"���nH��t:���	��={�0.�2n����q�;��L�J�ؑ��2��\)-�ۭ���0�QdY�Ç)$�Ɋ�KE8�2�G���q��Fi�yf����5�:����O?�4�{��w[!^����R�k� .���3�>Al�8��A��bEKKKE�H�_�V�uW�D�q��Fi�yf����%=: `[F"�2~��85z�Ƃ2�0zT�_����ʸ�˸Տk�F�gƭ︕�+���B���c�4z T;��E��/P�e\ƭ��N�h�̸��\z&t@/�$2+H��7n/]��(�H"�ЮY,V,..buuuW�>���(�2.���m[��3��w�R��LꈪOF��!�J�:6�~�b�S���)���n?����q�v5�<3n}�ݭj$t �_U�,��G<��M"""�ZW��`RGTu�(��C>S&�DDDD5��	��������H3�N� &uDU��6_Ǔ�C"""�ZcDB0�#"""""҄	�����Z�p=�|�$����IQcRGTef��	����DDDD�;Lꈪ̔	� ��C """��X� Q�1Y�rn�%H�0zT[�v;���vumkk+�2.�(�Qm�����:�*��}g�=+��BF� ���5zT[Z[[q�ر��J����ʸ�˸�5J��3��w\3��K"���)������ڊ��8��V�'��˸�[y\�4�<3n}�5+&uD|�6:�0zmgƽ���v��_��r�2.�2n�q��h�̸��̸��� 6�L���u��vA�ŧ�!Bſ@6�@v��2.���(�6ό[�qk�:"��3ro]�U��JG�!�"�V+b��2.��X\�4�<3n}ǭL�$B��w'_��f�}g�=0Z͘T�dY�Ç�q�����q�;n-��:"	@�5#1:n�V̖s�.b�Z񈈈�H_L�&�k���j$v-��]VIs�%Q�`RGdJb�rnܥW�}g�=L興���`� jE��q��U��A�M�,��/�P������ͦ(�CG�����7��O����v�e\�58�Qm�����8?jH~Ťn���Q5�2�eɿz~,\���
���C�����
0*�c�K"<g�x����k2��r!\��汶�q�^��#���Q�cRGdb�����uX�c���k��0)*	��^'�� ��p� ٠Q�1�#�������G�f��DDDD��/w�ҽMDDDDDT�d׌�ͤ���i��@DDDDD&$`ʨ�L�J C="""""2��(��ͤ�˙LPF��������C�q-��+u5��X\��ݡ�DDDDDT�2��72>{啡��ũl�x"""""jd2pq�����1�RW����f�""""��&���L��sq,���ֶ��������Y��=��/+�v��|� ������d��$��αfR���q{���L�������|
 ,A
��=�|�����I
    IEND�B`�PK
     �a�[$7h�!  �!  /   images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     �a�[��RL  RL  /   images/f093df24-6efd-4d47-a863-17c5645b3aaa.png�PNG

   IHDR  �  �   ��ߊ   	pHYs  �  ��+  LIDATx���}�$w}��|����͌��F �%�!!�aa�`־[{msqwqq���ᇋ���%��?6�6�ݰ��q�F�= �H�f��a43�~�zȇ�}3�W��_gfUO�H��KQtUfVfV�П�=f� ��{:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:�s�������kk�V���L�8�?�t�n7��$�$	<��i�z���AN�i�i��F���Zi�$�,�iD��T�۵kW�̙3�{�7� �\ Ё�!O<�D�+�h���5^���|����˭���w,,,��t:���K{WWW���u._^]��eބz����J� ȼ,��,����Z���{*��4Ra�6MՒt��I�S_]���a�m�Z�;��δZ�����s��S�3�v�;��ҕ}������o��N��m�|��]��x�;vl��W_�������������������io�KZ�׵��}������M�q<��ل
�VE�0��N/T�H���*�*����Y�Ga�gY68��L^eYV�h5�2�K�12�H�EWm�B��Q�[m�k�Fs%j6&[�YU�?�љ?����{��z�[.]z�[޲t�7.z �:�8r�H�l��c�ĉ�ӧOO?~��O~�o_^Y~��ss�w��=*���z���FS�[�z>��5Tx�Bu6��S��4M�$�yi{��ċ��f]��,�T(��
h�rW�-����������q��f�Z]a����o��uUI��v�~��+�V���Ԏ3SSS�������|�e���ڵk媫�ZU��e�G���s_r�%Ӈ�>s�̾O��o�=7�����۝�>U�ާ"�
�iU�PAۜ���[�V���*�����a,��,��		ky�r������ײ�\��������A�/TǕGK=v���j�:����bgaa��N�<����#���q.lD�&'Z������������yU��x ��l���?�������C_{��gߵ����n�sy��=�6�VA8�~J(6U�;_�Q�����PGQ��E�`��:�=i4� 6�@�?�t���m��m�z������^�o}�(
������b�̓Ϡ�5�Ӧ:�i�����:��Ͳ���l}hv����>t��h��{��g>�'�x��^����n^���;�mt`T���x�{_}�ս����'��������+T��k��;�$��&n]�֥o]
VA��,�%_��,Yr�������S�\�W�{�s����\��[_L蒼�90���+���4�[�v{��|W��7u���S�N�w����|��C�NL������w����S��~�Z� �78?���+��r���_����N������ޔf�ժD{ M���nwR�0�B�T����[�SWk����z	N�z��/�f�jz�f��ܼx��1��/̋	��܇Y}o~V��'�
��^�򪵵���kk�;77�/~�ԓ/�����X��u��2���]5O�y`�t`�����z���_������F�X�ߢ�|F��Taˈ0i7�f�m���z�Ts���~����ҹ��,��c��(;O�t_�9�����T?�j�n���N���^;u��g�{���~r�e��3���/��s��K�/x �B�c�җ����矿�S��ԯ����ވ���`�����Hg1�6ץ�ͨ
d{�ӛ��|oY8s�����û���e����$���'h4�{�˫��޹����W^=��������ƭw�u�W�����Z:P�����#�\�������t�	�覉V�,KvJ8I��m�:��y�������
qs;���i�eǳ�S�O����P���:^o�l6��I}��MK�C=�K��V���u���Ͻ����w��?��}w���{�9]L��F�%~���������?�K�<w�z�*�_��z�h�u���l�mY/Ǩ�p�̼h0k�ڿ���j �R��ެ	0z�ʎ�����>��Y����>j�t��h���z��z�-O=����{���{����/?�����}�0�@�j~��߿�o��?�ĉ�l�������K�w��_�h'�ҥ�>&��;���eʪυ]-��a�{�WU�WU�ۡ^u�fo���S�ň��^�cǎ�EJ�YR㻓cKg�f�9��ޥ����sw}��c��ğ��]��{���~7U�@�����W|�3��#/��k���wOLM^��|�Ĥ��j�A�$���8S%I���2{��Ϫv���ef�\���|�qmf/��P/;�8���0��=��b)j�/ �"=�/M%��F��E��N�s��O>��#/~�S���_��}�9�d5 �x�=����>�����_����݈�k[3I�x���`����Lc�7gk���ǀ�u�xviVO(��/t���-{^��>�ݮ]�ٮ�B��u*�z�y�����w)??ʗ�w�/��+++�z�_-���?w̓=��S����#�<���q9�/�˗}����3�>���v��V�q�
?M�ي�q�E(�z�)Xu�7�f'0sv����v�1}\}��/*��5ǂ�G3�c.7��Mem����m�e�vU��rL=&_���ˋ�����)%x���q:�^_��C����ĉW�O�����{��
c�q�"�q����?×���}nv�WVWW��q�<�����Y=]�.	vs�7s�z�e�W���9/��7R�/6[j6�g����W��}��bng����f��;��ּ�Q��=�N睯�9si�{��mya�O~���}׻�=�"C�����~��o~�[���k��Ue߫͢W[�t�J�znt�K��T��z}�����������<���lg�7����ו���V�,�������z��C�z��ceuI��V���/��<�ē�--,|���z����i��踨�=ȿ��#���?~�_��;wO�.�01�,&!���PP�U�z̹��<|��^�u%c{����#�^_vsU%~�|ƭ��zǛ�q�J_z�?�ϯX��s�vv���a���џΤq��������\$t\4T��g�?x���s~~���.��1��u�Hov���X��?u��l۶{�[�S[�����Nj��QVk`�7�e?�F��^7�#w�+���韫���u�q���.� ѝ���N���'ON}�ۏ�x��O�ʯ�{�.:.����ny���s��ݣ�3l��n�
6���*s��\�;��}���BϜ �JU�{��ks٨��	����Û�}�sn;
zC?��+��F���?2�P^�D5*ԛ����_�x>|�����~��?��#�qQx�����_�׳�gߧB��#]J���~� �wB�S��R����Ӳ\�K����d>ь�[-�>===8=��,����e����\�fn���}�ەmSVCPVBץn���dN�Zv\�������Is��~��v;�G�~��(Z]]��_��f#\{衇>C�:\G��y���7������>�x�����`6��l㕐�	�bv8o0w���,�u2ۙ<$\�d(:d���������� ��X��voQu�Ӻ��mS�Uc嫶���1t����.ɗ��,����.�J��C~��,ߩ�G~�&9ҹQ]Pi|��c��g��?�я�p�m��x��t8�{�;2�ȣ_����'��
۫�T*qC��V%��σ¬6kkk޹s缅�O��� �0�a!��]�釐��s3�eKKyo�|?�عsg~ ���<ץz30�ڝ�@�O�:x�y��'�џK���yOOܢo�"�|ֶ(*�����f�KY���Z�������mc��|�~��z�����U�+Ȇ���8�|��f�7?�ʿ|��K�?��"�ᴗ^z��������47�^���ٳA...z���y����K�v�Z��b�)��տ�:^.�)��%���o����z�N_ }��:�ف�k�-YOJ��� }�!ǔ��iAj�I�ں�g���J}��/�=�mS׿`p�Q�=.I{^���X\X�����k�>�虻���8�@���z��>�͏--.ܪ��B�P2ȑ�����q	h]Bסm2��uۺYR�%�ݻwB\B]W�����ݛoc]U�z�Ym.� �	f��0��钫ty���ϩ/*����̟���ݸ����dW�^��uA���ߊ�Ԡ'�Y]]9��+/dzz��O<�ķn����a�#t8��ї�����W���<���os��I?��;�I�I��Ozf�Nm��b�lP2�a���幄��V����R����	󩩩A�Լ�Ъڣe��/����l^��;��9hf󶯯��z~�={�x���˃]�ؓ��7�啱;���5�d`~�QC��jR�־�*.ڊ�e��	�����+/�����~A�~�C��I�����t����A��]�jׁbvJ3Z��� 7�gס�K��St�Vw���PzzX�!N�Ζ��������GYxM�9}�t��NJ������x�S�n?��R��s��+򋎲��=���!N��l;�}�v��싀�k��Q�8�z~�س������E��U_�Z ��p�
�����z�Z���,E�CW���L���XC�a�K�z�����r==��&U�C�.�� ��m�,���/4�����R*?{�����/^����5��t/��t�^���	N_?/�_�����T7��f.6�9��W�o����N���?��w��p�'-,,�\[]��z�f)ۮz���r��s�����rI"�U��7v��Gs�y�.y��C?�hW��.ƴ�achJY=�L��9�'x�\���Mu���8\M��{�yEQ3?�_+B=�o�CW����'�/t�v��]�j�׮Z�nc�Z^���ř�ַ��Wu��������^Թ����	�@�ct8iu��CEь
�PW�={� ��p�:\�2K|�R��U�fș��*z��\�����z)K�\w�~�p�nfff0[��޼({�nz��m�t.�$�7���s3ü���8��m����Ͽq�|������9��������D�߷��8��!��$UBW��<-��[z��q,�W9� 0K�e�t؛��CQw��6h�ä��-���}̺[�jRe��W{gΜ����y��l�6;ەuJ� ��t����iB_����y�u`+��n/��nw����J��j�s/~ͨ�,-O�Ξhx�ct8�ш�8IݎlN�2|'�d�}f��d�Io/ᧇ�	�'���l�e����vG�:zr)�K�y=����f�KX��={v�a.%}}�2�0ѽ��q�湛������o�/g^�=�Y�^��#�/dt�}�K\]���"��43���fI[�e�f��:��U	���f�4s�Y���U�2�g�q�r\O.,�,�lV��;��Y�Z�F^�/���>Ϫ��^u~v��k/����C��Q���m�y�u�<��xȶ��EE;����pR+;�~,%3��&��U��f��y!`�Y���u�tU)\?��d�]@�*��6~���\J��g�ǰ�)�߶<T�7�F��g~'��MU����{�wQ�㜃0��e��v��O��!��$jq��HVW�7T�c̽���e�Q����,����Qð6S2�t'>�֡���ef�����3{������Qm�em�z�f�>~U��f�2\�o��;���tv�Mf��st8�՚H'[����biI׾�IY����X�l�����<ި�e&{;s�u�3ꐮ��^���P��U}��{ٶU�1/��k����}�}^{��w������\�$I693��'��C��ISSS�Ԏ�����g@3ǡ�{�m��s<vYռ9{�]��;���e����m�J�v�u�s����o�t?܉l�tm���e�e秷��g��¢�v �9���M ��[�^�Lϴ'&&hC�st8I&;kM�s�����Rm1C��N_�µ��m�q7��3n W��y[T;�˖��/�[��u��_v��6����� .����g~�����X����.0�9�['�&�i��p�'%I�޵�_�_���^���a���iY#V�$�Bc�hUU�e������jC���c�풪��*���l����ظ�TE�{�?�g�����?�V=mzQ�m���>�^��Ȩ0g����Q�
'��.�%o
|/f[�z��	���'�ɞy��C�u��p<������M��ћ��$���j�?�j/��ס6��/`���y��Ԭ�ׯ���OBf��2���J�)���m]M�ݴPwnum�v�z��T�G];��<Ɇߓ޳>P�����ȿu����U��)�ʢ��d��<�W;�C�T]2���S�ykT[���k������s�'2��
F�yY��f�����a�nc�ۖW���wC�W��٧����w-�^L�SL�#��$ԩr��t8I
�Y�������%�Y�-�&U���X�J7ãl�Qs�9���nm����U�Wu�{^���Iy-Cչ�Ǫۧ~nN_[�}U�A�yV_TX�z�������@WxrŶ~�x�!:����_��>=��k��z+����q���g�>�f��C[�w%���mlf�W�@�J�e�<N�Q�m���ܟ٩N/���/ۦ�V��}>�7__L�oP#w��o�in%��$զY3����!��$��S������LhI�h�ց�o!j�
7��U�8���˪�u-����6m�8C�6"��J���q��� /kv�{���ng����u�{݈����^�[�¶�V~����ɿ	�N"�᬴��[W�K���
�P�i�4ﰦ@��%������0z��xY��0�c��n�7Յv3��:���൫�͉g�Ϋ���47�g�*��j�������۟b��y�>կ������E	�P�p�'��܍�a������Ef~:����3��f�i�J�uA[V�����xu������vv�z�~�:����<e��2�C蒸<:�n1��?�P���7��U�zX���P�Ԏvz�kt8I"\�叿�a��:y`�v	�|L��L~��,������
�8�����J��n^������]|�����~���\n_��~�}xTi�|��1�7��n�7�c�w���F2U�oC79��mWe5�~������g�bŲ���j4���w���Akb}�8�O����.�u��q�:Dt�MJ�z���K[B@�u5�پ��Y�!�̇9�[Y;�8%ٺR��9���4�[w[U/�����h޼�������>��w�7A:��/~O��;��;>��a}���N�d�����~ճ�����e�����]�[^B]C�����PU˫�j�.[�v;yɴ�#{�W����|����1�k������|��#�9�P�Ό2C\>��k��zcJ����C:\��Ü�Y%��E���rC	t]�U�:�%�V�����t+c�ʫ�ū^۟�j���4��}��S6n���8��ì�/�Qѿ���%si;7����@���C���E:.
�R��,��0J��5$�ԨK�L��%�Z�Aojs�y����0+_?��<���ju��[�������i��W���Fn^T�5��9�}�u�G�8="A?�u�������|�߆�`����pVY�	��זu�wt>V�_2�!���{Wײ�,dz�w]�/cmϾ=�>O3��f]3�k~F�g]	�V�f��2e3╅�� ���F���n�9���n�~�}�߭}�;��_:JN��p�'坞2o�jU�]�+���W���ɫ��ޠD���g&ӓ���m�u�������m�e�1_Wu\նnԁ.I�M��f���߿n7g�z���?>�����@��Zkkk:�C��Ii�S*0������.�m�Y�t��f~'����R�������.a�2�{�W��y>v	�*����.�b��.���f�u�9��	}�c�����t�C�{��~nf�:��5��6g\(�ȇ(����p�����4�#U���p��5�r7C@T��%F=�Z�IwZBo�{fO4[���v�f���ߊ����2K�2�:�՝������x$I�Kݪ|;x^ƜD�j�y�3YY{�ݛ~��Y���F:���~��Y�s�=a�u}�T��M//�����gC/�ׂ�C�y�%�}?Lӵ��� ��$�'����߷�fn���p��)�mn'��t 钻9�JB�<�ّKLN���?�ݬ�th�������6�j�n�s���!o���g3C�^&�1ü����d�3kE��Uu�2��a�{Y��L�s�@���4ieY���i���׺*W�r7�[��'.�׋��0+J��P�T��ץRU��<I��z��Jٶz}�o����M��N�E�nZ0{���2���u��"k��[V<��D����|�1Y��S�"�Q������ovP�n�y�k1�D؋;�烱�f�}��K}t'�4�{��D�K��� ���yu�_^ʵK���t ��<�,q�jV��cٝ�R���yT���0����(����}����z=J�p�W�R�U�Z>U%PaO(c�z�n.b>�x�^c�����뒲�6���uS����C�> ����U5�v�쳙�/���um��q�Σ�	��Ϊ�@/+��}�Y&]&�X�!��@�ҽ���.v�T��.+�;�t@���b�K���������1��Y��!a�zG���p{&6;l��(;O]��۵�>�}�dv�3_��,���J����U�-�=��N��9:����/���벟e��"Pҡe�D1�qs���m)���>N�.H�y����?"/���w�Ҽu���c���a��7����������]m_4r���o����`�b��>+>y�O�8�~O���lx��.A��J�9��R"b�!��$�G�5�Y�T��O�z{Y��A^�-�6��-E��}��*��Rh�[VV�.U�uwd�;�Y��������M��uh3?�]�7���)[Wv<�=e��?�$`:�C��I�4	�(����dNR��=���6_�w�
�����{������g�6�$-J��nYQ<5��Vv���.���l���wT�V>�9J��P��Ual��.on'/�^��=؍&����2�!��"U<�N����~T�p��R�Vj~����J˛=���j��_�166A���n�p���%|)�AB	�!��$?�>����߅����s�}���+EN�(W���K�1����jtH�n��}��g��>�n�8������n�F���*��]\�P��z΃=u9m�Hg�T%��T��s/k����x�)�PUPW�_UB�:����i��k���}p���"�ݮ��ن���7�T>���\]����i���M�i{�z����c�3�]����G�;�C��E��ݷxe���B�|.��/C�|��~~U�u�ƫ���v���q���[s�u!Qv,��K�x@�MB��9�I,�^XVB�S��r���}#J��÷t���w��������6N[��0���`]p���ZXu���2��9�Cw�oS�tS�c��@�s�G=?�FU��ެ�v{H�`��]J�U��s��Н��}WQ��W���K����I)��"A��9ǃ^7�0��q�B�E�ǥˍI�dh��*�+f/��U�ö����iQ�^�_B]B?��3#�_���Ƥg�c͘�ǁ�c�������1��1���]�
v���X����A�P���������� �3]P���O\Ŀj8'C_u0N	}��:��
����u7x}��Z�ý���8�����V;�](�j�����a���o��?j8'����GI��cYY�����o�{�{�cJ��Y�ު6����Z��n�X]���`�N�:5����ajz�?������t�z�ױ8�@����v��_���uPY"��K�v��3^�{�������ɬm�h��	��U������o!\[��z�����p��׵^�V�����B��>U�K])�.��Uӗ���j2��c��$����>G3Х��a�$�F��|���mD��9g�#I�ָ����*�:����wv����6m�ㄵ��F�kX?���r��V��k���@�St���iƽd��Ӆ��[��l�Wm�/ަ�\54���ٽ�G����gܡ�r��uҨo���7��E����,����笭�I7�5x�0�Lh��P�6��Y�-k/�0(s;��}���noW��jf�LBq��WO^c�RdoF�#����D�l�:^�tjf8��溺�+���ڙg����^ƓۡY�k�l6ϧ�4n.�:�����;ם��q�>{��ap����+AW�*�mk�6O��nfX�߅����۱c�>':��9:��X��S�ڡg�v]){T'����� �L/w=�NU�}PqS:��_�z�lWUU^������m�?�u$ц��pN���8��?�U�6��{t��i�MTF%FY;qq��������Bw��]E_��[{��"��f����o�Uϳk3��!��Ή:aЍ���?�ڕ���oD'������nU;��}{�%\3�SkJX���}�~���f�׾H��A0z��9���*w��@�sz�n�&is;Jav�U] lf_���9ŪP�K�fsU� ]�^W�m??���sd�����<?˸e�C��9i�Di�5���*󪒧ݩL/+���C�n�V�qIU����
�q��B�Po�;,k���EUII�@�st8g�kK�z�8�4\���3��:ם����1W��5��n��n�Y�����};.�~e;�cT�����?�Y^��7�Z����e���aT�E��lU�7����U��7s�� �ϣl�fj=Fu���g�}�+�8�@�sf���V����d�5�����}�=/��c�?��m�v�ږmƈ��+�#;����T���O{�Z�{������o&�떗u�+[6h���c�[=��r�;Y"?e��f���k�'�C��t8'��bU�j���ó���o���������U�U����~�����n�:�Q�s��_�!��V���ܟe�vR3��ڥ�J�S����ۮF.[VW5=�٠�������l�}+�c�_��?��3��9B��9�I��u�SI��U=�A�՗4�v�^��k�zU�\WB�k�Q�޶.��:�������7���x���"Ή�8���ۣ�8U�KWm7v�M��}�u�Q����*ԫj%�>S�g����ۼ1n绺����H�ڵ�D��I��F��NkV������ێvk��_]s�8��}�ǩ���of?e��>?K�*w��@���,���Sܸ8*,�J�췪��r�~ͺ��nf�-㢧,�G��@�L@�q��~��߄��QJ�[t8I�D���C���B5��6���Ԭ��=��<���,�WU����F����6e���/y�Fc��kp
�����2Ը��l���*.�b/[^V%=n)u����o�^�*����n~^}��S0���[�z����a����F~��_ϲhq�*w��@�s�N c�T���*Z��L�v������l�Q!汪�����j?�7�;�f#��j��ϒ$��yn!��5��*�Ū�+��Fݶv'8s����,VY5��>��ZW%^v>U��v�qFͫl3�ovgr���ߣ���=�%=&s�st8'��t���?��8ۏӛ�j��v7�6�q�n{�6��v�����R����#���ԍ��p�JqU ��0�GmkWKۏ����4��q�ᅮ]��g>�lS����U��EJ�R��oK�4�����d�B��9W�޽:15qxmumM��5j���k�>_ea^W`^P���ou�V�W���f1����gn��=/�v�e+�ι馛�����?������e�����Gm��*������mʪ�͠�S��߻��~]U_7�m��l{�d���ȗ���Z[����� ��p����W۝�[��^M)}hL���lhօhK���0{��\�u�����M�B��|��뎿*��G�z	��h~��z2����gfff�<�1:�tٮ�����#�p���w�?��j5�n����<�q'�?v�-��73��T��Z�=�7�G�/Қ`'4��Λ�� �y������7����=�n]v�`��1�i�u�m&7:W��$�~�aC�GJ窔6Vgg��������~���=�1:�t�~������g_�z���{��zؒ&��SYi��f�'۽��sU�P�)p�ޚ<ޮڋ�Ie�4Ο�o慏<VW���Ԕt�K���������;^� �p�}��w�|�S���O^����˓S������?�;v���y�ũK�{y��wY�v��I������7�����m��������D*u��_g���n���̮o�z�ۿu�o�� �p�/�rˋ�O���ǎ��_����TImJ�R�ڍ��voDǯQ�3��Q�������٪�����}�z��PFJ�kkk��q�;w�q��/��W=�Q:�v������o�8����G/i�&ޡ��7󹽷�ڽ.�֗yo
�<.��yq�=ݷJn#g��r��`PZׁ��z���k��������ʿp���s�=�����^;s溹��I�G�`��jlWzU��<،eoFI��M���+ǩ��w�Ʃa(:#�T���̶۝��-W}������Ep�����>���������������ٳ����ĵ��˓�ovu�8��īT�r��GU��xS�W�Wz�K�������BM�ə(j~��W~�����q洛�y:.���p�����?���}ciye�Q�����ne�U3�����6���d���u=˫�_(�a�z���J�����;Q���]w�����=�<�"@���[��['��կ��c�}����_�${�ӹLB�
�b\z1J�D�ݹb�|�]ֺz7N^2,��F�{���כT7\�r}~v�@��7��k)A����7�쒻���C~7B��(
��2�[�=�q��n��`5I��&���r�ͷ�����#�,y�E�@�E����x�G����^��w��?%I������]�Qnmm-���	O�}>i�,��V�Id�,�����e-�fV�޲s���X?^/z�f:���-�GQ��JF)�H~?r���8������}���=w|�w�w��cs�T\Tt\����_������o}�{�=r�����v�T�!��P���.��=�u&�\f�eUښ��}CU�gͼVtu�����6κ��{�{ǻ�h3�K�cd�|�rQeV�����f��n����G���������ɏ��������y�ņ@�E�c���C�=�կ>|����?�V�~��l^�J��%4$Lt[��iNBEJ������y>���a�.���1�{�֗����w�y��$%ty�woԔ����� 🙘�|��w��������P[��������7���������W�������*8ߪB��*�O��J���*g�br��"�Ǩ�.k��+a���^�u��H���di���DչI���0�^�{��ϥi�S�;��m������sױ_��_?�o���z�Ō@���~�ȑ�����w���[\Z��n�sK�f�T�L�%uy^�d��Y7�jU�������P�����|�9V����}�]xLOO{�v[�n͢(ZPT'���n�ᆿ�����w~�wN��/�����o�/>��O=��|���?�����+�Api�ј� ד��,1�+>��}��ᠴ{�W�j��U�^V�-�^�����>�3�a�k-꿀���l��=�|?xmyy��k��������w���w�~���= (q���ۋ����<������w�:�ꉏ�q|����U�H繡<��3�����T�U�7�>U�fvU�u�{�~�ھn�q��G���i�{�Pe/���Ν;Nu:�^rɾ��k���?���?|����m�:P�߾��<>�ٿ{��'���_<����[TZ]�f���f��y�{i�zaP�n��>���=(U�rG�~�m�*i��KӢ��ш�Ҹ>+����?SQ��s�g^q+S�N��@3�?��=��C�F�����W�)P�K�vA� dy�܏\:A�D���ey���8~ٯ,�l�!�+q���hM�1����~��}���v�:����{�[�1:0&�iN�8���=������Շ?��s�f�Z\�G��\јh4Z����u����U���B_��{��|+Řv�lz���ev�3o*�u�~��4K��������r��BBj$�嶢�,׭�r�Qצn��7�:����v�c􋋁�����I7���7ő�2J@>r���k���={��}��{���=w��ڭ��z���?� �F�����}F�8s�ȑg�|�k�}����г����*����v7/���4�li��-3�I��>��R�zg;݋�n���4袹<��;,*���x�sʗ�r
~�3)�����7�G߼����Q��:�C�Q^ji��?�u�@:�u�ͩ����w�ջ��n�~l���~�~���8x��O^<���:s��.�y�[f2~�%ռ�4�j	4	}�3�.��Z�r1�N����½h���ot)�+J�z��n���שg�lŪ��&]e��]���D��ЋuM�y�$�&��W����[[��:33;�e7�tӑ_����/����= �@���n[y�С�o�����s{Μ}�u䅣�s�Νm�'VVV��V&�W�w���L���T��z�*`76����w2��T�kK��7$��y(�IU�*�#뇻�%`����~����ӽA;�9�����p�`Pj/^��EI�η�.�'{I� ˒ �:�3�6�����PF	4���5�\�]y��ށ������=� ́�!Ёm�������ۿߕ��۳c���������z�T��?~z�ɓ�/=q����O�v��������4Nw�i�����P�9�v�R%[U�UڏT���O�f��G�)-�!L]��C������Л7o�?���j]"�(
cuы��'qG��Ν;v�^�������}/_y�UG���K/ݧR?���[�M��>��O}7����q����6�lEo����+3�����v�={��j�Zs�_��^�G�d���ɕ'�T��������������/_XX����z�Z�����M��ܭJ����۩WJ�SI�����L�%�U��ϲ�/�ȇz�^��uM��Ey��4oF��Fo���|ԩ
�D=�4M�Q���z�N'Q�Z�h�vL�\hM4�,X��5yz��'ffv�����������k��bi׮]k�\rI��K/����������굓����}2
�5�S�������:t����v��W�a��TS�n4�ׅRGm��F_�屡z�رc���-y���E���拇ʹ�xoG|�ӛYYY>���|e/�'	x?h�AI��
�@����@oPtf���m�;TRG����T��Ժ%��륙ڕ��˂�*���M�ԵZ7����;�v̪t����;'^qp���n�i��ɩ�����
�v�OA��k���.@�F���L�h0O�:�=j�[�/= ز={�D��7�^k7�(���lMD�}c�LZ��?aJ�)�����V�
U�?�Z��4I�ιsa�q��z=_]H�Q���Q��	Μ97���MLL�vRr�/���;��
�$�Չ�)��*\cu!��ϕ�߿?��>�ٶ�Uo�f����{���	?����A��= �@�(I��^��(���1�����wE�h�Zt|;�ӟXe�����.T�?�V-�ߩ���j�y?��� ������*j��ݯFN=n���R����=��4(�������F�[�q��ɲz�^�Cʔ5)�{ȥi��~�VAދ�f1$/-��z��تkU���~�����˄-~1����SN7Aڈ�D����y?
�v7�K7�� j���,�q��0�F�wa�C]޽��ĹO�УL"<���y��Q�֖�w����[��lQx*����*q�2���{�~�ÀL�d�Aa��mr�9��"Ё� Ё-���zdQ�rC�<���gb���b'�ߥ��P!f��]���ɳ�Y��*��X�kR/jE�P�$�{�,��W�y�OF�0�\��FV�ԛ� ��z($Ё- Ё-�^�~��L����N� �Nrmϧ�W_>K���i�"�,zU|o�>��:�ER��RUo��|�, �J�����H�~����@�HơY��i�M4�[��I櫜��O5r�
pp.My��;��b��Q�l�l��̀�����5t�m������U���-�2���s�`V���
)�[C�[t�7�?��sk�,���A���,�Gk&�R�C��<��;j�������^|��ٰ��O�$�t��=?hqz�e��>?�<Hӄ�ܽt�@��@��Ts�\;Z\���q�
�a�J°�!Wvm��8���G���D���y#Ёm�B���v;I/ɢP�m^/��v����������O�=M����K{ъ�B	��� �@�*Udjr]��b�$)��x�^ѹ���w��Ǳ�4ll�m�DI�dYҐ9�e4�]β(��������|�����>`�\`�t`DI$7b��3^��m���%�?!}��\�9ܳ�o��y�O��{i&��~��y�-!Ёm�l&I�(������qdy���_�a��*5�~C.p��jy~Kw�_	`+t`�i+Q��n~C�^QM�8T�P���_�O�>�-+�t�$\� l�l�D��T�í�(M�*f���k^�QpГ]W�K߸,���l�l�b4����/5����K[�GX��+	�T/�@ς �� �<�R>o�Z=I����8^���V��*:z�(�(SS�����jrW:�.Ͻ���թt*� �7���8��e]�4����͆J����ξ=D?+�o��]^��=?����p�t`̤3�Bv�����Q�o�*w��,����+����ߟ@�<��H��ďO���x ��lU��|�O{i�7����$ɲ����7��q����O�O0#U�A�)�/���H�[@��@�н�Sy���Aѱ]��7x�n�����l��m?ͦ�����m���7O{ ��@��ҥKq0לO�n,A.�^���*�w�T&�o߾αW^9ҋ��a�O�7��{Ǣ��`�:�E:�n�n�=:����^7�:����td[z3����w�=��N��x#�≉�j����T���믿~��%:��fk��~U%�b�׻���zk�n7˲�ZM;z_��y!���Lοx�љ�駯��Y����6��T'��̻\=�Q�K��u	{��o�Y��}����{ ��l����WT	�ө�uZ�
u/x�oL�������K�ی@��W\�z�ر�MƓO��3���r��Ox � Ёmt��Ai3?���@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�����%_x\�    IEND�B`�PK
     �a�[2)h�V
  V
  /   images/72f663bc-d85e-4d27-9085-2f4219a623d3.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��+  
IDATx��{pTg��}�n���	6$�b��+��_�Hg�qԡ��mi�S�L��R�h)"��2V*4>�S�MK���S^�-m�1P$aw�;��s�ݻ��������w��{�o�s���� a��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0���~�6ml۶:Ν���0-�up��AeU%��� K�>
��)S&Ík!�?��=�qg>p~��ضc+tuw�[G�O�x�%�U�(��!�Lo��L�S�߼v����,��X/���>�0L�0��RH[[l޼�m������K0i���L�lTU�����Ϝ=�w��n��$DU��欙�4]�PQ�c��kh����g�LUTV����,\|w>Lnjn��q���ǟ�ښZx�W����pE�������X��ul��<��+���SgZ�%|^FU��'��)//�g�u�Л��:�6xj��a��M�زe�	VB��	{�_��á������wE��w��B��8��CH���m��t����^�[��h�N�e�߫���]�X=����W���n�GY\`%��_߂,��`pt���^���,�.	2� ��{�D�V�:+LAy	,w\k����3b�M������?x���+!�550n��`K�kͦ�n��A*�#����c�EUWW���O?$�IԲ�2�u}PpEF�a�:6�6��d>���fBc��HOOgK˟���tvvB4�j:��� 1
!��2��
���>���n!��?NH��[��
9$/������`4�Iyy��JH"�Ŀ�����Ax�B�t�J�ES\�8���<B�|�!0��Hq ﯋]�@,.�
�0�a��Jd�x6��\��iT�=�5�s]�ؗ�5L����	u���.�2|����4.\���u�>��@~fU����	�
���[z�{�4QF�Fֹػ@(.��d�%����/ �H|��0�>�p]n�[,�(NK��4z��X��UʃA�(�$ܓ�6B(�+�\M�f5;c&���x.wuc�V�,�h�(G��HQ����"4jH��L�a�`���D�mۂh,\`#�p�(��X4T��mB*����8���kΠT�Jͦ��T����
/���TQKr�=��?�D��K��Κ�N.��H�{>�'��t1��[`�u鴅�~K\�b�W1�:�Ғ�=�j�
�MQų��	L%��6Bz�-/��A=���'���bL��������0h��ˎ���G���M(p���t�
vݘ�]Ǡ�i�f0`%CK5tF�v.��fY�{�EZ)YVq�M�>G�?��%�.�M��
,���E.�v(�s����$��Y��4��4��CE=�������;��:.�7�-]�ua�Wͥ+77Z@���K�#�U,˼�t�z�F�B���}�﬽U���2���
��B�N�s�4��8:��J/�FVo�<;�-�n#�=G~T�q ����M�t�����K�����_O�I'S8mUIH�;�(P���oF�����ׯ�)\.�G���k�\`#$�Aǂ�13-�k/�N�ϔD��_4��y�?�1�=�I
��?��e�Ce�6BLS������8\[S�ö�{��?8�q�*��[^�*�����Ϯ[���+V�r5�a���c��ѣGZw�ȳ�Tz=v�cr����4卐�R\ĳբ�A3/����?�ŋ���r���p���.�BlX�.Zw��h;s�Պ�ʿ`�� NM�Vj�X�����(�⬐���^C�ͲM��}�4M�3�,�|<�ױx�#�EaƜ9�i�F�+!�����e��ɓ����US6~��i/�nrߩ�g.uwE�c68�[���4T04��(�8�͠���Q<�qUMe��o�ؤj�WZ���;�	o���.�=�w����7��{�O������So��=x���k�n��j����N�c�]kg�e�EB����8�M��ب[n�����V�������7�k߀��m��{�¬Y��#,�xl޼��������c����>��eۮ��IwY��E��b�^�O)bi>����XCǿ���E#Q?�6?۹Cl\a-�� :&8�O7�e��a���ߥ��׬���+��oD�Qx�����|vl����H�T�CYwRrK0���O� �fu-����7��5njƲ첡,��T�A!��"�`/�jC��It`+����$.��`ِ�~���J��k�v|`d�S��ʧ<�LQ���k�Zj�{!i+�`,G]���~�C_�bO���>�C�� �/�"P��y0t5-����勗K^O�:��^��ѣ��{oa/��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0��}jS�R��    IEND�B`�PK
     �a�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     �a�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     �a�[�łk_k  _k                   cirkitFile.jsonPK 
     �a�[                        �k  jsons/PK 
     �a�[�'���  �               �k  jsons/user_defined.jsonPK 
     �a�[                        }�  images/PK 
     �a�[P��/ǽ  ǽ  /             ��  images/0b351edc-7875-4477-b820-546ce15be531.pngPK 
     �a�[$7h�!  �!  /             �@ images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.pngPK 
     �a�[��RL  RL  /             �b images/f093df24-6efd-4d47-a863-17c5645b3aaa.pngPK 
     �a�[2)h�V
  V
  /             �� images/72f663bc-d85e-4d27-9085-2f4219a623d3.pngPK 
     �a�[�c��f  �f  /             6� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     �a�[��EM  M  /             d! images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK    
 
   �4   