PK
     l`�[����s  �s     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0":["pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_4","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_0"],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0":["pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_5","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_1"],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_1":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_1":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_2":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_2":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_3":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_3":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_4":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_4":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_5":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_5":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_6":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_6":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_7":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_7":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_8":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_8":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_9":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_9":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_10":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_10":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_11":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_11":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_12":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_12":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_13":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_13":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_14":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_14":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_15":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_15":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_16":[],"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_16":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_0":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_1":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_2":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_3":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_4":["pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0"],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_5":["pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0"],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_6":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_7":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_8":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_9":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_10":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_11":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_12":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_13":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_14":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_15":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_16":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_17":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_18":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_19":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_20":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_21":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_22":["pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_2"],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_23":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_24":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_25":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_26":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_27":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_28":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_29":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_30":[],"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_31":[],"pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_0":["pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0"],"pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_1":["pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0"],"pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_2":["pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_22"]},"pin_to_color":{"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0":"#ff2600","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_1":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_1":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_2":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_2":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_3":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_3":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_4":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_4":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_5":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_5":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_6":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_6":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_7":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_7":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_8":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_8":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_9":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_9":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_10":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_10":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_11":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_11":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_12":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_12":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_13":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_13":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_14":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_14":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_15":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_15":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_16":"#000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_16":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_0":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_1":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_2":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_3":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_4":"#ff2600","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_5":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_6":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_7":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_8":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_9":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_10":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_11":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_12":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_13":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_14":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_15":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_16":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_17":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_18":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_19":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_20":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_21":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_22":"#ff6a00","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_23":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_24":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_25":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_26":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_27":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_28":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_29":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_30":"#000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_31":"#000000","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_0":"#ff2600","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_1":"#000000","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_2":"#ff6a00"},"pin_to_state":{"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_1":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_1":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_2":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_2":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_3":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_3":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_4":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_4":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_5":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_5":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_6":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_6":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_7":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_7":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_8":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_8":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_9":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_9":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_10":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_10":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_11":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_11":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_12":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_12":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_13":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_13":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_14":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_14":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_15":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_15":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_16":"neutral","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_16":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_0":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_1":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_2":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_3":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_4":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_5":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_6":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_7":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_8":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_9":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_10":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_11":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_12":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_13":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_14":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_15":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_16":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_17":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_18":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_19":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_20":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_21":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_22":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_23":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_24":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_25":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_26":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_27":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_28":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_29":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_30":"neutral","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_31":"neutral","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_0":"neutral","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_1":"neutral","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_2":"neutral"},"next_color_idx":3,"wires_placed_in_order":[["pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_4","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0"],["pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_5","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0"],["pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_1"],["pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_0"],["pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_22","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_2"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_4","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0"]]],[[],[["pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_5","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0"]]],[[],[["pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_1"]]],[[],[["pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_0"]]],[[],[["pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_22","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_2"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0":"0000000000000000","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0":"0000000000000001","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_1":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_1":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_2":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_2":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_3":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_3":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_4":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_4":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_5":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_5":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_6":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_6":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_7":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_7":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_8":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_8":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_9":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_9":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_10":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_10":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_11":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_11":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_12":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_12":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_13":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_13":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_14":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_14":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_15":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_15":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_16":"_","pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_16":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_0":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_1":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_2":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_3":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_4":"0000000000000000","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_5":"0000000000000001","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_6":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_7":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_8":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_9":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_10":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_11":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_12":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_13":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_14":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_15":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_16":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_17":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_18":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_19":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_20":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_21":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_22":"0000000000000002","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_23":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_24":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_25":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_26":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_27":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_28":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_29":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_30":"_","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_31":"_","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_0":"0000000000000000","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_1":"0000000000000001","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_2":"0000000000000002"},"component_id_to_pins":{"880c9da8-a61d-42e9-aa03-4974fa913200":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"d7de94c8-b632-4e7b-a804-76d3686565db":["0","1","2"],"1f741dbd-aee8-4a67-9184-a02a7dc435ac":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_4","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_0"],"0000000000000001":["pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0","pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_5","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_1"],"0000000000000002":["pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_22","pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_2"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2"},"all_breadboard_info_list":["1619011d-0a6a-4db5-a57f-2bf7743e6a5d_17_2_False_730_415_up"],"breadboard_info_list":["1619011d-0a6a-4db5-a57f-2bf7743e6a5d_17_2_False_730_415_up"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[1146.25,522.5],"typeId":"b269da49-8c00-4ebb-bd25-5859ea0c7cad","componentVersion":9,"instanceId":"880c9da8-a61d-42e9-aa03-4974fa913200","orientation":"up","circleData":[[1127.5,665],[1142.5,665],[1157.5,665],[1172.5,665],[1187.5,665],[1202.5,665],[1217.5,665],[1232.5,665],[1262.5,665],[1277.5,665],[1292.5,665],[1307.5,665],[1322.5,665],[1337.5,665],[1073.5,380],[1088.5,380],[1103.5,380],[1118.5,380],[1133.5,380],[1148.5,380],[1163.5,380],[1178.5,380],[1193.5,380],[1208.5,380],[1232.5,380],[1247.5,380],[1262.5,380],[1277.5,380],[1292.5,380],[1307.5,380],[1322.5,380],[1337.5,380]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"8121d10b-aa01-462f-b512-c9e041cef6e1\",\"explorerHtmlId\":\"2c90d537-8abb-4e31-b993-0d96a3bccf79\",\"nameHtmlId\":\"8e2b9390-2a11-4242-98d3-e0f1a5ca7114\",\"nameInputHtmlId\":\"50ed457d-9bf0-4af1-a9e0-b3f116633426\",\"explorerChildHtmlId\":\"613f2efc-f32a-4427-af03-caef438b8426\",\"explorerCarrotOpenHtmlId\":\"e0d5828d-06bf-405a-a113-396603ce2d99\",\"explorerCarrotClosedHtmlId\":\"ef1e73a3-7240-4f3b-b00f-16a7dfadca03\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"f9897fd1-c64c-4b16-a0dd-efb8fb0fedfa\",\"explorerHtmlId\":\"f9527990-72bd-4973-93b8-f8fa75c21baa\",\"nameHtmlId\":\"ed748e69-112c-4f9a-9480-e153aa26320a\",\"nameInputHtmlId\":\"7f7c1e70-5f81-4714-8e47-950db47e39e3\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"bdcc2d1e-960e-445b-b7e4-807a8561b6d4\",\"explorerHtmlId\":\"60fb520e-6d26-44a9-a033-bb24aa7b99b2\",\"nameHtmlId\":\"e7815527-5d5c-4661-9966-67d441576d35\",\"nameInputHtmlId\":\"8a87bec2-4c24-46cf-a58f-33bec0334e7e\",\"code\":\"\"},0,","codeLabelPosition":[1146.25,365],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[783.4530505,155.6357345],"typeId":"d41d5606-8708-4dc6-b0f7-7b5da01a1617","componentVersion":1,"instanceId":"d7de94c8-b632-4e7b-a804-76d3686565db","orientation":"up","circleData":[[782.5,290],[797.746633,289.9991315],[765.3475,290]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Servo Motor (SG90):\n  - Red (VCC) → 5V\n  - Brown (GND) → GND\n  - Orange (Signal) → Pin 9","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[978.2041015625,232],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"1f741dbd-aee8-4a67-9184-a02a7dc435ac","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-2.08142","left":"677.25000","width":"700.25000","height":"692.08142","x":"677.25000","y":"-2.08142"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0\",\"endPinId\":\"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_4\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0_0\",\"rawEndPinId\":\"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"692.5000000000_425.0000000000\\\",\\\"692.5000000000_417.5000000000\\\",\\\"625.0000000000_417.5000000000\\\",\\\"625.0000000000_702.5000000000\\\",\\\"1187.5000000000_702.5000000000\\\",\\\"1187.5000000000_665.0000000000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0\",\"endPinId\":\"pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_0_0_1\",\"rawEndPinId\":\"pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"707.5000000000_425.0000000000\\\",\\\"707.5000000000_380.0000000000\\\",\\\"782.5000000000_380.0000000000\\\",\\\"782.5000000000_290.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0\",\"endPinId\":\"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_5\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0_4\",\"rawEndPinId\":\"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"857.5000000000_425.0000000000\\\",\\\"872.5000000000_425.0000000000\\\",\\\"872.5000000000_342.5000000000\\\",\\\"1390.0000000000_342.5000000000\\\",\\\"1390.0000000000_702.5000000000\\\",\\\"1202.5000000000_702.5000000000\\\",\\\"1202.5000000000_665.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0\",\"endPinId\":\"pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_1619011d-0a6a-4db5-a57f-2bf7743e6a5d_1_0_3\",\"rawEndPinId\":\"pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_425.0000000000\\\",\\\"842.5000000000_380.0000000000\\\",\\\"797.7466330000_380.0000000000\\\",\\\"797.7466330000_289.9991315000\\\"]}\"}","{\"color\":\"#ff6a00\",\"startPinId\":\"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_22\",\"endPinId\":\"pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_2\",\"rawStartPinId\":\"pin-type-component_880c9da8-a61d-42e9-aa03-4974fa913200_22\",\"rawEndPinId\":\"pin-type-component_d7de94c8-b632-4e7b-a804-76d3686565db_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1193.5000000000_380.0000000000\\\",\\\"1193.5000000000_327.5000000000\\\",\\\"765.3475000000_327.5000000000\\\",\\\"765.3475000000_290.0000000000\\\"]}\"}"],"projectDescription":""}PK
     l`�[               jsons/PK
     l`�[�5zU       jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino UNO","category":["User Defined"],"userDefined":true,"id":"b269da49-8c00-4ebb-bd25-5859ea0c7cad","subtypeDescription":"","subtypePic":"e30496d1-6e1c-40fa-a66f-2add70ecdc94.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"a7fde0f7-2836-4f0c-aad0-66dcccec46ff.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":9,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"servo motor ","category":["User Defined"],"id":"d41d5606-8708-4dc6-b0f7-7b5da01a1617","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"b3e67e62-159a-497d-aba3-70fd70f56319.png","iconPic":"ab942d8a-eab6-45a7-8f5a-30ef729b6f10.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.29614","numDisplayRows":"19.69562","pins":[{"uniquePinIdString":"0","positionMil":"308.45333,89.01923","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"410.09755,89.02502","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"194.10333,89.01923","isAnchorPin":false,"label":"SIGNAL"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     l`�[               images/PK
     l`�[�R�W�  W�  /   images/e30496d1-6e1c-40fa-a66f-2add70ecdc94.png�PNG

   IHDR  u  v   ��:   	pHYs  �  ��+  �	IDATx��	�ם�����w�}!��l��Zhz��@?aK3�`l���-Ü1���vws�c�w������=��-,��lt��#��%K��� �ElE-Ԟ9�ݪ�����̈��ܾ�9A%��q#n�ȼ_��"!�fs]uD��$�\B�0$R+�B!��� &�t���4H�BQ�&�뿿6�m��#�B!$71��_�yd�䪰��s˚�u5��NC��-�B!���&��E��]S($7	!�B!$/�UaGQ� �7玕�%�7��t����˒i�(���F��C��B!�B��EaGQ��u[7a�����������!y�ђiF�����!�B!�&ׄE��l��emM��8If��?�J���2)K��̙3�ih�kB!�B�p䒰��s@u$��X^e�������r!�B!�&W�E�A� yD!�B!Ğ\vu`�KB!�B
�lvu)R���B!�B)H�Y�Q�R �b�4I(z4����±ȼP(6Mb���hB!���d������gL�ۧ���ή��^7n�DB}���'�;"��|���)*�Hqq��_����}�Cr%�$���';e��a6m�/J�l�V�,7D�Z�Kk�B!��Ad����������'��s/^��󘢢"Yq�d���������_:}2�D�\_(����uMN?۵u��.�-��-��77�B�w�B!��6aGQGH����6�>�-^���u��f�Κ"%�ֈ�,����3�z�����v�.��]�X���vٮ���@6	;�:B�XL��D�~w�>Ow�u]s��ڪG67�%�h|y9��1���2���ns����,��v�.�e�fڪG�G��)�R�zA��pϰ��S��]��o���ϧ��lvu��8t-}х�İqsi���u;+ݼ�(nr#�!�B�lvu��0qA��?A���B!d(�vu��(���˥�:+vU�ln�H�gB!�B�@�2�6E!9JT|��K�b�<�uk:�S����̮(U���]��v�n�+�Ѩ���z��P($�)��a�l���n.@QG�����S���������:P^^������%_n�leڞX�3S��F7��ܺa����tww�},��%2r���8d�l��]/���������%W�^M{_�pXƎ���e�l���n.@QG���z�����ܬD��Ç���9������v�T��0A*jj���Zjkk��#���m��l]�[�ym(~����EZZ�?&ҙ�ab6v�X�%����]��v����D"ERQQ�քTODQw5��(�e�l7�vs�� ����Ւ
��w�Tg��@̝?^.�=+'�~[�����bn�!�ʌ�!��%1��?�=��5^�?�W�1y�x]>n�T]3C��~���4IF��D^&�(��yw����\����Q$<�ǁ:v5�lݒNҔt&hzb�/xL��.�e�l��v�"�	�y"�v�.���l&�Άx�\B̝<|X>nj��C��Q#��j���s����i@��a)���R,��v� o��5)�6M�/�s�6w��3&���Hn�h(�(�C��Y����<1c�l��ݠ��
7R/&�l����t �Έ�n��s{�Jǁ�2�s��e�q�t:��]�q�`�.�H穓����rd�T��?�/2�����^�3���J$K�G���D��>Jy�Oz�'3��v�.����^�p!���k��Γ�(�e�l7?�O~�qŕ+W佷ޒ#��i55Rk��+��K�"�G�ʸ��"i;}J�ܺE.�志ًɄ	�8 &M�E �f�#[�xQ���=�'m^�M�]��v�n����J����a�l���uDA���.W^��\?�^�;&}==��qWq�ʱ�~"��2e�!�a�I/a�͐�#�B!$#P�%�~�{�D��'�*�����(~ �$Y_V&�엽O=%���i�K�h8�$Y�f���B!$cP�8����C`���ʩS��[Ɉ�"�|��4��?ɟ��*��B!����Y.�񆴿�[�PV*�t-�.��7������+�ň$��7��/a=K��B!�d��Y.O��_�5u�r���(nP®�Hξ���;�]'�.^���B!�BR���@���;;��Z���C�
���YR"o�h�L�9S&N�*Ğ�"��.ٕ3/�pB!���AQW����_K�'�'��Ύ����G�R��.����e��մ�B!��"uHgg�m�\S[#�?�P��;�,���W_�O�/�q�&	���e��θt�B!�d������Rc���u��Rˈ����K�2��P!Y(�B!$cP��?u�|~�ti��J���Q5���"= hj��UUr��i�&`�+�D�Hӯ������L��,P�n��J��3fL���W�]��v�n����K�������]��E�fu2��J���P���}\\/;O������ ӥ�v���r���y�g��4!�ڪG6/o�޺��E�^�g���r�5�8�L{{�tu%@�v�.�e�^���\.X���gp�8��v�nf��F(�
���pD:._�l�(Vֺ�R�% SB*+D�AC�;�Ĭ�������6�4��v�.��8��c�:�\ii���vB�v�.�M��l�����x��T��I˙3���6�غO��!��BrO��Ӻ��;���^����t��vb����g\�.�e�l�i�^�v"�q;!e�l���n6CQW`t��H��2^�`8"�R�t�!�)���$��uk6ׅB�-n?�DdĈiM�4�b��b)�5�]��vٮ�v�"�,�iND5zB��ő�]��~�� E]��z�Ttg���7l�E�p]tw&c�j��ӱ�Iww�\�xѓ����]��v�h�+P����]��v�����("��^�v`�#��pcţ�^��}A�1i\�5��#���Yа]��v�n������]��v�:BrXʊ��f�Bٺ�9�6Q� 5�$�B!YE]�Q\��<LK]J�BrSM$������+����M�B!�B�%7f����ha�����\1�r	!�BH�AQW`�"ER\^.�L�:MuN����z��7�>�5�Y)��fs�@R�1tg&�T�p,�u�|��X�j��t`�l��]?h�%o���n��׋�]����+0FL�,��[q�X_�d#�XLjg��X�B����[����ۿ��)���:t!%覊ϼxe�d��v�.��/�z�]����f#uF̈́	r�w���L����b�!���O��;(��q�JL���}�3�x;5/�D��pmb�B!��E]�1a�l��g�IyMMV�:�>c�<w���I���"y*��&	E�FCrԼ]8�g��i��p����B!$7�����m���Ei�L^�{��U��kJ++���LF������6 �:�1�~�mB�C	<cQ�톼9 �Ƙ2Kgϐ9F�׻���!�BH�������jI���U����<o�Mz����/۬u=��9g���ds&���|Ff:���[�çdE�.�ґ��M����>-�&��i#���xE���D_?(�9x>�BH!BQW�\w���jӯ�v�Ȭutݱ�|�s�B����R���2�<�z�{fLTbo�S�$W�3�g�ßW�BN8��M���E�e��?S�B!�E]+��[�T"}�Uֺ�hTb�2��[��lc��k	���n����D�]r�52��F�_j�\ �®�!;��h�{v�.P�,��}�8�K�I�/��Vgg�kt�⵪���l�

����%K�x]F�-��@�A��Jw���BH62e�k�@�-���z�{��qawǌ��#D,q�"��Ϥ�CއuNY�6|Y�ϽV���wBH*`+���&�1���
� ���P�6[�*ʔ�0�	��xcz�O^�J˳>�-/�����KnW}��e�p�X�q�k������~5h}���Xi��l|�ׁ=PjZ�����X~�l|��� ���E���1�����u_f�3����(�
X����"���[R9r��_t^��+����z捴����,%]W��Gwi�|0sQ��6��(ǧޜ��%�W��^�p4�z�N�M���G�NT�~�0yHֶ��m��#)�]z��������k�'��k=Ld1�����'�j�j�O���H��bw�R��8�lu)Ʊ�_^?ŗɽ�O ��O��BM|�=����^-00&������t�w='ZLڡ�����n1���O��y|��ϸ/���>�p6�86W&~��@���-R�~��v����𙄢����t�����d����~Uz:;?�]�4]W8"��o�F��:���v�o�-�zE��ًmw䅣�o*�n���������u���B�_k�>��>�)�ښɤг��W���	��ǰ�a��ɒ�Ƹ�$�1�!��ˣ���6_�E�_YA,�Řઉ��>�q�jf���)�t��z��p]О��Ax��%���7=̖;e�B�|?yٓv��8�����x�u�/�PlZ��|�=��z|zu��f��M7��3����7c	�m���~�}�o,)�
�������o�������Gv}}�J�����/}�+a���Rv^�����RЙ���Ϟ��o��ՙ�x��#i��%z�ݐ�A���uB[i�� �u�fr�uz��, �yjV'c�z�����gF	��L�1m0�_Y��0��x鎨,9F��1��A�d��m��7�S��w�����ǈ�hA����B���ĸW���Ό���z}���8?�+������1lN��7�74������񷖢������kk�7��]�0i�\9y*0a��^����ZXi�	;��N��!�4��������M�T� ����g_2<tC
�̮ts���~���νmZ}� k!���D�ڮ~�~0�����X�(7[���t�u7��>��
��ۆ��n�����z��A�,fk�c|`���S�l�����_��,�;�/�+�)T���3��H���.�ʊ�"��%6���#2j�t�w_T	���������ꀅ�S_]-��Y|I���&���];a秠ӄ� +�<*s�ޗ�����Dx�Y�nH���VgGܽ�C�:e�o��,c⌶!�!Lp]1��>�߫k�����/�ԡ-sL�H��7Zܩ{��)����DL�7������G�[Q�^N�16�����\@�v1Np~]/|��G�Xt�N�PI_�v���9�c:p�xy��ݍƘ�k��J������Qň��kE?$Ľ�,ۖ�E}}���7(��n�?l����q;e�\�xї�)���t�E�/���~#-t>ⷰ�X�]P횅]�����?��>$O	
L�Ryr�I�����ܐ *%f��ۧvGN���ަ�_b���ya�:L�0q�rB�bhD�.�ؿ)_Z2H8@X��DN]+�
�Mu �cU�K��Ճ��X�u��	�����"���@�^�D?\~=��y@ kwD�}���xy�hGd�wf/���OQ�Ǹ�A�-��a��Ȭ�V{�Pԑ8�c�Ȣ��[�����+R?m���?�I���tG���Iф�x�7T{��m2a�A[�~]�� ۅ��-*����t�vOO�1��(k�%p�n���S�$;h
�IM�&A��K�i�x=�18`��dj�O.Ov�Ƥ�j��Ѽy_&&���t	
s������o.��N��^�� ��NFa��^6m���!~��g��D��8�y����>��I��'�;�vPI��3u�Eb��X�ZN<(��~Jjjk�j�h��N��h,&��R���J����	�t��!�ۓ�v+�.*���%�,(7@��p���+AYhnHzb��?0Q�F�vu�3��`"�[��,�WɅI�~=Â3���A��*�@z�D����&���_�gɚl���������	���w��_���Dj��$�"ᆸ�2�X��D.��=��9����ɍ���#�D&k��5%Yjo�5�y:���2i��㔂�쎘�:k׻�y�,�B
�� �{��}�8i�Ln�YW+������w�?.��|"��쑳o�!��=RZ^.��s��q=Ʊ����װʕ�+�fϑk?�X��e�HD�r�t�K��8���}pD޾|�>���rdu1�KL�G�:����x=�/D7$�~aԓc�V��l��˥�BH栨�������'��/")ӢN���y��+r��u��Yi�l�7WTT$+n�,��1VUU%����y+��g���d�	��KW���.9�Ijc6�v��,���fx�r��nHΞk��v��Ep�q>p9��h��=�p�U�.�[
��5�t�h?\�
�)��_I6�1g�h��ٕV�F,����������,�q2����:�f��m�GTIEE�||�^�@е�uH4���Z�(�ힱo�V��mF��Ew.��+���Kn�O;�a-,R�<~�]�`�D9x��,���\�e0��ص�����$;�|��6m�<����E!��1#�K������ܦ���H�(l�;8وj�V��n������2�&d*�?��]3�^|CV�5O��x�lX|�<���B����`\��w�,���������8Yy�Lyp�̂'��oճ/I!pǌI�/Ɠ�u]�`b��{���d��7��|����g��9���A�B���ۭ�����B��v�]� qn�Ə���L��g��>,���55�"�&����Sn��+WL=N �
a���)#j��X¢Y������T�>&�:B!y���a�T�L��g�������d�xϝ_�B'�t��fA�?����X�w<�$���[��:B)0�����<����i͸��g��up3��E�aJ}���z��#��{���8)�����վ��½u��I�u���JQG!�NL���7('T�s;2����	q��!$�8p���\aÀU%(��q�J���B�/`��=a��{_�s��:x�s7Ld����e�=w%�,`��G(�)p.\h�ʲ�5��L-m���nSK̻vۤ�|p��)˥��5/�5똝�J�������������l7V��o�ض�m!�b� �N\nl�[h�P����Ҋ_n��]6{��8[���<NNCQGH��'����G"��_���M���;���.�]p>9�*�	^���t�ty�ݏ���L�k��-�J���khX���E'�@E���g�(�qR(�k�vi�O7�U?~I��_1��.��HP�ȏ��H~}�tt'/��S�ejU�oA��G_> �p�X�I�?u�W�[%�X,�p�k�����O����n_��n$q�ӧ���{떑�v�G�{��A`��(~nqY(q@�SP`]̚�GOv�"�]��B'�~���.���e�/���3��.5ur�r�ZR�����b!��F�3�BD���	����3����v���ue��'!��������/b�T�������?�ӌ��N��iWM�{l{u��B1���R��Iv�/\+\�c�z����B'H�s���Źٹ?��+�cϿ��1������E!�d *X�t����)�����+��%���.7�p�l�_s{:���맨���8b`�we�1a����@d {��	������+�qR(�q�K7$�5?)!g���B2�v}��!������z�WE��K��@�!^.YLl�v�|!���ڤ*��Z�nj�6N
�|���u�P�BH�����
��Ec�K&�����VAa�6��a�öX�0%=��b�L������m��84\�$�������)))�p
	C���3�t�d-���\O������:gwV�"R�9
���2�&��{�-�T*�L�}����M!$(겔�HD"���]6��P(�����z締C��;��a&���pE����e�C�Tbě�dm���fApB�'(겔ʲR)-��������d�7i�<�ٛ��B��%����H��!vo�O^��Y/����!�;��:��U&8��"��(겔_:#��?����.I6p��]	LB�� ~A�,�5����q1�R*���z�3o:p����!�!҈�JG!�E]����u��6N�td�Ő� �5K�u�u��%IQ ���	qg�m������r�j�Q��R��[f����p�BH!AQG!��#v�jAǯ�
��t�<:���Æ�d%(�|۷��MQG!y	E!�d��[�Mi;���f����B����T̘('.�����(��<}�qu�������8S�BH�$%��^OV�ض��
<��{��];0��Dۄ����	�
�W{��vU=X�4_C(��L���	�GL�d̮U��X̟A�nX��y�`���i?����X�q;G���m�,38�T���"�F݀�����	�VӇǅ�6��!I������ yPV3h/ȶ	!�I&��CVg�}b|�Y��`���w6�uy���0n(��^�}�qȓ�i�dJOO�yd���¯�L>q5�}@�$V7�T�h�D���"� x �3N�}Z��$Fy��W��{�V���>��3�Y��2�6!��Ȕ�B���0�x�6����7�E]� +/n2u��ȸ����y��3�Aԩ�}	�^B��%e�3X��%�����G��.�����j)��	!�E&�~Ga�H�/��bN���|����Ж8�Y��MR� _��B��{?f�a��o�b���e�B�V2%�0�ł��{(��S	����)E]�I�6��z�UΘt��͈xB�3�?>�u#�OB�q2)�0'���]�Q�Z��U���k���u�ʠw��x�+�a��l>�M��u��;'n<q���..O%o�I��m��t�
���po�>�}ń(�Br�L�+�0�p�[���y!��E]��ڌ��p9�D)�9�?�3��e����n�n"�=k�b&| ���a�����U�"D�'��KdR\��Ƃ��AY7����i<ɘ�曰���C��/1�a)�ൖH5�h�Qt�X���g��F'3�%�c��
��`���	!��
��+/1']Q�7m~71n���@5�uyN<5�W���v��TQ����e7�Nɞ�O?����,��?�_n���Cr�\3���`�Vp�<�wu�Br�D�J�՜��q��06����:Y>z�P�9�Ϊ��-���������TC��cIC��N�n�tC�NS�����RQ�����}���M��*��p�'��BH��J��-fڃ�A���aP�--� ����R��ytd�?I�!VzEƗ�%�� ƍ�B��%��q�<��a�k'֍�U�@�;�S#���?qi��K����B!$U2i1üT%�3�=j�nr��3D�.��C���������@Ow׵�����	M��e�� �7���x��͙(�%�����,���칋�օBl�B!�ȴ�L�+ю����_�f>CQ��p����8�$&l��R�
J�J�.a鸎��!�BH�i��99�O3�:B!�BI�LY�̞d�J�e����:B!�B��m1�xӮ�?|!���c�^�����ˢ��E!΅mRY>8�㔉����*�W;�.!�B��L��`�����.�X �X���7|r�U:;:$bI���t�ty�ݏ�Ӈ���.!�R(d�b�6��vj�Os��|�������V���J,I�͵ӧ��ߟd����P`2kEե|��!$����5y��bҌڱe	1>o�Bm�<,$�&��,�zbng���I�Sk���c���=o�6����Xp�Ȥh�}>�����.�4o���z���.C7��m�r��s��H&�Le�b��2������#u�(��|f�ZZ��b�*�0߸�v%2�Ց�b�f=i��b!`Y+��Q��DYqL9J$�ʛ�O7�%��˄�2&���p ��b� �͢"m`тQogm��^��˷I��K�%��1�'�wӇ�n����7�������|���%��#�B� z��Č1	Od1�d��:�HC.��v"
� �����Tn��T�G_����a����)���1���1�zhf�����?���
s&����Uj�J���y���e���&+n�)e�E�7����E�3�q*V\��������	�ځ���{+_k�Q�B!�dL��.�=n!�COJMԭ�hݢ�_eU���@(b_N\��W����O��2-�v�?�D��?&�X�Qh�� u�z[��,� ��D.�A1��Fv��Wj�J���Dyp�Ly��)ٶg��>xX�_9��0�^�tve�Z�)T<�3�J�~���4u��!ݥR~5�:,}E�i���^J��$��x���%v1fLL!d�D[��(ڃ0H���#�c׮�f7MXӴ�(�����f�mq܉b����	�K��`a,Y���Q����P,rpfLTKKg���"�'���[����a�S>�c����}���93u��!�\$��h���@��*��#3nS��l��irz�ra�t���I8�h���5��w!��;���范N�qfں�8>�
��]
{��X̠��&�ɹ��iˡ�J*17`�3[⬨�+Kn�[q��LZ��P;06��٧��x�}��1c���k�,1D�t+��%��|���� �"(1��.�]�:@QGH����Ł,:�t�Vǧެ^w�T��7�O�;s���%����٦��ٲ�J��d(��I��]0X�Rbb�Nh���c��N��ר~���cj���""�1b=D���t��\���:+����Ձ?��)�� �~��[ԙ�w�E!y���*�j�NX!�(�!~2�,��d�.�~�}C�4`1�;��D�, � �pf7Ns{U�`��=s�%�S�K$ˀ���x�G(��s�X����'��vt�?��PI>�qS5�P� MW��AŨmzz��x]:����tK�uG���巆�7�s��S���[�^o�$S�dsL�S ��A�	�f��k�N�J�'���o fk������X�%�WZVv�'��.\M�~e\HH0��rLN�� �V2A�W��+?�!�OT"c�9\9��0�5i��-�4��3����D�Xt&�t�� .�IڡV�׃�Cܟ!�e�4.�Y1���w0����O��P(T�F�4S���y���|�d9�`%��z]"�O+h#��p��7&���,%]W��2\"K��6���������^I[�9i�BR�L� K�X*�	� FH%4�ǯ�׫Zl)�K��&J��\faf=�qX��ݢ3]ډ�e邔�� Z��x"p�2Q|B*B�Jz�*��N�X��awp�_!�d���}��)oߐ��I��$n�ü���}�#!���y��Úf�P�tnu�$�W��֤,��;W����ʄE���U���#�B!���$�ʹ!Obֲ��$w��#�B!���S�}@��J�W&PV:S�ARP�B!��@�k��X]eIa@QG!�B!9E!�8S�kdʈ!�B
���˕<+|NQG!̜	�e��{���D!��B����t�sy%�&N�x5g� *++�kkk�������B�Pv<����BHA1{�(y���dճ/I�@K!y��o=�
�Z��Qd��^Z��>���Mdl���Z�A�2c���`��/�ׇC6�-/�5h�(���梴���~����ˊ�v�RG!������_�|����D/�2s��	�a�u��z��^�����,kafʹ�m��P��r�O^V�v>�y����a�;��\�k��/��lqw<��1u�B
��Br��-�-R��,� DX]E�_���[��.��D�U�A��3 �O%}2>A��! ��@`BB�xj0�ԢB!��&u�`py�����Ġ��9�BDc��uS��s��B!dx(�)0�K�x�2���->�YӇ�Ӳ�Ab��2g`L!�BHr(�)0`�j����3?|A�l�D)���0�IR�hft��Y4ڶw�l%�Rq�$�B)t(�!I��S�S�E�o�Pg�T�Ol����*�bF��g�C�X��~�B!��:B
X�҉UӂLe¼�:ٸ��x"s��d���@�S%`I��G!�R�P�R`��HY��F�(��jZ}�e��.90h_�|��S�_?eP�:��B�]:�!�B)4(�)0��R�N.�o+�t;����z;�N|�*n@�ڃ��N8B!��ᡨ#��� C]8U����+�,n��A�i�I��-v(m��%�A ��9�PG)4��ר��S���s�$�r���B�N_����`��3g�hc�^O�33�c}����#B��#� �{�W�����!�l����ֺ��z8��O	D�Y*!!վL�a>N����<�d��k�h�3q�Ԕ�������!^�>)�Q�/_�p�}t��LQ��3dh?�tv��9tR	�|�#'<~�]��;��x��WdǛ��n�^6��g��;{ze���&?}�C5>w<�L�9��cϿ��ͺ~E�.��a�-3e���������^���������}j=xl������o�_o>�m��-���F�c�1c���gʉ˭������w4,S�֯xj�:v<8�~�g��Ot����r����\x���#��?,�[�z�\	�Br��U|o�z��l����<g��=i�Ng�L�T�[���v@,&+o@��S�Je������N�Pq��G$
��FGw�t��Ji�a	�'C}�=r{�a�W0y\}�<C��H*✀I*L�1��}�<cLn!dr�eF-��O���ƾ��0�Gm3DF>Z�0� v�k�!| � �c�!n��t���H��:-r ���t�s�{����o2����Ȃ�t�Ѷy=��zX�1V���m�1b�pXf��m+�c����C��1O��Ա����|�����_���*��G�|y���~*�qS��'�U�Ͼ�\m�q\xb|��1��u�B$��%]���nҵ3��"��$e*�$�ʙ��Jg�Y˛!�7�V���]��"���y�1!���K�k�&�Xc۞�s��R�������P�-ܬ�Z��*�cb�R�Q.�X �*֐��N�=�}�;�v�Nm{��59����q�և���hA��7���v�6g��ScWO��2�;�B�_�	(�!����vJ����HQ��yդ�k�L�6|�6�EJ"���o�~��l߳O�� Ŝ�'�R}ѝ+،vc���a�^�"j�,f�����x `;/�{DY~a	6�_�,^*\�l�X��} C�����"iuK��cv���p�4o�s�;���h4$�.�wʫ��&;|�YY���ߕu~@�O�;)!~BQG!9�.9�.`2z�;����j���>c镪�	R\Z+d(�
�Z�e.0	�t�]j�Mna��f� ��{,G\�0δ��������"��e�qiE�~�&�W�yQ}�f�8�M�|#�^�m����/�c��Y�#�N?X���B뵘�k� sL��c��b�������a�1AP�عUϾ�����S��Y��[�����/�ԭ|z��{�<���xL�'�W��?|AV�2k��D�b����;��*L��:B!�Ģ}���+�XL�Q'a�3�>4&5Q5�)�-䏮o^ły�v���L%w���+Y����d�!H��}���97O3D`œ��k��XQ	D��Ԑ�Xv�!T��J��uvV+�cL�^%bf������sJ�����������X�;(���ڕ�����(��P�B����Dj믑�1I)..��2���弜9sH����ȱ3%�H��bN"��@t��CJ�m��eɜ$#[��|���D��L�������E�hK�C��	I|'X�,�#�x��x���P�B��~�)�9d}U�h��>�_Ξ��L��))*�P�uwwK��I�9�_. �	��#j�4?����g�u.��̩�3�ϚIr�qL86�����H2,����鑋W����_ƷQ.��Zs6S-�N(�!��b�r��a9{r���t�!�
'�
�u��\Ǯj�m�7wL��7gd�50)��ʤ˪]vH$��u˴�$�����Y��FKQG����B�kƎ�A���������qR?+�.�4���s��</̍d(H����eu��{}�v@p_��ms���O�Bc��3Q�OBܒ����B|e��OI��c�u��T�^���1�tV�)�/�N��d_�㪷���X�襰��'�l�S�Hh�,��9C�j"��hn��Jة���e�p�5'@��Qܛ�p�EB}_�h���Ol��qW�,�$?��#����f��핎N���>ii�Pƌ����1a}�R�@D�>xDձzͦ`s"��i�;F�8��W�Ώ,�8�g�	1����b��uA����.z�
c|�S�c��2�Ȕo�@Hn7^Ǌ{Vr회k��AĹ�����B�k*++����~�\��WN{�vb+�}��E%׀0���aiy����3���c��u� ұ�+�0I�5ˋ�(~�ъ[f�b����*&�~Ʋ�Ya}�M�˼�d�b�E!��G�d┹r��>5�[J�륻�\Tu�@�/�\� `�I�M/�w��
��ҵ�Tf�ŷ�v=LG�y����>B6B,�|��܊;��ç|Y{m,�t��C��BP�m�b����k�6�	�/�K��c�I�:B!CGJ��l��!RT*�'�$��~(}�HQ$&�e��s��~�#��v���?��{�᳷)WQ7�v�l
b�
�b��7�d�n�������(����Y-�ee�neUی>I�X�5�`Q�*N�\c`��X,���p�������z��1�����B�@�8�!�p�9�N c��㇫0��z�m5&u�AB������B|�f�Jع��Q� �����6)��H(��r��8r+X0�D�[B7`��:f�n,Rv.�$I7)
&�8���M�2���Բ���dܫ�:�K�!�&�ւ֩ �c�^&��k�����9"�za�����0���N��� �-�)<�I5�	�@���k�W�߃v3HaCQG!y�ƥ�b��-�ʾ����/�����q��?�S]����hTB�L�+U��	�`����Y3�������25at
\)!x��X��8_XU~�A�B�ќo?�,�fW*���8K/ĉ���|N��s�}2k2=zU~V6X[q�ZHa4q�1�u���P�B�3�"t����¡6);s����$*�Cm��CG�����=+�b�ܸ]B��J�X��m��l��3��):#��K��v"75�o?h*M�)�Gp5u#��7^�:klU�V�L�sŽ��ӽ.���_��K�-�ΪJ
�:B�a���wjI��WE��UX�u����".O��e�-`1D���2�� ��jw�:Lt1��&ᢅ���+��"
�6���ǞE	o����+�a�M4�f�W;p�c4[1FP3.�v�n�R�g�x�JG�BQG!�XX���=&�?��L�:Q�a��붵�I&&�n,��(�48&XQ��I,چŷ�up��c`"����'R+��U�l�
. ���ڼ��eELtTɍK��Lpq@��q�
��Vu�l���y��B$}(�!�Ȏ�<��d]*@�!q�SWL=A����|tXG���qn��̻��Ä}ת/������l�3�*"�m{����J��v"�q�C���h�����b_XplڵY[�i��-j����5A�KQG!����q"\tz�\ ����%D��	���mpզW�Κ��چ1Z��\6�G�eV�Ź�춧
�ϟ��	k� �~�H��(�#��۩�����E�N����\;�.�*��z�i�CH�ˆ����E!�bb�C��N�e�t��ǉAܠ&�Y膋qD<�W�7T��o<���Ȅ	�O�V�+��o��6P�M�uy�dXE���ƣ{�i-�0n��ֺT��%La��$��B ���
[���uK	;��cN�ݖ����	�7ե��q$
v���r�� ����|g��S�~1t/�C$c�ML)������t�/�18�����S���⌱`���
�_�?-�(�!����t�b2�	0q��C;���,��aӋ�;u��:u ��*9
�]@w�3q��"��Y�L����1��W�b y�5q
\kO�Bk8w�h%��ͮJ2K���B�N�����l�v�
�򇉦������L�� ��V���N@,jk�)�x)]x�����uA~׮õ��F쵅.���+o����C�`[;�M����ݴ��,A	;�:B!d '�s$x�u�f���|����!LSu�QL���f�<%f
0
*�]�ᒉ>�+ӣ����A��ZE�3��RM��qg�bF�~���r� �E!�2�5{�p<��{�@�͙8ʳ�)�~�R����с	�q���d�Į�5�NHc��!��_������!�c����DU�.��|-5p�gG�w�vu�B��#Q�'�n�Ŝ��&�n-^&N���k�O�פrmR��9q^�Z�`�Lep�4�\�1�"��~�� �����������gm/�񡱳���"�㧰��#�BD	���M�[;ae�n�q7��gJT�9t�?���7{�?��87Ba�1�NU��i���%y�\-�r	��9�l�����3�{�Ə�uv ��J�r���cOu| �p��CY�<�K�Q�B!b��.�t~���L�MPHۭ%�0�K?�����H�X��:�Ŏ�������~Ԯ���~Ƨ��^�J]qxk��7�J�o�!�(�!�q6�Ǥ<�0ۻ~����z&�Dpp�1O�~欏Ȋ�WY���c��d�:?���͙�,f��9D.�,���uy����BqȕN�ie
�ab���@1���M'�Gkm2;V��n�]��k@������e�;l2_��hg��SH�_�L"C2����B!q`ep.�r��8����D�l����If^�[x%�(�!���ضBE��IA�)� ]��$��ɚ�U�:���	Ɔy���u1Ib�vu�BQ�:�^��{[����&b�PDz����"��lz�Kf�Ry�vhgIv���)��m:aE�.u�Ȓ��R��B"]aGQG!�8�67��0�|ͧzS�=(��a�m�>���Hn��5a���;h��5L�e4t�7���iRM�����1XDQ���KX�En��V}!����u~�U��=�N��]��\�6�#�(�!�q6�a̙��l��W���t�yX�|�)�e��L��}��a?k���).��p�3g�D�Gs.	�Ar<�CM����F�)�C8I���~�����*q@aW�vu�B�8���7wC�]�~���&��|o��M,�k�Ǆ�N5�섃X��j燨���c�G?���,jҭ]�(%D����ڸ_:)�ˤ9[&��p٥�/�;�:B!D��.t�~T> +�V)LFw<웋i�,�}��ʱā���u07k��	���_�m��֮�&�;|uw�<`�X����B qY��Qa�����s�
X��
���iҘ�)Ydq�%s�=w��Ch��hY���<�bj�X�b�L$�Y9� !�N�:��U��J�u�<�+?�����n�[�p/�f�˂ĉ���#�B������ŕ��k^΋:�+D��`R��=w���$���[f9�>մ�p���K �:^�Y½���&�i"��?�]�_ԁU�ڻ~E\ܤS�n��#��% ���K��6�O_p�\B�`D�"�x@}N��T�E!�2���f<��UWCX�y��/sU�BD����p:i�eԜ0���MYo��y���jy
�R��1�̶W���A׮s
��Y�q���@������3o���>�᳷Ƴ�"��	RH*��B@���?��a5X����k`b�{ս��`���G�DpA3'����%��;��	IV[#�J����������@H�p�m|ة��� ��&i��u�_WV�4��W�0k������v�C������6A�/�	;�:B!d <��S/�&��8�)� ��N�3pG��	��aB��J�ɂ"�oV�򖙆�IO�-�$�A�
E��Z�g����C����)p{5Ǫ�t3kj ��\��Z���f�$��]D
��E!�bt')��!W��zr���eF	�����mϥ�?��W��q"x���T��5՜��+^����[f�6Cȸ�7��;r&�,��j��s#v ���z_���n���
ƼS���E��<�$K�#����#�BL`��$f.%A�x7�.19�0��]�F��W��o �pP�@$8.�Hq?g�(%4�\���M���&c�f����\��u�E׮�L�v1vS�/k��X���ͩ�����5x�/_w�����{�1�>���N�Q�B!6����Y�@b��քl���L4a-YѸKe#t:��a��4q��x)3xx������F�i`��Z��o�FݷT���!�.Z���2��}��k���ƳٝSa��(!�L`�:7]�~��9)��XK�����j�xVaGQG!�X��w����L�1�#&�n3]��'�zB��21�,� |`�r
�t�d&��6' �k��i<�EV?�~q��e\K�?@��K����V��S1�kdWcd��h�@F�T3�&(0�����!!��XUl�����E�!DX�{ ���T��2gC�;���4��I�Y�Q�B!68����lv8�:X}��Lpa�q�7@;X\�ʊ�.�Ļ�
a�=M�lm��6�M`�k��*� B �ƣ�\!�!�>��p�*U��N4��w�\<qcm��ƥy)�����O�-�(�!�0�[9���lv�Y��v-��>��2���u�M�r%�V��Lgu+耛x)+�������	��$���c1��)�VAg�L�v�4[�܂qk%b���m]9��_nBR��BI D�]�M20��s�$e�ʄ�!�J:Y.SqC���q����D1e�g���K�A����:��"=?���7�U�}�����֮�p�����;�[�Z����:k0n����;�҉�n�:�k��̠�>��D�mY��Ld%�E!�� X'0�vc���l��Qj�dZr����(W���\� � F�Z��Fw��TeلE�1���4����������P��3�6�86�,�Nȸ9w�h[�O�1Ch�Z�eb�ly���K�Wh����$�,������J�*17`!�cJ��e�U��u�B�0@�����*�]1��ㄏ.U8���F%rp�.]�$A&�v�[���"�S�T�)��#X_��t[���y���Eg���jz����.���ע7�[�y����bH�[(�!��$�M���-3�q�'�^&	���uN�YтΩ`.1� ���ۦ���[&���nAp�x��3�?-f��t��BQG!�$!�T�f���dq��#���aW"e��*C^:V'�[A��J؁�b�w�V�]F?�}Щ��d�ѭ�e���B3p�����s�}\��7�N	]X�P� �l�@I܁q�4�3kL`�.�$?��#�"+���ݓ�(V.�TIsU�Ģ�!�V�*�J*�5
IkW�L��:p�C���H����O��(�.9�}�hA>Lܛ�I�Y\�b�"*]k��t�F�tNX�(�`�귞\�G 1b�C!E�bW��[`�k��g�^�@&��^ƒ��0Ǻ➻���\�t�A���t��#��F��[J�.I��Q7Nr������*��#fI���ɒF�TɌ�1R_\麝�!�||����Q�Q'9���Όj3$p����px%�4iX��
��(�84k/�=����5'/�w����fe���W�|��G����K�b���"�p����핮�^)�8�~%���_><u�߀����E)-�����M#MkHi�}'?��[���^^7Y6�~M��j�B�<쳮�Lm��;X��[��m�"Cȉ�$j���Z�(M?���e�vA㶦V*`�H��@y6��L�<���k��C  >�g�z/+K���V�v�V첏zJۇ��V��O�ȑ��F=k�:��Y�l?ky'$�B,&�KS,�i6��ɴP(<��	]
�M~E!��?|A��m�l\�@	���Nz��KKd��ý�'/�t�Ģ�r���?wD��kd�\�������-쐒<l0��uֆb���9�G?0�'�.qh_gI�˞�����x�r��N=;�=��5�F�!,��xS<����fi��� ���ZJ��%��C���iYx���R��d��C����3x��a���/��,��:�0��~���D[�Xט��l���DB��ZC�N��(�!$C�������N�x%�aB,���ݷHm��4�sƏ$�^��=9�P8"��r��n�T�ǬO�����˄)s]�ǿ��Aaw�;dGò�q���̠�`�>2ǆe;z�şqS�yX��/a��
d��x\�PBB�g�z�Y����k]� .��I~?T����j��6����Y�k���bL��=�I��f1�� ��h����v�m� ���E7�?���񇷮k6~����T��l���F��E!��l�Q��~ ��	���y^P5�Z)�?d���7H�كr���R?z�2:9
Yo2&n��9����̡����6��v~��������+�]�_�j*�>Ix��:�N�uՈ=�GK$Ա�ec�#N���������}Q�����f�9NJK�d��R\Z��1hA��)���C�Pr���p����'v��.MW8�"f�f�Xhc�_������o��5EJح���#��D9� �%�^ď�ȱ3�ܩr��o���D��HIi��D(���#k!&x�f�C\�zg���N'���9����\��:7����:	���~���Y��� 2p��%&�-�[C�!�c�Z*����Xo���z�p ����UŇ%Zo����_= �P�P�w���>��?K	W���0#�,�������9a���v�:\�s��M��?~a��W��񢓜��4��Ƶ��+�5�4����-��r������j	G���弜<���Ս��Q�����i:nO�_~e��]��z��EŔã%���XL��D�~w���խ뚍o�U�ln
K����L[US�BH��0_���#@��Ek��_��ܤy��vB�z��s2f\���a�G0&���������nX|[�-R�:m{u_�ʓ`ҌI2ĂrI3&�w:�^};�b�`��u���Ч8s?�2��Å�!n���Tv�\*��J��(��\Q-q| �М,�q,��q7t}�:�g�ƏG�Z��S�ں~�w�04'ځ�����h�$���87��קt��z���Ei�x.�*����HiQ��A_��W���uV��ij��ˈ1Cc��jF�����KW�>?y����������<�hDD�U�!� �y�a�߿wt-}х�ĺf���Y���E�pS���BrX>�Z��C��MU�4�D"���c�%%�3�� �J`Ʉ��dV�l���.}P[������eV��K˦_���3kL$��Y����eW���09�v�vq|�L[�2C����u=
��?5�(�	�ڰvM���>!��YJZ`=�����8f����Ht�:��,������];wXX�̥=r���>%��Vc�� %eu���%��J���:/nw 
� ��6=-~t[�tX�vu��� �%2����e%���'r��{2f�L)-���s.��&���z]�M��ܮ�G��}Њ��a����~<�O)A%�	
�DD��:�\&?{� ��c��Z*}����Gb�Dq|v�y��n��S�����U��Bf�=ރemH���ǃ�f���\�'��;���^���k*,}ϼ��%&F��^N��\m;穨õĒJVJ?x��7���w~<�D]W_ty�NaW��憈��vu����Ee���)� ���RZ1�vQ9s�}1j�T׌�&�*��ٗ������aV�@�`�	Q��������@�ud��y�$ی���I;��~�m�|rV�� 8ஸb�a�@[oͥ���J��5?����4h��cC�S�o�|cH�����C|���a�������hF�ˏ�O�O��i��8��c�z}N8fm13����Y*��"�������S�9(��~¨��<�o�z8��GyE��Ec���7��z�������9X�𛇤)^�aF%�еu�Q	�b�<�u���)u����	%�Y �t����}i�,���>Ǡ��.f[\Z/&�(gO�+-����q�IIi�tv�I_o����O�{�;�P�N !X���R��6�[�E�%�w,�ﺯtY�������/���1�|�d�8��+%��g���h^���&Xo�R_���eþ�YdC|Zף��P뿶���X�;�h���|���}��e��rN�DKK���뤭�tuu��+��	1)���~�QY��{q�b�3ǔ[K����=�n�d����ƚ�p�7L�:B�1�J��hA��a�L�aW��i�I�)9{� �?���Ĥ��Lm���Duo���t0��|��d
��q�h=D�]�����,���'�7����\���J���f���땓�ޖ1c%ma��^�O��N��*ɬo�r�zEW_�A2��uͱ��׆B᧜~���Br<�D�8��/�K
���?�}� �1�k����늴�����΁���W!�d7(y0i�͆���!����}g�Y��j�n�����y�����$va:6�R`�\�5�x�d�b�|&�.���]�#[�8��Q�BH�J��A�Y�d��(k�����3Ӡ�mEu����D RT*�+a!���\}�n���Ⅳ�且�����y-;U��lvMkHX|\ǉ�"� ��	�w�E%{h��uu��#�GOo5�����E3�v��B��/���4�όk(!�"5#o����?_^Q+�ܤ^_�xH�B�bє����&�ıX1ǉ��.l��x�D%�%􆣍��0E!��*e�R4�'�)�47A�-}R:bp����}�iU���"Ο�Z���޾��K�IiɈ���KH1~D!�xO8ҟ�S'�rC�!ގv\��{;������W1N*�[%U ��bib*Fn����.�4������e0R&&M�E��A�#[�8q���#�"_�����@!����<2^��¡6	������{]�]�>k�+cw�;Kef�j<;�`]s��k���@e���'%b1�'��fH�Ius�:B!�B򈯿|ɲ搐�D��&�2 4Cu�B!��D:��$%B���Vq�ِ��B4u�B)h��A-��t�*�: N�?��APZq;�����7��/a=K�Rݞ��B!$�h�u�O�!�xE!������ 0�wm�z	���m��zw?kmB�(q����뺯_HrT��E�%.�[^~K�;BH�PY$��%�2`���⠬+E!���+��$��M ܏^��jj��B�B�@QG!�� D���\u8vZ蜃~C��pi�	!����e��.�yN���#�B���X &�MkP�ސ�F�`��N�BH��T@BH:ٜ��BI���ar�DX0��K&�7���z�1�-�N\�F���_8P~S���y���:�E!�Y9�^�\����*i�*�X46d۪X�TI���B!i��	�c�U�u��]v[�t<�NTq�Lԩ��-R��6x��<�|�?�bжX���2-�}�D��|�D�R��`u���ie��:X"�Ȑ �*z�X?����^aB�VB"�U�l^���u;%(��F!�<t7����?\U"�G̒v	K~�F�TɌ�1R_\麝�!�||����Q�Q'Y�tH�a�v�?�g`�N��6�_��Ab�襖�k���w�L&,B}fp8_d}����j>?��ZQI�!$�	ǔ��
Qg���u�B����zۥ�r"1�®��V*J�=�w.�|��oӇ��a�J5a����2�-|m��ji��e{~a��c�����8&}�Zܚ+��gt_�<�4>�ϛE1!�d���S�f󴮭�f�8��on�����(�!�$'�������#RV^#c'��zWϼ!��.] `�3��Q�d	S v��Ѯ��7�����.��l-`~bv�8��� ���A3Ě>��%���f�����[r;E!$�)���$��uk6ׅB�-n>JQG!FOz�3��A:6
�[�����R�/]0d��P8"��r��n�T�����;}|�L�2��>{{Z%WЖ2;+�ov�.a�]�p�2� �jVЦ��m���ǂq�q��h���$��S���猯#�d+��ܝ�غ���F7V:@QG!Y&�:)��pC$������%C✴�&�n]Ոk��r���#F� }gʥ�K���ϘE�-�t���D��oZ}���k�������D�K��)�N[��p�i~㒢��̈́%�X���W��n_��BL�n���S�BH�0����DJ���D�v�3'��d[�@���;SΝ: ��V��K��~���VKQQ�J���k���H�0�3K&b��2M]EY�u���a�� ڍ�B� KYQ_�Q�l^([�5�&J��F�i@QG!Y,m���n�=�o�*�ރ��v�H�O��P("�&͓����sU�Z�ɘqU�%�I>��tN�g�GB�}B!��&nj	@�A�E�Mn�.5u���������b��=�o�j�I$����Hoo��DJ%_��Ji�V�T����%����K�ߖ1�u�l��X���H!f���}ts�_��p���.]A(�!$�Ѯ�p��r�gd+�q�DN�|Oƌ�)��5����t ��M%�p�L[gFתõ�u��@G��g�A'OA;*qO�̖�w��#��v��U�����'��*+�-k6�$EqCg���B����zx���Kx��02)e��%�Ҋ�2aRHN�x_F��&�5c%��צpis�:'�"��ە��>�(��|LUV7[�(�]wO�ډ6���LQG�5`E�b�k�o]��nl�޺�t���Ѕ���*BQG!Y&��7!6�Ƅ>�K�F�"ŵ2a�r����r���w���VJgG�tw�KG�e�]o��I52���޽�u�g��u�F�$ ^,RwH�)�%ږɲMHv��e��Ue'k���k��5�d+n��$Y��쌦*+��dU^'��b{[2�SQI3�K6%Q )RE��w�{�y�n6�@_��sN��S�>�o������v��t%@��_n��Bz����������ņP�3}O����oeQz�~�:m[�����p��4 H*mw�l����ϳ������ηӦ�MM;r�pW�a�#�@L�~�P�͚e�=��/���
j��*��knYk]�A;3zԎ}��M�6?7c�T�֭=;�j6�T�ۛ�7�W>��t�s���_�|~ۊBzl���O�*��a,������������i�80�ʫ��7_�$S�KYz{g�=�U��ڀ�2������6m˅�n�Z��q�����P 1����j����cbjɕ,} �֨��W�Tȋb�3�����2�5;=b�G�"*g�K��c��t�c�!�/�R��r�M�����3�v���3Xd�R��9���{ k�ͫ��G����v�s/�Q��1 �$.����v�]��j�'�P 1��AA�����2����{����w#w�(��uZ��y����}MXSs��F�g�֙Ry����
��z������n��_8S!����\�.u�
�? �vu cj$�\s��qK��5��2����q�W���*��ī�L|U�������ﱗ  A"�@���-5�MN=3>�ySKl_�˞��^w��0���vk[�9����옵57Ys.�Ukzn���3�n�bm��/����{�  @eu s
n~�O8pxq��V\jޗ.��0�����/�~a   �u �R�p�W��+)e�  H>B    $�    �P    	F�   �k޴iӖU�VE� Z[[������է��   ���:    H0B    $�    �P    	F�   �#�   @��     ��ޛ���eT ���徎[��Z�j��ի;g3Y����c�T}�Sٴ�6Fg�   �W���s�����z�W֯_����ı�U�����7    ���K    H0B��L��`G�}�   B��d�[m�k�   <�:    H0B    $�    �P    Q.;��u��~�����vz�Ł��   @b(�m<9hI���ӹo	,��    �Ԯ;>d��ٺ�졲nW��2��    Ԍt媧@��u    B׵�����{��6p��\sYɷ��@��u    B��w��Ĕ���?Y��?]���9�y�;B   ���?���~���\t���t���L��m|�ƲoK�+AKK��}�n    *Rn��5g�������r�5�<��/�ۋ߷q�   @��J������7t��w?��^�2    ��k[/��_eMM����Դ���q{湷,w�m���\����N���=j�<��B�+����a�    >2Y�3���eK����q�'��С���_�;?og�L���P��׏Y63oa"�   �;~|��o�tA��+��L&��)�P�?>d�ׯY��#�r�6B   �:���ǎ��|��K3��w��(7�@'�:    H0B   ���}�G���     �u    ��ɡI���;粖t�Z[[�-��H���s�mj	�\!�   �o�k�O�wy:�d]Е�)�����;�r��(7�+w���P    �R�-�$���c����l�K�����fs�Y׺�&B   �D;�����7;r4�r��x䰅�P    	F�   �#�   @��    ����]ikϜ�F�I7���+�-�   @,��pq��[������)нv�'m������    �V��j��    �Z�� ��    �^�����    $B�� ��    $�v��;hIu��P    Q֍��Փ#�TkΜ���:    �C��Ɠ��dg��޲��X=B   �D��@��u    b���T�#�   ��zt^��P    ��9�y�;B   �X���+u�<��֏��ڍeߖP    �֜�F�>>L�   �FC�   �h���B�~�U��T<�LMM�˯�g�{+��"�   H�L����m��e���G��i;t�e��(��   @����ö~C����Q��z�2�L�0�UT��
�   @����c�mn>s��+�r�"�   @��     �u    �`�:    u��ФM�̝sYK:c��-uY��    ԅ7ߵ�'�λ<�n��.���N���\�P    �R�-�$���c'���3�pU��u    ����K8j���Ѻ(��    �P    4{��zo���V���������d�   @(�~�N�'����OX��N�uǇ\����'� �   �����^��G�x��{?�.Wo���rN��J[{�5�L��F�_X�m	u    �s�e[z
q
y�.��]���sz�Źo��z�@���������nO�   P3�C�e_����@'�:    �V��.�@'�:    �Wo�.�@'�:    ����a;n����/u�8���)��tB�   �SW��Z%���S6�wВ��
,�	�   @�/�ޟ���oS�uc'����w~i�/�@`�G�   ��S#n/��]v�9�xrВL���Վ]|} �G�   �������ꮅ��!�   M��6���	�z��e���z���-�����+Υ��@�]�喪��   @(�]r����.�i�q�t�����l�(:��D�#�   E��?�kn��+�]w|�:��)�)�����N�niPρΫ6��    N{�uo�t�.�����w]�{�����i�{��W�>�y
v3���˾-�   @���J��y��PKm]���^���U��ǚ3C�H�Ǉ	u    ����׏�C�   ��)�]C0����)�g���۔�׶^h�o�ʚ��Ǜ��i{�����soYP�*��   @�|o�F���'��K�7����[�ߦ\��ٙ�Q۲��Z[Ϗ8��v��Q�f����-D�   8��i>���-��i�KͱSo���=z�����ö~C����Q��z�2�L�0�UT��
�   @(v}�	�3�P��
���_8����r�x��*���ǎ��|��K3WT�E�   ��6W��}�G.�:�:    �Q��6��(�s�4�N�/�KW��8JG�   
ma�M�5gN
C�.�1����U9��q�    �B�(��!�O<{�������1���){��̓C�6=3w�e-錵��X��*Wu    �a��[i]�վjq(f5��1��?1t���t�]tAW�pVT�z�:    ���2�ݯv�-��B]�6����e�+�d��؉a��6\EUn!B   ��OL�x��=�Ɓ7��pԼّ����-D�   8�4�n�P�B*�@��P    p~�V�\)��a����    N�ϕS�R���חB`5��42B   �P���nh��,����F�u�:��~xf�x��]�!�Z:3o�n�m������nK�   ���i����;o�7n]f�i�����-4��n�]�ɺv
t���oO�   �5�S�/�3'
t�̡��`Wm�B   ��P��d1�zvA:!�   \����K5p���0�ނ]P�Nu    �@���O�u��G�V�,�^�]��Nu    �a�Ŷ1X�6+�����;�T��rY�   @��G	��]��(�u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#ԡ*�O��G^6ki���dldU����   ��UI��ܻGlÆW�m3#�  ��P�3gθ�qv
t'O�4�p�   ��P�@�`���iq155e�N�2   ����������1   ���-����Ӂ�_{[��tz�   ����6������V�ܴi��ޓo   5B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�5���_e���N	�~���O��mz�k;3d  ԃ�-[mt�U��:4�������\`��~z� �����w �z0ٵŒ�P��06l��S��x   �"�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:4��-i�⥭��ߦ�������   Q#ԡ!��ͮ\���6�m3    u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P��0�1;8�	��F�L   �:4�S��Gf���#�   �:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P����)e���~��Ρ   �F�k�;8>k#��@���l���u�)�� CݦM�u   �B]�8xf���ա������   ���     �u    �`�:    H0B    $�    �P�Ě�����)�d2���d�W��T*e   @#!�!�����,�ͺ���͹�u���   �PuH$���@�)����X[[�   ��P�DҐ�r.   ����9tn���   @#!�!��(����9=s---���j   @#!�!��JGG��C�W�$�  ��X
v�.�rl:c���Tp�x�   �8 �   @�����q;u��Ess�uvv   P�u��ɓ'-n�w݆   �W�:T-��N�����v   P�u��l{��u]`]�.���fl�}�   ��P���n����{-�f   �O�:    H0B    $�    �P ��ؖ�6ٵ�  ��]�-Iu ���n��  @4u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u "u���?�j��Z�lr|���W߱7G��> h<�: �Z�����T��e��Ykon2��� ���     �u    �`�: ei��#G��d0�FO���>bsss��MNN��![31S��gfglv������X�>/~�)����N<�b���-��,^�������W}��S�vf����}� �x��Pw��w���ޠ�o~���-W�u��kÀz� r�/���)[7L��>d�����uZ0�^{��_�/'���P}ڤ����]�7��`J�3��5{��]} Ш�6��(��yPw�>i-��r�PO��T ���ٮ��zkoow��袋������>|������CCCv��	�Fww�vs1
"���U�V���DC�'  ���Cݢ�����3��9rĀzSm Q������mݺ�.��[�~��.�`���y�fggmffƅ�~<x�~��_�L�D�P�
z���� ��5D�kii�իW��U@�K��O~�~�7~�� �.?p^SS��]�v���7o��o���8���ةS���^������z���� ��T(Lz}  c��0���G��m����*i浸��[յa��f�-�И��o��� r�ڗ��%��C���J��
&�y�ץ�^���v�m�ٱc�\X�>�"�'  �.D�Sǭ�����!YRss6;9i-s��8;H�:�� 
����k��~���f��׍��K�N
%���'���_1�DD*��/��.dEY���/�b������v  D�!B��h.I����5kָOÑ,����u۸q�ǩq>::z�r���� �s����	s��%�Vٴi���SQQ )��A$���!�q�O  p��ujt��4Tjݺu�a�dч jH��4I��S�+5�h�������=DԋT��QHa��+�t���ۿm===���]�A�����W���Q�  �T� ��� ��G�Gv�w�@�!���\�e~��_�����+��f�>	v  ���Sj ��+�����2�q���Y��'O�^�k���y�%�#�P�;  j�P�� �}�v��?����I�ya�@��O�ľ��o-nĝ/� B}�  �%B��J w�y��ܹӭ��\�ri��B���z���/�2� B}�
� �� ��� �T~я��D�O�  Q ԅH��k�˹��Z��A>33��V:.��}�)�xa�` @Tu!v�;��K�m���J���_C{��뮳���߯� ���g��7���q���l}>���gϞ%�#� BЀJ	 ڣOa���'n��JD.��"������kK�A$���e~���?��l};v,��  �!�huk��72\�z�n�!�Z�p~~�������̙3v�7ح��jO=�Ԓ�)�=�βo������p� �  ���� ���O�n��7���w��7ߴ���߱�^zi��`Ah��ܼy��a�'  8��9���j�җ�T�D4gR�n��u�h�����K���_�> ��u 577�=����!��a���\5,R��������4b}j~]X�	  �F����o��۷�U=�����p�|�w�}��/�l} ���B��H���h_�z[�g����`����~Gջ444d���'�����>��`�  G�Q*�r�h�m.����s�aU?�2/#�%׶m��p�F�U�BN�<iw�uW !���> @q��)���<�b�I�Z[[]��sW��A��g?�ن�U�|����ȲK���> ��u����][[���k�mRhԍ7���A|Æ�����>���B�yVP�	  �G�C(ԛ711�z����d��$���>g---�Un#�.��N�8Q��P�gU�  `y�:�J�0���\��B^�a���f����:;;�رcv�m�������oO}����  +#ԡ&�&''�'��wG�7>4�Id7��Գt���馛*
!�繪�O  �2BjJ+�jHZ{{;[#���?�qzO�h��ߐ\�nccceݞ�<W��	  VF�C�)ȍ����իݰL���*��_~9�A���ڒ����%ߎ�\��S�`�[�  �4�:DF�1�"*Iok����>粗�o��Sc����!�R�h��+�����Q�竴> @iu����t];=���!K���.���K��U@�e�֭eݎ�\Z��	  JC�C��%�%х^ȼ�"�������,���  �!�!���Ӗ4�k�R�>hа�rP��UR�  �4�:Ć��iULŵ���|�Y�����Y\%�	  JC�C��`�>v��J��i?E���y`�<�zI��>���> @iu���MMM��Q6�������cY���  �(�;�ӧ��   ���f�繯�l:�|�l8��tֺS��6�ZO*e7��Xu�%��i��   q���e����_�v�u�kj�M���Rf���u�%K  @\(�ͧ2{��=P����3ۛ�i���r�.�'�pG�Cli^�u �ѿ��oڗn�΀ �N��]����K�޳��\G�?Ͼf��OJ:6k6�ͦ��=���A��z�v���hv�n��P��Ro���K������d&>���ˇ��o���^��9��V��7�x���P��UR���/��8�\��cU����>�����Ѩ�:bK���������e��5E_�k��N|c��>�}��s������7��t���Y�]�kZ4%�NǾ��Ԧʟ�;���[�Z�9sư4�k��r��,����W/ƨ�GaN��8�\G��t~*Ѝ�gz�����3�ܽ������Lz��`G�C��f�<�B3�7==]��N곸J�^��3���3���6�����M��\G\�t����7�^�����<��u@v��s�}��������nG}.����gjL,נ ��:�Fs��3;j�<�����6Y�{������!�I�r��	ۼy��W&'�·<p�@Y��>�Vi} Pk��N��=X�r5���}�*]<�P��S��*����������]x��o���q[�v����Keݎ�\Z��	 @-iۂ3��U��s�=���J�a���_��(�h�JB�+��B}��>�ֽ��z�����z�  �mz>��ط{8{_߮T*�p�7%�!���g�yƾ�P��3��~��n���O�W��U�sA��5��_��^?b��F P��Y�~�.i�����-���P4��'O��N�^{-�挎��ᾕ��Ҽ:��W��O  j!���[|�[�s�uH���GC�^x�����mnn����uvv�O�ӊnO}�����U�g\t�nsC1�����,#�������.y��^�]�}��s��]w��n+�ձ�Cs���y�}�C�.`�����/9��W����7]m�_�t�Ǽ�g�������=N�I�<��	C|���?�W�����λ^��^瞽���Z��v���%o���}��ӹ�O�n�ۭ�^Uʹ^x��K.X�L���'�]�,=Ϟk.[|.�>� h�K-Tb11����d҄:�z<���O�=����C��z��ۦpV)��,էzYM}����h5h�&9���^�2�0G��>�#�X�ԈU S��u�.�u
{���Fr�S����]c���j��q�k�z
t����K)<N���+�qc��x�y�����U.�K.��^�R�\ra1wN(�W�*�\�?�{C�;�����������_�^�<��dm�bD[tܿo��!��:$�B]SS���������SO�G?�ц����{ϭ���c��1�>�
�>�QC�	O�#5
{C����rz��^G5Luu-�֩q�Fna#S�X5�ըu�s`}w��5�������!�u��U#</�U��u����a�ნ�PJ=�K�:��
G
T{K8G|��,(����s]���u|�{�������?�=��\�9^��J����ō�f��.�pB 7L�?��m߾�aC����
j�o��4�����>��8���,��@԰�A�5J�xv��\#:���5t��o��P���hw=u�������{
���!��{������F��:��Jy�ѹ��T������[ι�WK=�bCKWR��J&���Q�L� �뗿��k|_w�u9�Q�h�����'�ܟ�S+a~��l�`t}�� ���z;Dp��z�
�\���?�R��+�=�Oe��}T���^��R����+�Z)������T�ܳe�#�uC�B��YN�+�\_�ia�f���"�!47�yuᚚ����뿶����j��`
]
!���r��Ͽ����o���L05X\/�Ĕ���G
����<�K_5�ESw�BC�ͽ\��+��a����\,u�_���{�D��`ņ�\԰��#����W˝����A��z�^a-@���_%��������T�a��^��:$F�0C���7�\�cǎ��ի]�l}.E_�;�F@>�*�]�5���䵜��`.�R��0�{���?S�<*}/��Q�B)~�}���'&c�=j��?7x�綐��/~8b!�G�78/���,�}��s��{b��K}h�ܪ��Y�y�|�:$��Ԇ�=��Cn��64D�VgԊ�~�i���p�ҩ񪆈�����_V������]_t�g�B:�PWw�9��ł�B���o��C�<݇�~5� �I�~�(�����z+_Ƙ�S������9���ߋ
���M�u����,�}��s]��yr^h��w��4۶q��
��L��ҥO�C"dzY3�N���~���.�s=ӰH�T�����|'�2���}�j��3�O�Y��q(��!
{'\p�}�o ~�\a�ׇ8?�-(n��>�zF�CS��<��{����o���r�l���m1p����Ntn�+<�6�z �R��{Ҋ�GW���BŞ7�G�C"�|��Z���/�l�z�c��������v(��y�'�\jh�p���r�����]�6�2���0�{����[e�Rz�s�@��o���Ph�[f�e:�ԳV���Gt[d,(�Gn�\�/��R��r=���=��7�x��n�VU�g��J,����z�b�S�k�n+�xB��g����v��׻/4���l۶�n��&knn}�`~}����e�]-�s�̅�rC�)֐J��]��g>rvq;��T#x��N��a�����Vl��R�p�մ^�7cY>�-L�������W��=`~%�b���=�Z�d��]de�����:��A��Be�|b�g��C��&R�S��:Ğz�OW{��1��G>bO>�d]���n���m����裏֤L_�����π�O�}�F5DԘ��c���QH�G�׿U�m����_��b��󸫄�I�W��`�J!;.d�PJ�큘w���JC6�r��r��W:��y���CQf�
[�}�R+k�BbO��h�	ԞBH{{�}�pAdvv֒n˖-��/~������d�W>�gkk+�����n��S�������\ H��Y����v�����͙toٷ1 �O--|�y����$���^��K\ �bޗ�^R�ɡpX����߽��}-^6T?=� Ј�Y�b�rz˽��F���zvq
 �gr��'BZ�+S�����F5�,�@�(@�rMλ�v�uO��=��Xw__�z˽���E���]j�߻��VOD���'>���	�"��[�e_|ql��s�ƍ��O=���q���X�ƽ��Wc��l�<-��a���G��޾�D(A+�2�G[S��"�_���+�J�䦄:�ZRz����;���-[��U�V��>�1{���ȑ�/@���cw�q�e2���8�P̵k�&�>{,���4�o���t�?�-�}��{r{2��~�o���
wn�gd	�V��w����Ҿ\Z������(@�䚝ۣ�[�ќ�SI/��[---,�CSSSv��	��[\O�+����Ԯ�.�o��W_mo���=���G�@`bb���F}�G�c
U��������Es���[�ma_1��-?�k��ƾ.c	�`(4��L�ڤya�������j����L �t�}=���|-�U�����ޞP��R/�z?z]�p�M�6�s�=���n��Vף������~x�������g�*]F��Q��ˆkX��zs|O��S�SO!�0�燺��%�wA:���{�O�)k�O��ξ۷{�ej�t&Wfu�%ͥ��.���v:�v~��2��)*�/M��뮳W_}�~�X�P��P���!s�s��
r^��'  ��J�MM��;��Lz��a�����g���5������.G�S��52�k�f��뮻���_��4��𡡁'O��|��jP��ѐ9�ysA��#�����E.*�6�^X8C�mǍ[�����Ш�4Գ��;�r	� ,����k(��\����@'�:Ďz*��hs��to���<x�:::�s����Y��)Z���k�uy_q�v��i������˙���t��o��g�J��Ri(���K�+ĉ������^5C45oם7�ysn���B
Q
z�c�r�������������=��
7|�ֆ�Q�	 ��ԋ��o�{�k�J���}]��T<�����@e]�ɤlUkk(C\F�x�7'��nsaGC�4G��@��^�_��_wD���>��[92,����z�5�\Mժ>����ի]��^�T
X��la��k��G=X�S ��_E����_��S�{�����O.D�Ebr�ٯƩ���R�/%�ߣ(@2�-���uܷo�|*�g�����?�]���-@�:Ć��Ԟo�;�����W��Ұ��f�n^�(�|�����v�����GV�_j�G���/mr��".��R�k��"r~��[����܇ͷ|f��jU����YAY��~�z{��W���{,��Jܐȼ��n�d�2}�}�G�-Z�zs���_�>�|��[~/�׿��u�.��Pņ�Qn2�V���GV<N�r��@mh��fK�,�~��L�ؼ�/u��65omjڑ���s��2��������+��ȻvIg�FFFB_eT��رc��W������W����y�fף��ﭷ޲�G���ZR@�ܶuw�w6�~Ӳ�FU��N�էz�4�qfff񶱨϶ա��`T�S���D���W���PV��^{>��Bd�P@?ɣ׵�zM��<��p�����f{8����Ke3)�?.�mږqݖ������q��S����5���[��.����̴k��z	8�t��o�iq�zP������ r�m%����e���LOQ�*��j9�M�N=cjt����]_�=?|r�gG�R�S�~ΠGa�R���zE�U��e���LK� z.����v�]���RB"G����+>�ֽ��5�N�BH�-�QK�]k쿽�s��|�O��읉�����1k7�\�QK]vm��\}��U[��P/�B��WM
�P��ڹu�婜Z���Q���ϸ�Q�79wC.s�_ϱ^�Q�\ũ�L����~�?�"B"U/�Ns�^��K*�J�%�쳿y�9�Gh����e�Ƈj���7r7�炀��X���9�[,��E��nS�\��:\=���.|�Q�\ť�LHh�U�s � h�:DBaNC�V�.)���ؚ�v���� C�R����q,�H=�@�a���F�蹪u�~S?S��T�z���:�\nOI��M��{T{[���,ן_���'�5���^˿hL�C���{����#�F�_�R�/saÅ���!U���蹪u�~���v�EE>�y�|���U8�Y�Q����>���^g�ޤ�ʿ?��ms����x$��+}H�r�3��C�׊�"�HB��E��n�΅�W�{��&�b뙨�P3������ ����O��x^�����M̱�E%�>����C�G<���yznK��(k�)��TY*[�}�a�FLX�*DUn=WQ�����ܗ�p��^y�� TaG�K�g�;{�x��:�s����"��Q�QL�!^�W8��-�p476��k�Ø��-�*��q��u}������[����.W���?��~��^ޏ��?�A�;���zE�CM�;�b@�����`4Z}��Cr&5��/����	�f�¥6����h�o��j�y5Pܢ(���k�}�3�1)Ć��e�Q�\E�[�yQ�CZ���X��X�7nue�įt6^<o�ӽ�_�p�[�=e>䨞}o���?�¨g=W����P���|���*pz��<��P�P)�i�z�; >�'����y=F>�(x�J�qmp�aFn��\�M��Ay=�E�U#��E)���qs������~��^�b������\����z��ʵaЇN�}�=��ĉ��> ���>�C�g��.Ե��~��-H4����|�P��)�i��0��"ņ �rטPO^�q5X��X�<�c&j��b�Y-ʍ"HG�]�7�WR/s��S�>ȅ߻�7M���6�p�@�>���d!�[������Hi��Fa���繑����U����;�T-������z,n���ߋz^��P����g�[�<9��0K��[�P�b���\j�q�O��	�c�a�]~�)z�~�q?R�*�O��*�P�v�Zͮe��R��z�%��7?�i�!�a.���O�]�y�����p�?����ͽo��^a���
�ş��{]&a���ɇ��^c?3L�����ܞ�C�5�U�ר�zF��z��k����)+��9���8 ��FB�m����U4&� �'��F�_|��SQ�l��A����Qܜ�\�8�����\X^���y.����De*$�h�����sɯX���lj��U*��9F��?o|�Q>/�`L�<�d�zN����}�E���s\�%�5����Ι���{~�d͞o�u!����Ş, @p�<�\�*�@��V3��7:����A�:��[���WI�����q�XT�_ �phg��}A�勢L)܇p�,��W��
{��X�)�*��u-,7��^��*W=Xz�U=�!��Baa��Z���3Y�����#�: @"�/*��e��s��~uK?���Z�����*2o-̍�����a�����'~�<?-��/k]��� �����
�;��!��N��[/�F����P H,���Х��9ao6��?�%5N\�]�5S ����Bm�a��i��ד��	�F�~��r=Vn�b�q(��H���|Q�%�K��É��n�\ʭ7>��gB  �
����Z7��Z��HX��}��6Ȁ�XX��-E�+��綰a�/�os&�x�S���(ʌj�Z�y�6�Ν_n���s-��E����r���P H$�s�����\�j����σ��\n�Ͻ��+��޲��\�
��_�����J��T�]����.���	jq�(�\NT���-�s�틋���R6�\ʍ[�Q*tB� $�r�D�f��ׅ�"���x��v���ܼ>y�߰��9Uf�\�P�ϛWX��w[F��s=�R��"4>H���'�Q�����!�_�ޯ,�K���:w)�r��R�Nu �D����Ԟ,~>��G�c�sH�z�
;~���h��}��\��y.X�\5�t�~��9�z˂|�(�P\��_E�m�P��ԝ�!��\ʭ�ߣb�Nu  Ĝ��V�e��>�x�r��;������[#���}��|(势O?�0_�\�$�)Q�?dY_~�B��~�iX[�P.�&�r�Nu!�>uڣ��6o�L]��OOO�xܺu묵��  ,n���?o�u7��,�^����-����(S#̇J�x�\�<�2��0.|�s�2���Z�F���+:!ԅh�@�����Y�k� �M����Q������Q�r�J�
�5쵪u���C�h�W��e��\ʍ�R��   Q5�)�r��@'�: !�Y�y�k�R��L��Kg���R���oO*e7   ��@'�: �\��L�ؼ�}���9t��ж�����iG.��J�]n   H�r��R��Oe��?�{���N��=8m�7���u����R�=�;  ���$�	����/�H6��3����qc�}�;�]��i@ >�y���͵س�Vʥ\ʭ�ܨ|�חr�ܰT�!B��А�>}�&e]u�U�?oܸ�ZZZܶH��A{{������Yss0�F٬�0ה�����-H�v���Z{�@����p�i@k�N����ǼW�}��C��K�+��܇>o�����[�Q�U�!B]T�����.yִ��ի�=nvv�2�L��)Ѝ�gz��e��U��7w�o���9� �  �C��Nu!���6�z��������B�̴��^�e���u����|��^���H�  �� ��6B��ު��A��C�͡Ӑ�0{�
)ح�������3   D"�@'�VBD%c!̡+��bvܿo���b�!�AI�Rn�1�R.�_nT2���[G�!�@'�v�m[p�����*t.���9��0L�D�Kgf�mbb�����͛��ň(�r)7�r������:*7hA:��Pw�С�ܷTP������fK�̀�L�gz#} �vg��ەJ�6`�$���٭[�R�T+Ɩ�G�r)�r�/7*)^_ʭ�r�F���u@�e��}m���>v���KoJQ���?��K��[�r����K�uTn��
t��w��dR�~��~cnJT�� ��R.�Rn�����K�uTn��t��w ��*���Kg�[2iBJ�?�'O�����ߺ��@��R.�Rnr�mM���[G�+�@'�}w �*k#Z}���}#�D9���sDK�t4��
�K���\S���[G喪�Nu@�e�V�-V�����   ��U�BPc�tf�bFA3E�  D-��      �tB�jl|.~�/�{����   *E�B     �@'�:���4۶q��
��L���  �"�   @��s�b1�K�l�   �u@��2@���   �H�:��b���ۖ�X�e���U�V�t�5k(�r)7F�F��חr�ܸ!�5�2�\{ߎ3�ܽ�b�9��5���x��u���i�\ʥ܈ˍ�^_ʭ�r�PD �uA*�.�׀���͛˾][[��^�Rʥ\ʭ�ܨ�����:*7�u@R)��mg_���݃Q>�u�����ЀT�ԫ�)�R.�V_nT���Rn�g�: "mM��i�p~�ξ�T*�׀�R����z����P.�Rn��F%��K�uTnꀈ�ޗ�G9���9��^:�"�N[ss��:u�r)�rVnTҼ��[G�&��P������L|c��,Wa2�vP�l6k333�K����r������:*7	u@��S�<�}=�o�p-���L�L   �B�T�n�hJ�� �)�5g��  ��: |��{��7���r�:  @}!�1�`�^�u�}k�؃_nUʝ}]��0�+:�n�=���/{̧:˟�>4�bώwX5(�r)��r����~�ߣ��Q/Z*���oߎ�Tf��7wTsn��t���H��K�	-7*���K�uTn��v͖�Y.��<k���y�_�|;mj��Դ#w�   ���1�����w6��Y��X*3�I�`�q�lӶ\�붬�h��~   @c �	�^���nwޕ!.e   h0��inS���    
e����&ԕ!�B�pvh    �IY(�R��PW����S��3    �3���GU6��c����}�y3    GC/'�����Dط{8�{��T���     G�GY>��Lc};�hch��   Ț�Ӣ�Q>B]F�3=M��   иr���o���� �Ub���ѝ}
v���   ����.�Nu�R�3�Yw߷v�RYO   @.���Lo�C.��4�����ξ�uM�#e���   P?�r�2��曻�[���kQ�f핹    IEND�B`�PK
     l`�[$7h�!  �!  /   images/a7fde0f7-2836-4f0c-aad0-66dcccec46ff.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     l`�[�W&��*  �*  /   images/b3e67e62-159a-497d-aba3-70fd70f56319.png�PNG

   IHDR   N   �   5�   gAMA  ���a   	pHYs  �  ��o�d  *#IDATx��}ip\ו��{7�Fc%v$����"�Z(J�,��%+��X�ؕrMy*I�&5����W*���5�Ԥj∶5�����D�Z(��. �  ������{.�`/�~�z%�SuQ�~���{�{�yZ��@L�!�(�ώỵ2�V���<Ո?]nE:��{Ct�4����ɴ����6��b(J�����Fa��#6ء4HZt�el�ȓ� qt����U�DXCM����3�&��'�Δ�`����DM�X��z	?���%�Kd�b��,�h@�����ޛ���H�~��"X�<��ƲM��8��Y\�˖�d���KZ�w��O�o��,m�V�F�/c�1����,_:u���8�2�J����M�^J�4�N++���3j��i��P��g{}~x|�_�`$aș�6.�V��V��������^�Q1qz2t������Ob`{jK�j0��aP�1=#�g`W�b����l���SD�A��"-=�_��������Pf�ä'-��O��ݓf��"
����˦���5�L�8�>��T��''N���U�>F-qI\�h|0 ���qk�6@5{�*;E��9��]D��ES0�T���T���r���[�u��O�V���/�9��j�d翂����1AZBJ���OĲ*"�͘�3*6I��b���9�rɣ�P�tj����Zt�._b��2���`V�,W��рnii�$��<ş�ȣ��:����ơb����Ec���b?�Ť��]GJV�p��o/Y<����.��3�+]�
� ]HVXIR��!���o.7��cL	E���%1Ar(���o2B*N��F3˖�������$� Y��>xf��D��A����B�Nh��B���k�����<���g��D��2Ub�8�H�8ZY�&��u�ˁ�PL�&37����re<PL�Zk�7��\�l�	��b�t9��iJ���=ޕ�o("��(M�o*�2��!K6qdTz�[�֑<
��!����:��,�8��~S�H �'1%ĭ +�)�
q
����{`t�B�A���_��W�	�>~�#3T�e���@�|'jT��(+AMY�l���a�����6F���֯�O�ǣ�e%.�1�Zg+�h+5�V+<�ˍ��8w�7U���
��X6∴m�V�ǟEi�tb0�q��n�V����x_;��0`9�,�i�Nlp��?��gc�������Oc��/q߰�˅e!�2ߏڀ�2�r���!�T*AR׬Y��vV���t�Vc��v���j��G]����|>?N��c<u�Bv������:n��z|���5����r �gչ�a��B���YKK+��Б����i���ذ�6���|[2`���aX�dCډ3�fQWj��j��k|�Y����.xl�%����q:�<<^a�^Q^�ڛ_a�i�u��a�7[`�A�`7��8�.�$�o����gv���}�����E�ǖ����:��Bډ�1���D?_����bA�~#_��i'N��@��!Q�u,���v��v��Z&qI N��.$�	�w��6U���[���Z2�jܹ	�u��A�~#[�Xq`"H;qY?��§���Ƈ׻p�]�ˏ����c���"ژp��}�$.@���ѱ1\�̓7ka1��\���
�c�ej}X.��V�E�jN�;�8�X<�����ܵ�����NI��+��6m܀��ȸsM �j։�&:&���qP���h$�9t� �l��������dU��G��d�yM�XP���ju�f�U�i#���n�84��d��Pn6Ð����!�)'������F�9������ǹ[��e�Z�BC�Ʉ�%%��kqϕ����,3�VVbr~���wz�+u1LLL�w�� 2�^�}p?z�9X,�S�l�c��ɐ�-k*��1���S��w'�Bʈ+g�bw���/JM�ũYFq}��݋��}0mm��8��Ӌm[��e.	�f�9��tH^J���(����%N�,�I�^�csy�{�C�j�K�'�ɺzN���$n�� UH:q�A��&?�Ȝ�S�ԬǕ;���3Gه���?+z<���p�L�>"�TJ^R�J�I����:��HVV~��g���U��uG�Aw_,��愉�[S���><���T�h�����0���SJؼI��i�V�u�B%/H
q4H���K�8���|iw$�4�oJ�΂+�'u�&U���I�N���P����T�?	OOy��ǐ�%�LzãE\�,�6�^:*0<)�χ���E��8o4�g�j����OS��nF��4����E^��Ք�Ĕ� ���0--m8wo-��|�J;�z�� h���͈�>��GnJ2E�đ��`1OpI�p��vx4zhsK�w;�37-� ��MUJS�IZ2EB�Q�N�C��8�h����[K;��\�	��t����9�-\��Kd((� ?3Q$D\h�#�d���т�4�[�a)�bG��Ousn��D��uى��F�ፄu~Zr��P]]�_r@δ}~�3| iKV��8R�d�F��d5)"H�8��� �doM'�AQ�?�_B���OrCc�S�Z{Pɨ��}�e@���\W�>7�&v����g���L���َ��͒�g��1;7�̜bY�HV�N1qd��1�c�X��)yLgg�|�*޻3���g���Xx��̲��&eG�Ur��<x�D��8�B�:Nc�����1���ۿ�?o��#���Y2Mx`�A<��jU��du�̪q�R�JgFrss���]�Y�֚g���{��Jx��%�� ���đu���8���[���ƍ�x~|���>^�&f���ū*���U�Ѵp�lS5^���P���C�öm��mQ�l�}|�9�Y�5$4�e5�G�]:����R+����h�/?��!ũ����>�B��o#*dR��Y!�%/�����%/[�U�J�����.?v�ՠ�@��1�h�i��S�B.Z�M	�#D�rr\���a6U�$�g����!�骸q�q����/I֒PF��,p4Mi�7�̄b r&�f��¤�I�Xzzzq�]�iS�;7�EOo/��l�I���0r�923��uH�绗�8(X��k"���>F�_��5Z��7�A3kw���``7�b�⋳���g^�$w�,$Dݹ`2S$iD��hv�EKX���Y����aq�1��<'���K~ga�ֿt�=��	�Gӳ<���I��B�h������_2�I0ge�g��@ww7�j���J.`HǙ�RI7�$o��ǰv]�>.�$	Gw�^��?T�BA���XU�ɈM����3�J�(��o:?ݰ�λKҗ�:��-Hi�R� TI�	�N+�S�n����7�?����0��_I�,�9�̎�~��vԸ��r@�Z��^�ϤT����ᨆzt#V��a�$�'TR��l�"؏�j��svr|���z���1j�07Ώ��m8�Ò�!�KӥL�������E�D�=�?I�jm��K�8��'D���Y��4�Q_Kk�=E@͓������z�gM�����jaL�l0m��@���M���T2��%D�i�u;PX��**q���fc�(��]f������ �-����؝6�k�W���w��5u����k�(GM�"ISg����t!��j�����Te�l:�\�6Â9g ��P����31���2ŕ��*�)Z^1\�M)!Oq$���ֈ,����+��WH<H%��ء��:~��b�01�e��=(*Z�{:^Һ��
�L3j�J0i����'D�6#'���qGj�H�DEnxF�J�3�j}�:��dY��$�5�36tCuL�<��a�9�Za�ܮX��M�0d֔����E%���䮩�"ˤ%Q�z�$.��o�E���v�?���(��Q<e��xw�^#�I���R�L	��RG���h�$���<,��% Oy4e�z��F�q]�w&B�1��n�+F���[$�x��۰�x`�L���LM�1�ٔ���vM)%��-ұ$�F.Y1��\�kVKU'�5k*�4����f����I4��躹�� %�3�M\d�a�6R�\��/�x&:����T"�>44�{����0'���~TTT`�����
�|Q�*��&���3�Q�y𦒥�;�ʎu#^�$.z�^#�9i��,L�wv����������믑�����Z�ݻW𸾾>~���<<�u뢭���?aN�К�]J+ј�ٔ��"%��=A��4�/t�L������R����5��!��
�X�l7q��}����{�=ޡ�ĉ1sn�W��/�Ӊ����K����Î��\���8�ٻp���R�3ª��㵻��#LŤ<���g���X�"����BgZܣ�QA3|�qt��m�eE�X���Ř��n�P��v���رc���H�h4�ȑ#��>�z�-����a�!� �gE�<�m�n��������v2C����s~9̲��ͱ��[mĀ#v_qCC�h��%��U��v�3�T����=o�H;t�V�����uff&�~�m��F���i1{����w�P�:Q|u����wаg�h	Fq�ͷ��t�w��{��?��صkWB�Q^^�.Ԇ>��O�d 33��V�����6^����0#�D�͛M������EM�d��ݻ0��LU
~NS�����&P;[*{-..f���xE�$o`` ���l�V'u�%l�=w�(>��K4^������q⺺�����s�=�)5�󯱓���+��ݸq�_|}}=�m�����0�*rG�l�^_%+{�ԩ�G�ť��:���AA~���3N\��k\SEZgg'���.J[ʟ~�i���{��t��;�<�b�����Af�c������];p��z8q�K�B���W�;w�`���Q�ONN2i�������3g��U�'�|r�����ܹs�G���7rU�
���jm��Km�u������ᶰ���qR��q
�Qho��J�t�X�lzz�;���r�
wK"A����H�T�z�j�$�� ��2���=,
Q��;::y�NJ�F�V�褏q�D���vn�u���'�}�G�I౵���+/��|t�ڧا�Bh����C��������,�frA����ۂ�Dk<Ǣ�w?8�9S%O��=��O#�O�>��~̸UX���O<��5a�Cd��>���Z�6&��%����5�V[��i�h�X��6Ƭ_��,�7-�Q^�j4߻E9��F�͜�Л@A4�)F}�� A�&��AK���1�Y�B87�{��z��,$^�����g�6�7�F���Qđ�h�?\�ЪD���R띇���{�{A�}~�!n�Z��.)�Mz�JMMM-}��xx��M]�uY�;<i��#8�]0����}n���Ha����^Oy_k`"K����k+Q��5�jL�;���ȳAP�Ԫ-��>ì���ͨ�=M�R��E����K�s�:��1ק���_�_�K��v'��M��aZ]>������sK�S[������Ű͇�-��G�`PTa�%����/��UB����̕ �P�B�����;��w�a�ڍҺZ�qG�.F�b�T��*��&	�7�[��?y�)^�IRS���E������QԮo�-��Y1M	�2<,��R���@�+ ��^bа��uk�%��bѿ�hhh�~܁ ���a.JD�T&��R�ed(ĺ���7�\�ʥ��6T�7�����MqU{���)��z��E��� (	YPx��-�D`����}?� B�ر��c�F�	�w����M,�����uuu���-�=��8�<���I��4T2)�mjj�Ⱦ}��	�9~�Y�8��t�k7����>7�۷o�Y�^\�҈�{R2 �� ��ȣ`��[rS��������������&T���(az�&�\wɟ8r�0>9s_^��=�]!�+���<y�Y�5�QM����ɨeDBA	 z�Ź����ï^]��):��D��g�l���#��;�Y�X���^x������_�
�H#"Z����k�%m|�[���&��.&@��κDe���i�CoƯ���a��K��k�m�Di^�	�x���~��6eT�m�`cUE�Z�W�����?s)�'�
���(.\��o�PF�
���o����BA�sz��.�P��[��<ӧ�� �|����dŻ��CV�����,�c��������B��ݍ���و -�L��VW3�Ww����<~��/��"ϱQm�֭������ū����Q���W_�J�μMP���K�0�u~�,���Ew��Kn	��	�\��B�J���/an#.?����Z��a)��l+��|	��/q�h��E:��7��ŋ��?��+^2b"(�hmm�y�M�6E�3q�/pӾƺ}���^�2�SqÃţ������E���&8*^�"���|��Qx�{wD?f�_z���裏�ĐA&
Ղ� �4D�n�hB�#Ƶ�D��{�|5�ʾ��Mdg,ݸ���E�m��US%���Q�-�O	�(A7��r-YU2z�[�o��m�k�*�.�����$E^��&N#P:@��MY9\�j�J��,}�\��>���ٸK�6֞�H�W��dAmގt��4;� ��c��.%�qU+EI#qn��W�K�d�)'�8%�L�]%��Pa�g�wx����)A\�ѝ�|lp��l�I�B!_֢�{5S�4S'�m�:#����јn�Ȍ����K_E&=K�XVc��k���@5(�"έ��R�*�]n8�9") ��q�B
	|FԊ�$�v��^�LӀ����;�y.��Š�$�V�i5���`ˆu�i� �.'Tڇ7�,gA��K��+��@�eV�G"PD��v�P]Yym��ʼq��榨tF��b?jll��SE�Snw�������ƴ���U`R��mz4�4�R�
Ņ��먫`d��t�u�V�CF�B���ủ�����Ma�d�^J�L��,J�IeT<�m�\TyI�Ý���'!c͎���H��9�#"ɣw�{��t���d*�62�Բ���m�c��t��<8�����S`���d��ǚ�ɣ��H�A�ʴ�`�X�qo�-��5�hj���V5>d��X8v$��Fgf1�q��[���H����z"�v����A��S�h�	��b7N�H�������j9�]�[V���w�?��]�NO:-��d��`k_(z���q���%x�󘞑ײ��^n��A<��,Υ	pјH����mا7�łl��A��N&4�����B|=� 
e�9�9½8rn��4���r�h���m��N23��Y��|z�8�����A>��c�2**5���9z�� ��X��ڑ�ulj�&����󋔪0�ϩew��4W��K��K�K6$u2�j���X�\rt�Ϛi����ܻf(`���)E���u-�gv�=��������@dk�r�����D��8�=q��EJ���^�Cb�8cĸ������>_>-Q��\�.�H)PU����U���c�*�+��,�t3�����ŹcH�����1ܸ�Rk���aU�t��b��N����r �8��Kl���CWg�d�U�������,���	6n����9G��$�IÐ�4b�0�)�4�1k��� ��o�,���6U�	�e�`djnis^:�6����"c����8��ud8�g;�m��[�z=���i�8�H)�wt���a��kh��bz�W����F����8��Z54�}��������e�vI�#�c�0ݼ��w��]�/`��I�f�m�SUŢ��z/�8�4F7����T(&ΤW#Sz�U00"��9�7jO5]���t�ټ�<��/�ی �GV�܉|���P���H��}ߤװJ�
zv�:M��i~�r�g����v�A��ц�ϧ�t���I'N�ْ�K�v9���E3V��T5����� z����U���8�>F�O&uvO ������E����B����O+O)iè#�a�L��wz��)"N��wL�v���Hde�.,����y����isa'�&x*��v�yk�f������YT����9N���2��ĸc^_�t�A��1sr��6sxfgQ�{�䂴��]�B��I�"�s����|0H4�r��
�� �
�?x�Н�4�Z�>���/��'��$�S	<������%A��H���͚cV3��$����8�[X��4Zx��BD����A��Y�M-t���ӌ��~Q�ȡ�wo��q��0i��H�����I̗S�ǹ�ɧ؋`R�T�L���0S�N�=OSPH�0��K�Zq��"�ZbG���@7��:&y��\�x��(I$r9�E@-���T���O`*'z��*��A4���cW��F���G
�H_"�a�!-q䷽��7y	U�Ӧ3��o/E��ǩ���gJ'V�j~I�䀦ꔕ�Uj�WHAq��W��s�6+�kk��#d��B�*�_ʺy�.D����"�^X����ȐFQg
��i74��<T�{���A	�2!^�&��]����i�%2���$����߹'^}Y|��ǻ��1�x H\y~6L����J-IeH���_|����|��ڶ�a�Ȃ49������cAT�^ڷ�_nM*y|�AªRI�!�X�Ԕd����U0�(~y<��]Q���}yOm)��O���s�p[�y҂��M�a`��}b�;{�b��=��.�����
�h�)KL�5���,�������
�����O�r�h���$��38��lٗ�]�RH��r��e���Ժ�R�45����r ��Qc ��ˉ���q����n��8s����Y����a�U��f$�������v6�
���u���s�33���ޡB������H�]�����O�sEu�
�z����y��S�M�S�����"A�2M����b��'ǲ�EZ�sv7CǤ�W!�u���6d-�rS7�P���*�[�����з�8%�J!��oGFy9�ns�+ܹ�7>�MI�k�KXǭ&Tm݉t"��9zn���`jjZpVmm5&_<��ټ&o�3O�F���bQÂ��h���4Gڈ��u8{o���,�u|���غmώHu�5�.>�m9�\���fG��~��ws����;�455�X�t빴G�����Ô�xƖ�.9g��.��'�Uϥ���/�����V��̊784�k�ݳsؼ{�E~A�V�!+\����B� *�`����(�|�wП����i}�Y�����ѥ^n�<�!��ҭ��B���'K��R��<����O�"wz��L�-� -D���\�D#���y�i!.8M	f�����т�6dAڣш>x��jOx����	�~K��92���sC<�}����{O<�)���/g�Z�ދ޻J=��LW�#�r6~r����i��)'�;;��*��w��x;���R������{A���=�Ђ���70�|:ot>]nIJ�#�0�L���:'�._@u�֨N�T�TS#��r��ݽ�S����kU|-�!�ą�P��p�p�ˋ8���Z;f��B��̈��P���s��s)%.r��b�����Y�S��`O�N�Z[
�����khس��,�����ݏH�[���8�iD�o�:�������.^Bqa,f3,e�<�I�JF��e�Ӳj���1����E	�#�;�\ʈuz#A�q����u���ŕ��p��P/�m�MM��v��_�5��>�r�ĉI�?�2���!k�Ѩ��2�?��b5<�Y�@߹�۶���~:���'�ߌk7{R}:�֔'��h��$��6鱩o�b��~K&r�JE-+E2�zJ�4⺻���768ğwcԩ���P�� ����m�Z3K��{��=�o����3���
�bzɻ�s�j~�xJ�:766�ܝ�>0)��#?�}�S�.����"��3���t�Q�[��1#�<����GF�?39�I�.�4ó��ۿE�y��!-^��ǯ3w�{H&����x�ߣ�+�ɝHݚc���p�4bXD����z����~��_^Q!�>%H�8zt��ӑ%�ԕ�$�)N���+�)�
q
�B�B��+�)�
q
�B�B��I'�J������~_x�O�t�bu�I'���$��T�{���b�8�X!N!V�S��b�8�X!N!V�S��")ĥ2�I�=Ƅ����x�G/7����8���؏䓃�HeC��x�G+:N!�N��l��>�����\�������x��h�E꩜��F����{N*�T������9qb$<x���#��D"M��O���!�0���b7�ʼe?�:^$�8���/R(L����Dm�USY�bϥH���������j
"����_#���TGG�� ��cY^"���B��yT��"��B�?	D%��`�7,L��qY"3�r�5��="3��+VU!V�S��maS'��I�>SSS���|Rp��h�j������zoo/��"!�G5���ޗj*O�uuu	.I��S�S�#8���`�u���4$mtL$y$iDId����BM�Ȋ�w�C5߂G��EZ,���C�w�<4=����w�8$�=I�8
��[�֔�D@ӝB:��� a�jjj��;�|�$�,�dy�0<4�7~�&�Z�,$e����}���q������g���    IEND�B`�PK
     l`�[�W&��*  �*  /   images/ab942d8a-eab6-45a7-8f5a-30ef729b6f10.png�PNG

   IHDR   N   �   5�   gAMA  ���a   	pHYs  �  ��o�d  *#IDATx��}ip\ו��{7�Fc%v$����"�Z(J�,��%+��X�ؕrMy*I�&5����W*���5�Ԥj∶5�����D�Z(��. �  ������{.�`/�~�z%�SuQ�~���{�{�yZ��@L�!�(�ώỵ2�V���<Ո?]nE:��{Ct�4����ɴ����6��b(J�����Fa��#6ء4HZt�el�ȓ� qt����U�DXCM����3�&��'�Δ�`����DM�X��z	?���%�Kd�b��,�h@�����ޛ���H�~��"X�<��ƲM��8��Y\�˖�d���KZ�w��O�o��,m�V�F�/c�1����,_:u���8�2�J����M�^J�4�N++���3j��i��P��g{}~x|�_�`$aș�6.�V��V��������^�Q1qz2t������Ob`{jK�j0��aP�1=#�g`W�b����l���SD�A��"-=�_��������Pf�ä'-��O��ݓf��"
����˦���5�L�8�>��T��''N���U�>F-qI\�h|0 ���qk�6@5{�*;E��9��]D��ES0�T���T���r���[�u��O�V���/�9��j�d翂����1AZBJ���OĲ*"�͘�3*6I��b���9�rɣ�P�tj����Zt�._b��2���`V�,W��рnii�$��<ş�ȣ��:����ơb����Ec���b?�Ť��]GJV�p��o/Y<����.��3�+]�
� ]HVXIR��!���o.7��cL	E���%1Ar(���o2B*N��F3˖�������$� Y��>xf��D��A����B�Nh��B���k�����<���g��D��2Ub�8�H�8ZY�&��u�ˁ�PL�&37����re<PL�Zk�7��\�l�	��b�t9��iJ���=ޕ�o("��(M�o*�2��!K6qdTz�[�֑<
��!����:��,�8��~S�H �'1%ĭ +�)�
q
����{`t�B�A���_��W�	�>~�#3T�e���@�|'jT��(+AMY�l���a�����6F���֯�O�ǣ�e%.�1�Zg+�h+5�V+<�ˍ��8w�7U���
��X6∴m�V�ǟEi�tb0�q��n�V����x_;��0`9�,�i�Nlp��?��gc�������Oc��/q߰�˅e!�2ߏڀ�2�r���!�T*AR׬Y��vV���t�Vc��v���j��G]����|>?N��c<u�Bv������:n��z|���5����r �gչ�a��B���YKK+��Б����i���ذ�6���|[2`���aX�dCډ3�fQWj��j��k|�Y����.xl�%����q:�<<^a�^Q^�ڛ_a�i�u��a�7[`�A�`7��8�.�$�o����gv���}�����E�ǖ����:��Bډ�1���D?_����bA�~#_��i'N��@��!Q�u,���v��v��Z&qI N��.$�	�w��6U���[���Z2�jܹ	�u��A�~#[�Xq`"H;qY?��§���Ƈ׻p�]�ˏ����c���"ژp��}�$.@���ѱ1\�̓7ka1��\���
�c�ej}X.��V�E�jN�;�8�X<�����ܵ�����NI��+��6m܀��ȸsM �j։�&:&���qP���h$�9t� �l��������dU��G��d�yM�XP���ju�f�U�i#���n�84��d��Pn6Ð����!�)'������F�9������ǹ[��e�Z�BC�Ʉ�%%��kqϕ����,3�VVbr~���wz�+u1LLL�w�� 2�^�}p?z�9X,�S�l�c��ɐ�-k*��1���S��w'�Bʈ+g�bw���/JM�ũYFq}��݋��}0mm��8��Ӌm[��e.	�f�9��tH^J���(����%N�,�I�^�csy�{�C�j�K�'�ɺzN���$n�� UH:q�A��&?�Ȝ�S�ԬǕ;���3Gه���?+z<���p�L�>"�TJ^R�J�I����:��HVV~��g���U��uG�Aw_,��愉�[S���><���T�h�����0���SJؼI��i�V�u�B%/H
q4H���K�8���|iw$�4�oJ�΂+�'u�&U���I�N���P����T�?	OOy��ǐ�%�LzãE\�,�6�^:*0<)�χ���E��8o4�g�j����OS��nF��4����E^��Ք�Ĕ� ���0--m8wo-��|�J;�z�� h���͈�>��GnJ2E�đ��`1OpI�p��vx4zhsK�w;�37-� ��MUJS�IZ2EB�Q�N�C��8�h����[K;��\�	��t����9�-\��Kd((� ?3Q$D\h�#�d���т�4�[�a)�bG��Ousn��D��uى��F�ፄu~Zr��P]]�_r@δ}~�3| iKV��8R�d�F��d5)"H�8��� �doM'�AQ�?�_B���OrCc�S�Z{Pɨ��}�e@���\W�>7�&v����g���L���َ��͒�g��1;7�̜bY�HV�N1qd��1�c�X��)yLgg�|�*޻3���g���Xx��̲��&eG�Ur��<x�D��8�B�:Nc�����1���ۿ�?o��#���Y2Mx`�A<��jU��du�̪q�R�JgFrss���]�Y�֚g���{��Jx��%�� ���đu���8���[���ƍ�x~|���>^�&f���ū*���U�Ѵp�lS5^���P���C�öm��mQ�l�}|�9�Y�5$4�e5�G�]:����R+����h�/?��!ũ����>�B��o#*dR��Y!�%/�����%/[�U�J�����.?v�ՠ�@��1�h�i��S�B.Z�M	�#D�rr\���a6U�$�g����!�骸q�q����/I֒PF��,p4Mi�7�̄b r&�f��¤�I�Xzzzq�]�iS�;7�EOo/��l�I���0r�923��uH�绗�8(X��k"���>F�_��5Z��7�A3kw���``7�b�⋳���g^�$w�,$Dݹ`2S$iD��hv�EKX���Y����aq�1��<'���K~ga�ֿt�=��	�Gӳ<���I��B�h������_2�I0ge�g��@ww7�j���J.`HǙ�RI7�$o��ǰv]�>.�$	Gw�^��?T�BA���XU�ɈM����3�J�(��o:?ݰ�λKҗ�:��-Hi�R� TI�	�N+�S�n����7�?����0��_I�,�9�̎�~��vԸ��r@�Z��^�ϤT����ᨆzt#V��a�$�'TR��l�"؏�j��svr|���z���1j�07Ώ��m8�Ò�!�KӥL�������E�D�=�?I�jm��K�8��'D���Y��4�Q_Kk�=E@͓������z�gM�����jaL�l0m��@���M���T2��%D�i�u;PX��**q���fc�(��]f������ �-����؝6�k�W���w��5u����k�(GM�"ISg����t!��j�����Te�l:�\�6Â9g ��P����31���2ŕ��*�)Z^1\�M)!Oq$���ֈ,����+��WH<H%��ء��:~��b�01�e��=(*Z�{:^Һ��
�L3j�J0i����'D�6#'���qGj�H�DEnxF�J�3�j}�:��dY��$�5�36tCuL�<��a�9�Za�ܮX��M�0d֔����E%���䮩�"ˤ%Q�z�$.��o�E���v�?���(��Q<e��xw�^#�I���R�L	��RG���h�$���<,��% Oy4e�z��F�q]�w&B�1��n�+F���[$�x��۰�x`�L���LM�1�ٔ���vM)%��-ұ$�F.Y1��\�kVKU'�5k*�4����f����I4��躹�� %�3�M\d�a�6R�\��/�x&:����T"�>44�{����0'���~TTT`�����
�|Q�*��&���3�Q�y𦒥�;�ʎu#^�$.z�^#�9i��,L�wv����������믑�����Z�ݻW𸾾>~���<<�u뢭���?aN�К�]J+ј�ٔ��"%��=A��4�/t�L������R����5��!��
�X�l7q��}����{�=ޡ�ĉ1sn�W��/�Ӊ����K����Î��\���8�ٻp���R�3ª��㵻��#LŤ<���g���X�"����BgZܣ�QA3|�qt��m�eE�X���Ř��n�P��v���رc���H�h4�ȑ#��>�z�-����a�!� �gE�<�m�n��������v2C����s~9̲��ͱ��[mĀ#v_qCC�h��%��U��v�3�T����=o�H;t�V�����uff&�~�m��F���i1{����w�P�:Q|u����wаg�h	Fq�ͷ��t�w��{��?��صkWB�Q^^�.Ԇ>��O�d 33��V�����6^����0#�D�͛M������EM�d��ݻ0��LU
~NS�����&P;[*{-..f���xE�$o`` ���l�V'u�%l�=w�(>��K4^������q⺺�����s�=�)5�󯱓���+��ݸq�_|}}=�m�����0�*rG�l�^_%+{�ԩ�G�ť��:���AA~���3N\��k\SEZgg'���.J[ʟ~�i���{��t��;�<�b�����Af�c������];p��z8q�K�B���W�;w�`���Q�ONN2i�������3g��U�'�|r�����ܹs�G���7rU�
���jm��Km�u������ᶰ���qR��q
�Qho��J�t�X�lzz�;���r�
wK"A����H�T�z�j�$�� ��2���=,
Q��;::y�NJ�F�V�褏q�D���vn�u���'�}�G�I౵���+/��|t�ڧا�Bh����C��������,�frA����ۂ�Dk<Ǣ�w?8�9S%O��=��O#�O�>��~̸UX���O<��5a�Cd��>���Z�6&��%����5�V[��i�h�X��6Ƭ_��,�7-�Q^�j4߻E9��F�͜�Л@A4�)F}�� A�&��AK���1�Y�B87�{��z��,$^�����g�6�7�F���Qđ�h�?\�ЪD���R띇���{�{A�}~�!n�Z��.)�Mz�JMMM-}��xx��M]�uY�;<i��#8�]0����}n���Ha����^Oy_k`"K����k+Q��5�jL�;���ȳAP�Ԫ-��>ì���ͨ�=M�R��E����K�s�:��1ק���_�_�K��v'��M��aZ]>������sK�S[������Ű͇�-��G�`PTa�%����/��UB����̕ �P�B�����;��w�a�ڍҺZ�qG�.F�b�T��*��&	�7�[��?y�)^�IRS���E������QԮo�-��Y1M	�2<,��R���@�+ ��^bа��uk�%��bѿ�hhh�~܁ ���a.JD�T&��R�ed(ĺ���7�\�ʥ��6T�7�����MqU{���)��z��E��� (	YPx��-�D`����}?� B�ر��c�F�	�w����M,�����uuu���-�=��8�<���I��4T2)�mjj�Ⱦ}��	�9~�Y�8��t�k7����>7�۷o�Y�^\�҈�{R2 �� ��ȣ`��[rS��������������&T���(az�&�\wɟ8r�0>9s_^��=�]!�+���<y�Y�5�QM����ɨeDBA	 z�Ź����ï^]��):��D��g�l���#��;�Y�X���^x������_�
�H#"Z����k�%m|�[���&��.&@��κDe���i�CoƯ���a��K��k�m�Di^�	�x���~��6eT�m�`cUE�Z�W�����?s)�'�
���(.\��o�PF�
���o����BA�sz��.�P��[��<ӧ�� �|����dŻ��CV�����,�c��������B��ݍ���و -�L��VW3�Ww����<~��/��"ϱQm�֭������ū����Q���W_�J�μMP���K�0�u~�,���Ew��Kn	��	�\��B�J���/an#.?����Z��a)��l+��|	��/q�h��E:��7��ŋ��?��+^2b"(�hmm�y�M�6E�3q�/pӾƺ}���^�2�SqÃţ������E���&8*^�"���|��Qx�{wD?f�_z���裏�ĐA&
Ղ� �4D�n�hB�#Ƶ�D��{�|5�ʾ��Mdg,ݸ���E�m��US%���Q�-�O	�(A7��r-YU2z�[�o��m�k�*�.�����$E^��&N#P:@��MY9\�j�J��,}�\��>���ٸK�6֞�H�W��dAmގt��4;� ��c��.%�qU+EI#qn��W�K�d�)'�8%�L�]%��Pa�g�wx����)A\�ѝ�|lp��l�I�B!_֢�{5S�4S'�m�:#����јn�Ȍ����K_E&=K�XVc��k���@5(�"έ��R�*�]n8�9") ��q�B
	|FԊ�$�v��^�LӀ����;�y.��Š�$�V�i5���`ˆu�i� �.'Tڇ7�,gA��K��+��@�eV�G"PD��v�P]Yym��ʼq��榨tF��b?jll��SE�Snw�������ƴ���U`R��mz4�4�R�
Ņ��먫`d��t�u�V�CF�B���ủ�����Ma�d�^J�L��,J�IeT<�m�\TyI�Ý���'!c͎���H��9�#"ɣw�{��t���d*�62�Բ���m�c��t��<8�����S`���d��ǚ�ɣ��H�A�ʴ�`�X�qo�-��5�hj���V5>d��X8v$��Fgf1�q��[���H����z"�v����A��S�h�	��b7N�H�������j9�]�[V���w�?��]�NO:-��d��`k_(z���q���%x�󘞑ײ��^n��A<��,Υ	pјH����mا7�łl��A��N&4�����B|=� 
e�9�9½8rn��4���r�h���m��N23��Y��|z�8�����A>��c�2**5���9z�� ��X��ڑ�ulj�&����󋔪0�ϩew��4W��K��K�K6$u2�j���X�\rt�Ϛi����ܻf(`���)E���u-�gv�=��������@dk�r�����D��8�=q��EJ���^�Cb�8cĸ������>_>-Q��\�.�H)PU����U���c�*�+��,�t3�����ŹcH�����1ܸ�Rk���aU�t��b��N����r �8��Kl���CWg�d�U�������,���	6n����9G��$�IÐ�4b�0�)�4�1k��� ��o�,���6U�	�e�`djnis^:�6����"c����8��ud8�g;�m��[�z=���i�8�H)�wt���a��kh��bz�W����F����8��Z54�}��������e�vI�#�c�0ݼ��w��]�/`��I�f�m�SUŢ��z/�8�4F7����T(&ΤW#Sz�U00"��9�7jO5]���t�ټ�<��/�ی �GV�܉|���P���H��}ߤװJ�
zv�:M��i~�r�g����v�A��ц�ϧ�t���I'N�ْ�K�v9���E3V��T5����� z����U���8�>F�O&uvO ������E����B����O+O)iè#�a�L��wz��)"N��wL�v���Hde�.,����y����isa'�&x*��v�yk�f������YT����9N���2��ĸc^_�t�A��1sr��6sxfgQ�{�䂴��]�B��I�"�s����|0H4�r��
�� �
�?x�Н�4�Z�>���/��'��$�S	<������%A��H���͚cV3��$����8�[X��4Zx��BD����A��Y�M-t���ӌ��~Q�ȡ�wo��q��0i��H�����I̗S�ǹ�ɧ؋`R�T�L���0S�N�=OSPH�0��K�Zq��"�ZbG���@7��:&y��\�x��(I$r9�E@-���T���O`*'z��*��A4���cW��F���G
�H_"�a�!-q䷽��7y	U�Ӧ3��o/E��ǩ���gJ'V�j~I�䀦ꔕ�Uj�WHAq��W��s�6+�kk��#d��B�*�_ʺy�.D����"�^X����ȐFQg
��i74��<T�{���A	�2!^�&��]����i�%2���$����߹'^}Y|��ǻ��1�x H\y~6L����J-IeH���_|����|��ڶ�a�Ȃ49������cAT�^ڷ�_nM*y|�AªRI�!�X�Ԕd����U0�(~y<��]Q���}yOm)��O���s�p[�y҂��M�a`��}b�;{�b��=��.�����
�h�)KL�5���,�������
�����O�r�h���$��38��lٗ�]�RH��r��e���Ժ�R�45����r ��Qc ��ˉ���q����n��8s����Y����a�U��f$�������v6�
���u���s�33���ޡB������H�]�����O�sEu�
�z����y��S�M�S�����"A�2M����b��'ǲ�EZ�sv7CǤ�W!�u���6d-�rS7�P���*�[�����з�8%�J!��oGFy9�ns�+ܹ�7>�MI�k�KXǭ&Tm݉t"��9zn���`jjZpVmm5&_<��ټ&o�3O�F���bQÂ��h���4Gڈ��u8{o���,�u|���غmώHu�5�.>�m9�\���fG��~��ws����;�455�X�t빴G�����Ô�xƖ�.9g��.��'�Uϥ���/�����V��̊784�k�ݳsؼ{�E~A�V�!+\����B� *�`����(�|�wП����i}�Y�����ѥ^n�<�!��ҭ��B���'K��R��<����O�"wz��L�-� -D���\�D#���y�i!.8M	f�����т�6dAڣш>x��jOx����	�~K��92���sC<�}����{O<�)���/g�Z�ދ޻J=��LW�#�r6~r����i��)'�;;��*��w��x;���R������{A���=�Ђ���70�|:ot>]nIJ�#�0�L���:'�._@u�֨N�T�TS#��r��ݽ�S����kU|-�!�ą�P��p�p�ˋ8���Z;f��B��̈��P���s��s)%.r��b�����Y�S��`O�N�Z[
�����khس��,�����ݏH�[���8�iD�o�:�������.^Bqa,f3,e�<�I�JF��e�Ӳj���1����E	�#�;�\ʈuz#A�q����u���ŕ��p��P/�m�MM��v��_�5��>�r�ĉI�?�2���!k�Ѩ��2�?��b5<�Y�@߹�۶���~:���'�ߌk7{R}:�֔'��h��$��6鱩o�b��~K&r�JE-+E2�zJ�4⺻���768ğwcԩ���P�� ����m�Z3K��{��=�o����3���
�bzɻ�s�j~�xJ�:766�ܝ�>0)��#?�}�S�.����"��3���t�Q�[��1#�<����GF�?39�I�.�4ó��ۿE�y��!-^��ǯ3w�{H&����x�ߣ�+�ɝHݚc���p�4bXD����z����~��_^Q!�>%H�8zt��ӑ%�ԕ�$�)N���+�)�
q
�B�B��+�)�
q
�B�B��I'�J������~_x�O�t�bu�I'���$��T�{���b�8�X!N!V�S��b�8�X!N!V�S��")ĥ2�I�=Ƅ����x�G/7����8���؏䓃�HeC��x�G+:N!�N��l��>�����\�������x��h�E꩜��F����{N*�T������9qb$<x���#��D"M��O���!�0���b7�ʼe?�:^$�8���/R(L����Dm�USY�bϥH���������j
"����_#���TGG�� ��cY^"���B��yT��"��B�?	D%��`�7,L��qY"3�r�5��="3��+VU!V�S��maS'��I�>SSS���|Rp��h�j������zoo/��"!�G5���ޗj*O�uuu	.I��S�S�#8���`�u���4$mtL$y$iDId����BM�Ȋ�w�C5߂G��EZ,���C�w�<4=����w�8$�=I�8
��[�֔�D@ӝB:��� a�jjj��;�|�$�,�dy�0<4�7~�&�Z�,$e����}���q������g���    IEND�B`�PK
     l`�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     l`�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     l`�[����s  �s                   cirkitFile.jsonPK 
     l`�[                        �s  jsons/PK 
     l`�[�5zU                 t  jsons/user_defined.jsonPK 
     l`�[                        W�  images/PK 
     l`�[�R�W�  W�  /             |�  images/e30496d1-6e1c-40fa-a66f-2add70ecdc94.pngPK 
     l`�[$7h�!  �!  /              6 images/a7fde0f7-2836-4f0c-aad0-66dcccec46ff.pngPK 
     l`�[�W&��*  �*  /             ^X images/b3e67e62-159a-497d-aba3-70fd70f56319.pngPK 
     l`�[�W&��*  �*  /             ,� images/ab942d8a-eab6-45a7-8f5a-30ef729b6f10.pngPK 
     l`�[�c��f  �f  /             �� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     l`�[��EM  M  /             ( images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK    
 
   �(   