PK
     $s�[����E �E    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-neg"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-pos"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20":["pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_0"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_24"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28":["pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_3"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29":["pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_0"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_26"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-neg","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_2"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_1"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-neg"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_23"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-neg","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_1"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-pos","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_2"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_0"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-pos","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_2"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-neg","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_3"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_20","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_2"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_19","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_1"],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62":[],"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_0"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-pos":["pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_1"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-neg":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-pos":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-neg":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-pos":["pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_1"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-neg":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-pos":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-neg":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-pos":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-neg":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61_polarity-neg":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-pos":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-neg":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5"],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62_polarity-pos":[],"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62_polarity-neg":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_0":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_1":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_2":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_3":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-pos"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-neg"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_7":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_0"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_9":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_1"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_10":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_2"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_11":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_3"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_12":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_5"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_13":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_6"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_14":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_15":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_16":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_17":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_18":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_7"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_19":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_20":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_21":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_4"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_22":["pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_0"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_23":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_24":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_25":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_26":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_28":["pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_0"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_29":["pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_1"],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_30":[],"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_31":[],"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_0":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62"],"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_1":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61"],"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_2":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60"],"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_3":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59"],"pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_0":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55"],"pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_1":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_29"],"pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_2":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56"],"pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_0":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_28"],"pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_1":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52"],"pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_2":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53"],"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_0":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8"],"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_1":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_9"],"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_2":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_10"],"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_3":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_11"],"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_4":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_21"],"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_5":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_12"],"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_6":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_13"],"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_7":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_18"],"pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_0":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_22"],"pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_1":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42"],"pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_2":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41"],"pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_0":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29"],"pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_1":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-pos"],"pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_2":[],"pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_3":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28"],"pin-type-component_336ab846-dec5-4cbf-8759-1d0cae8637dd_0":[],"pin-type-component_336ab846-dec5-4cbf-8759-1d0cae8637dd_1":[],"pin-type-component_33827630-9a86-47d3-b759-b445a42e4930_0":[],"pin-type-component_33827630-9a86-47d3-b759-b445a42e4930_1":[],"pin-type-component_2183a60b-5a7f-4b57-a29c-94c67ecdb107_0":[],"pin-type-component_2183a60b-5a7f-4b57-a29c-94c67ecdb107_1":[],"pin-type-component_b49ac763-faff-4428-8cd2-1f59202c6272_0":[],"pin-type-component_b49ac763-faff-4428-8cd2-1f59202c6272_1":[],"pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_0":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20"],"pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_1":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-pos"],"pin-type-component_96269a28-ca9a-4d81-b0ce-f5da10a7f5a0_0":[],"pin-type-component_96269a28-ca9a-4d81-b0ce-f5da10a7f5a0_1":[],"pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_0":[],"pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_1":[],"pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_2":[]},"pin_to_color":{"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18":"#189AB4","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19":"#7544B1","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20":"#FF0000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20":"#aaaaaa","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25":"#A75740","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28":"#98FF52","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29":"#FF74A3","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32":"#968AE8","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41":"#189AB4","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42":"#FF0000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44":"#189AB4","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45":"#01FFFE","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52":"#189AB4","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53":"#FF0000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55":"#189AB4","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56":"#FF0000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59":"#189AB4","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60":"#95003A","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61":"#005F39","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62":"#000000","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62":"#FF0000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-pos":"#FF0000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-neg":"#189AB4","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-pos":"#FF0000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-neg":"#189AB4","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-pos":"#FF0000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-neg":"#189AB4","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos":"#FF0000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-pos":"#FF0000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-neg":"#189AB4","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-pos":"#FF0000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg":"#189AB4","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos":"#FF0000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-neg":"#189AB4","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61_polarity-neg":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-pos":"#FF0000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-neg":"#189AB4","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62_polarity-pos":"#000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62_polarity-neg":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_0":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_1":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_2":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_3":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4":"#FF0000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5":"#189AB4","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_7":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8":"#91D0CB","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_9":"#007DB5","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_10":"#6A826C","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_11":"#00AE7E","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_12":"#008F9C","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_13":"#5FAD4E","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_14":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_15":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_16":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_17":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_18":"#FF029D","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_19":"#005F39","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_20":"#95003A","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_21":"#C28C9F","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_22":"#683D3B","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_23":"#01FFFE","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_24":"#A75740","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_25":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_26":"#968AE8","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27":"#7544B1","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_28":"#00c7fc","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_29":"#FF937E","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_30":"#000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_31":"#000000","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_0":"#FF0000","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_1":"#005F39","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_2":"#95003A","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_3":"#189AB4","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_0":"#189AB4","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_1":"#FF937E","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_2":"#FF0000","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_0":"#00c7fc","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_1":"#189AB4","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_2":"#FF0000","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_0":"#91D0CB","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_1":"#007DB5","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_2":"#6A826C","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_3":"#00AE7E","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_4":"#C28C9F","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_5":"#008F9C","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_6":"#5FAD4E","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_7":"#FF029D","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_0":"#683D3B","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_1":"#FF0000","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_2":"#189AB4","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_0":"#FF74A3","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_1":"#FF0000","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_2":"#000000","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_3":"#98FF52","pin-type-component_336ab846-dec5-4cbf-8759-1d0cae8637dd_0":"#000000","pin-type-component_336ab846-dec5-4cbf-8759-1d0cae8637dd_1":"#000000","pin-type-component_33827630-9a86-47d3-b759-b445a42e4930_0":"#000000","pin-type-component_33827630-9a86-47d3-b759-b445a42e4930_1":"#000000","pin-type-component_2183a60b-5a7f-4b57-a29c-94c67ecdb107_0":"#000000","pin-type-component_2183a60b-5a7f-4b57-a29c-94c67ecdb107_1":"#000000","pin-type-component_b49ac763-faff-4428-8cd2-1f59202c6272_0":"#000000","pin-type-component_b49ac763-faff-4428-8cd2-1f59202c6272_1":"#000000","pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_0":"#aaaaaa","pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_1":"#FF0000","pin-type-component_96269a28-ca9a-4d81-b0ce-f5da10a7f5a0_0":"#000000","pin-type-component_96269a28-ca9a-4d81-b0ce-f5da10a7f5a0_1":"#000000","pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_0":"#000000","pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_1":"#000000","pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_2":"#000000"},"pin_to_state":{"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62":"neutral","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-neg":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62_polarity-pos":"neutral","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62_polarity-neg":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_0":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_1":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_2":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_3":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_7":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_9":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_10":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_11":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_12":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_13":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_14":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_15":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_16":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_17":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_18":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_19":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_20":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_21":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_22":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_23":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_24":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_25":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_26":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_28":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_29":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_30":"neutral","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_31":"neutral","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_0":"neutral","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_1":"neutral","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_2":"neutral","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_3":"neutral","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_0":"neutral","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_1":"neutral","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_2":"neutral","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_0":"neutral","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_1":"neutral","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_2":"neutral","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_0":"neutral","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_1":"neutral","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_2":"neutral","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_3":"neutral","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_4":"neutral","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_5":"neutral","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_6":"neutral","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_7":"neutral","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_0":"neutral","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_1":"neutral","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_2":"neutral","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_0":"neutral","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_1":"neutral","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_2":"neutral","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_3":"neutral","pin-type-component_336ab846-dec5-4cbf-8759-1d0cae8637dd_0":"neutral","pin-type-component_336ab846-dec5-4cbf-8759-1d0cae8637dd_1":"neutral","pin-type-component_33827630-9a86-47d3-b759-b445a42e4930_0":"neutral","pin-type-component_33827630-9a86-47d3-b759-b445a42e4930_1":"neutral","pin-type-component_2183a60b-5a7f-4b57-a29c-94c67ecdb107_0":"neutral","pin-type-component_2183a60b-5a7f-4b57-a29c-94c67ecdb107_1":"neutral","pin-type-component_b49ac763-faff-4428-8cd2-1f59202c6272_0":"neutral","pin-type-component_b49ac763-faff-4428-8cd2-1f59202c6272_1":"neutral","pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_0":"neutral","pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_1":"neutral","pin-type-component_96269a28-ca9a-4d81-b0ce-f5da10a7f5a0_0":"neutral","pin-type-component_96269a28-ca9a-4d81-b0ce-f5da10a7f5a0_1":"neutral","pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_0":"neutral","pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_1":"neutral","pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_2":"neutral"},"next_color_idx":27,"wires_placed_in_order":[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-pos"],["pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_14","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8"],["pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6","pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_25"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6","pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_22"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_22"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-pos"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-neg"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_0"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_3"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_19","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_20","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_1"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_2"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_2"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_0"],["pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_1","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_29"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_2"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_1"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_28","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_0"],["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_0","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8"],["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_1","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_9"],["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_2","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_10"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_11","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_3"],["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_4","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_21"],["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_5","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_12"],["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_6","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_13"],["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_7","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_18"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_1"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_2"],["pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_0","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_22"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-pos","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_1"],["pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_0","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_26"],["pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_3","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_24"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45"],["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_23","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27"],["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-neg"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20","pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_0"],["pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_1","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-pos"],["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-pos"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg"]]],[[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg"]],[]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-pos"]]],[[],[["pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_14","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8"]]],[[["pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_14","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8"]],[]],[[],[["pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5"]]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6","pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_25"]]],[[["pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_25","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6"]],[]],[[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg"]],[]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg"]]],[[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg"]],[]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6","pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_22"]]],[[["pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_22","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6"]],[]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_22"]]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg"]]],[[["pin-type-breadboard_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_22","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5"]],[]],[[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-pos"]],[]],[[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-power-rail_7f4e5b24-8c91-4743-bac7-b54846f3442c_0_29_polarity-neg"]],[]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-pos"]]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-neg"]]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59"]]],[[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos"]],[]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62"]]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_0"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_3"]]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_19","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61"]]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_20","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_1"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_2"]]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56"]]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55"]]],[[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg"]],[]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_2"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_0"]]],[[],[["pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_1","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_29"]]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53"]]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_2"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_1"]]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_28","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_0"]]],[[],[["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_0","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8"]]],[[],[["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_1","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_9"]]],[[],[["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_2","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_10"]]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_11","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_3"]]],[[],[["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_4","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_21"]]],[[],[["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_5","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_12"]]],[[],[["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_6","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_13"]]],[[],[["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_7","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_18"]]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40"]]],[[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos"]],[]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42"]]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_1"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_2"]]],[[],[["pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_0","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_22"]]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-pos","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_1"]]],[[],[["pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_0","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_26"]]],[[],[["pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_3","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_24"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45"]]],[[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-neg"]],[]],[[],[["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44"]]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_23","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45"]]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27"]],[]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27"]]],[[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27"]],[]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27"]]],[[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27"]],[]],[[],[["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-neg"]]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20","pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_0"]]],[[],[["pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_1","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-pos"]]],[[],[]],[[],[]],[[],[["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-pos"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18":"0000000000000031","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19":"0000000000000030","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20":"0000000000000034","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20":"0000000000000032","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25":"0000000000000027","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28":"0000000000000026","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29":"0000000000000024","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32":"0000000000000025","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41":"0000000000000021","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42":"0000000000000020","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44":"0000000000000028","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45":"0000000000000029","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52":"0000000000000010","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53":"0000000000000009","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55":"0000000000000007","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56":"0000000000000006","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59":"0000000000000003","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60":"0000000000000005","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61":"0000000000000004","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62":"_","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62":"0000000000000002","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_0_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_0_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_1_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_1_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_2_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_2_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_3_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_3_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_4_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_4_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_5_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_5_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_6_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_6_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_7_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_7_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_8_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_8_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_9_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_9_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_10_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_10_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_11_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_11_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_12_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_12_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_13_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_13_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_14_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_14_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_15_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_15_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-pos":"0000000000000033","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_16_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_17_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_17_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-neg":"0000000000000031","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_19_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-pos":"0000000000000034","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_21_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_21_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_22_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_22_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_23_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_23_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_24_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_24_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_25_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_26_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_26_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_27_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_27_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_28_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_29_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_30_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_30_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_31_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_31_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_32_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_33_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_33_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_34_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_34_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_35_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_35_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_36_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_36_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_37_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_37_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_38_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_38_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_39_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_39_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_40_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_40_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_41_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_42_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_43_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_43_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-neg":"0000000000000028","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_44_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_45_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_46_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_46_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_47_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_47_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_48_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_48_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-pos":"0000000000000023","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_49_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-neg":"0000000000000021","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_50_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos":"0000000000000020","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_51_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_52_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-pos":"0000000000000009","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-neg":"0000000000000010","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_54_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_54_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_55_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_56_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_57_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_57_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_58_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_58_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_59_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-pos":"0000000000000006","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg":"0000000000000007","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos":"0000000000000002","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-neg":"0000000000000003","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61_polarity-neg":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-pos":"0000000000000000","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-neg":"0000000000000001","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62_polarity-pos":"_","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62_polarity-neg":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_0":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_1":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_2":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_3":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4":"0000000000000000","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5":"0000000000000001","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_6":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_7":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8":"0000000000000012","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_9":"0000000000000013","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_10":"0000000000000014","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_11":"0000000000000015","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_12":"0000000000000017","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_13":"0000000000000018","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_14":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_15":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_16":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_17":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_18":"0000000000000019","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_19":"0000000000000004","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_20":"0000000000000005","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_21":"0000000000000016","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_22":"0000000000000022","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_23":"0000000000000029","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_24":"0000000000000027","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_25":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_26":"0000000000000025","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27":"0000000000000030","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_28":"0000000000000011","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_29":"0000000000000008","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_30":"_","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_31":"_","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_0":"0000000000000002","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_1":"0000000000000004","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_2":"0000000000000005","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_3":"0000000000000003","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_0":"0000000000000007","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_1":"0000000000000008","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_2":"0000000000000006","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_0":"0000000000000011","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_1":"0000000000000010","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_2":"0000000000000009","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_0":"0000000000000012","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_1":"0000000000000013","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_2":"0000000000000014","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_3":"0000000000000015","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_4":"0000000000000016","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_5":"0000000000000017","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_6":"0000000000000018","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_7":"0000000000000019","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_0":"0000000000000022","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_1":"0000000000000020","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_2":"0000000000000021","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_0":"0000000000000024","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_1":"0000000000000023","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_2":"_","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_3":"0000000000000026","pin-type-component_336ab846-dec5-4cbf-8759-1d0cae8637dd_0":"_","pin-type-component_336ab846-dec5-4cbf-8759-1d0cae8637dd_1":"_","pin-type-component_33827630-9a86-47d3-b759-b445a42e4930_0":"_","pin-type-component_33827630-9a86-47d3-b759-b445a42e4930_1":"_","pin-type-component_2183a60b-5a7f-4b57-a29c-94c67ecdb107_0":"_","pin-type-component_2183a60b-5a7f-4b57-a29c-94c67ecdb107_1":"_","pin-type-component_b49ac763-faff-4428-8cd2-1f59202c6272_0":"_","pin-type-component_b49ac763-faff-4428-8cd2-1f59202c6272_1":"_","pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_0":"0000000000000032","pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_1":"0000000000000033","pin-type-component_96269a28-ca9a-4d81-b0ce-f5da10a7f5a0_0":"_","pin-type-component_96269a28-ca9a-4d81-b0ce-f5da10a7f5a0_1":"_","pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_0":"_","pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_1":"_","pin-type-component_f740428d-a39d-448f-ac5a-24b4e88ade74_2":"_"},"component_id_to_pins":{"27375bda-91ae-44fd-a8b5-a4fede174c00":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"36f0ce75-1dbd-4c59-b727-b45890b5209b":["0","1","2","3"],"b730a454-d8cc-489a-b7a2-ef95453cd4ac":["0","1","2"],"fefd5a80-67a4-4511-8644-deb5b8b182be":["0","1","2"],"f43f5baf-10b5-4113-931c-ffae3f691543":["0","1","2","3","4","5","6","7"],"9a09bf79-7cf3-4d76-9410-f7a4311d8644":["0","1","2"],"d2d6d00d-6536-449d-854e-7729bcc5cce8":["0","1","2","3"],"336ab846-dec5-4cbf-8759-1d0cae8637dd":["0","1"],"33827630-9a86-47d3-b759-b445a42e4930":["0","1"],"2183a60b-5a7f-4b57-a29c-94c67ecdb107":["0","1"],"b49ac763-faff-4428-8cd2-1f59202c6272":["0","1"],"977f2642-028e-48b9-a72a-d1c123fab533":["0","1"],"d332df42-6ca0-4992-9d92-c982e107f43a":[],"96269a28-ca9a-4d81-b0ce-f5da10a7f5a0":["0","1"],"f740428d-a39d-448f-ac5a-24b4e88ade74":["0","1","2"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-pos"],"0000000000000001":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-neg"],"0000000000000002":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_0"],"0000000000000003":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-neg","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_3"],"0000000000000004":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_19","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_1"],"0000000000000005":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_20","pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_2"],"0000000000000006":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-pos","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_2"],"0000000000000007":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg","pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_0"],"0000000000000008":["pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_1","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_29"],"0000000000000009":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-pos","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_2"],"0000000000000010":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-neg","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_1"],"0000000000000011":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_28","pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_0"],"0000000000000012":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_0","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8"],"0000000000000013":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_1","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_9"],"0000000000000014":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_2","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_10"],"0000000000000015":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_11","pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_3"],"0000000000000016":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_4","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_21"],"0000000000000017":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_5","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_12"],"0000000000000018":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_6","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_13"],"0000000000000019":["pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_7","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_18"],"0000000000000020":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_1"],"0000000000000021":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-neg","pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_2"],"0000000000000022":["pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_0","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_22"],"0000000000000023":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-pos","pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_1"],"0000000000000024":["pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_0","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29"],"0000000000000025":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_26"],"0000000000000026":["pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_3","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28"],"0000000000000027":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25","pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_24"],"0000000000000028":["pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-neg","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44"],"0000000000000029":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_23","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45"],"0000000000000030":["pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27","pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19"],"0000000000000031":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-neg"],"0000000000000032":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20","pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_0"],"0000000000000033":["pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_1","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-pos"],"0000000000000034":["pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20","pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-pos"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000009":"Net 9","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000015":"Net 15","0000000000000016":"Net 16","0000000000000017":"Net 17","0000000000000018":"Net 18","0000000000000019":"Net 19","0000000000000020":"Net 20","0000000000000021":"Net 21","0000000000000022":"Net 22","0000000000000023":"Net 23","0000000000000024":"Net 24","0000000000000025":"Net 25","0000000000000026":"Net 26","0000000000000027":"Net 27","0000000000000028":"Net 28","0000000000000029":"Net 29","0000000000000030":"Net 30","0000000000000031":"Net 31","0000000000000032":"Net 32","0000000000000033":"Net 33","0000000000000034":"Net 34"},"all_breadboard_info_list":["7f4e5b24-8c91-4743-bac7-b54846f3442c_30_2_True_835.5_415.5_right","720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_63_2_True_1112.9999999999998_137.9999999999999_right"],"breadboard_info_list":["720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_63_2_True_1112.9999999999998_137.9999999999999_right"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[846.25,237.49999999999997],"typeId":"b269da49-8c00-4ebb-bd25-5859ea0c7cad","componentVersion":9,"instanceId":"27375bda-91ae-44fd-a8b5-a4fede174c00","orientation":"up","circleData":[[827.5,380],[842.5,380],[857.5,380],[872.5,380],[887.5,380],[902.5,380],[917.5,380],[932.5,380],[962.5,380],[977.5,380],[992.5,380],[1007.5,380],[1022.5,380],[1037.5,380],[773.5,94.99999999999997],[788.5,94.99999999999997],[803.5,94.99999999999997],[818.5,94.99999999999997],[833.5,94.99999999999997],[848.5,94.99999999999997],[863.5,94.99999999999997],[878.5,94.99999999999997],[893.5,94.99999999999997],[908.5,94.99999999999997],[932.5,94.99999999999997],[947.5,94.99999999999997],[962.5,94.99999999999997],[977.5,94.99999999999997],[992.5,94.99999999999997],[1007.5,94.99999999999997],[1022.5,94.99999999999997],[1037.5,94.99999999999997]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"5dcc0497-3d62-4b0f-b16d-dee4d9f57e93\",\"explorerHtmlId\":\"5c557c04-3d0a-4a9a-9f82-2c0ff585f5fe\",\"nameHtmlId\":\"301dcc05-61d8-4db3-a87a-5caff13ffe60\",\"nameInputHtmlId\":\"aa21ae00-4acc-4be2-9308-a772e882a14c\",\"explorerChildHtmlId\":\"e9eac437-d09a-4ad2-b3d4-477d85453989\",\"explorerCarrotOpenHtmlId\":\"5561a252-7e8f-4fab-935c-2eb6ee376ff5\",\"explorerCarrotClosedHtmlId\":\"f705d10d-7361-483c-b496-cb0aee82b59a\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"da896fb4-dec9-440b-aaaa-d82c8172ffde\",\"explorerHtmlId\":\"5c9ef1d3-e5a2-4f94-a643-1b690c7e36da\",\"nameHtmlId\":\"265146d2-57dc-44b0-8b02-907c6b9cb73e\",\"nameInputHtmlId\":\"a28b2b8e-e303-4460-bcf8-ee9f5ad64eb4\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"fb620434-0a3b-4d85-8cbf-5456d8fc7292\",\"explorerHtmlId\":\"ee7548ca-22c3-4de5-b9cf-4ba7f5381803\",\"nameHtmlId\":\"9e425e3e-6315-4668-bcae-7aa3e10b47b4\",\"nameInputHtmlId\":\"df075a4b-db03-4fd4-9c1e-6931c7b56501\",\"code\":\"\"},0,","codeLabelPosition":[846.25,79.99999999999994],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"SEN-15569","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"SparkFun","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[477.0136134999999,718.496435],"typeId":"f7a95729-a811-496b-83f5-7789de376adf","componentVersion":2,"instanceId":"36f0ce75-1dbd-4c59-b727-b45890b5209b","orientation":"up","circleData":[[452.5,785],[467.49922449999997,785],[482.49999849999995,784.9953095000001],[497.4984445,784.9937494999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[575.908,1032.5104999999999],"typeId":"8f4dc0af-d812-4c84-aad9-cfeab9e8c28a","componentVersion":1,"instanceId":"b730a454-d8cc-489a-b7a2-ef95453cd4ac","orientation":"up","circleData":[[557.5,1160],[575.4655,1160],[595.951,1160.2400000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[920.921077,999.3420785000004],"typeId":"905c0666-7ddd-4192-a785-7e454e84ab15","componentVersion":1,"instanceId":"fefd5a80-67a4-4511-8644-deb5b8b182be","orientation":"up","circleData":[[902.5,1130],[925,1130],[947.5,1130]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1336.672258,85.18009099999975],"typeId":"4898f56e-60f9-4315-8c2e-83ff52744e63","componentVersion":1,"instanceId":"f43f5baf-10b5-4113-931c-ffae3f691543","orientation":"up","circleData":[[1292.5,305],[1304.021389,305.1630365000001],[1316.4649255000002,305.1630365000001],[1329.1045000000001,304.9239634999999],[1341.7010365,305.50907300000017],[1353.4094635000001,305.50907300000017],[1365.5069635,305.61603650000006],[1377.5697220000002,305.542829]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1133.645833,1057.608683],"typeId":"507015a7-8113-03cb-aee9-f593197b129c","componentVersion":1,"instanceId":"9a09bf79-7cf3-4d76-9410-f7a4311d8644","orientation":"right","circleData":[[1157.5,830.0000000000001],[1138.75,830.0000000000001],[1120,830.0000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1270,910.4750255],"typeId":"01cc3eef-ba83-0e3d-7920-e5931d8f1e12","componentVersion":4,"instanceId":"d2d6d00d-6536-449d-854e-7729bcc5cce8","orientation":"up","circleData":[[1247.5,965],[1262.5,965],[1277.5,965],[1292.5,965]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"220","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[1165,680.0000000000002],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"336ab846-dec5-4cbf-8759-1d0cae8637dd","orientation":"up","circleData":[[1142.5,680.0000000000002],[1187.5,680.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"220","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[1225.0000000000002,680.0000000000002],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"33827630-9a86-47d3-b759-b445a42e4930","orientation":"up","circleData":[[1202.5000000000002,680.0000000000002],[1247.5000000000002,680]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[954.9923994999999,566.9295574999999],"typeId":"773dd385-6643-437a-99c0-a6e92849b80e","componentVersion":2,"instanceId":"2183a60b-5a7f-4b57-a29c-94c67ecdb107","orientation":"down","circleData":[[947.5,545],[961.4211399999999,544.8568969999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[1322.5625005000002,616.7614505000001],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"b49ac763-faff-4428-8cd2-1f59202c6272","orientation":"right","circleData":[[1322.5,560],[1322.5,665]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1476.7518610000004,949.608393499999],"typeId":"3ce813a8-322b-4f90-a9f5-e0d3b4eaeefb","componentVersion":1,"instanceId":"977f2642-028e-48b9-a72a-d1c123fab533","orientation":"left","circleData":[[1547.5,1040],[1536.600442,1040.060618]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"## Components were connected in the order provided below.\n\n**Ultrasonic Sensor (HC-SR04):**\n  - VCC → 5V\n  - GND → GND\n  - TRIG → Pin 12\n  - ECHO → Pin 11\n\n**DHT11 Temperature Sensor:**\n  - VCC → 5V (in the middle if not defined)\n  - GND → GND (or written as \"-\")\n  - DATA → Pin 2 (or written as \"S\")\n\n**IR Sensor:**\n  - VCC → 5V\n  - GND → GND\n  - OUT → Pin 3\n\n**4×4 Keypad:**\n  - Row 1 → A0\n  - Row 2 → A1\n  - Row 3 → A2\n  - Row 4 → A3\n  - Column 1 → Pin 10\n  - Column 2 → A4\n  - Column 3 → A5\n  - Column 4 → Pin 13\n\n**Servo Motor (SG90):**\n  - Red (VCC) → 5V\n  - Brown (GND) → GND\n  - Orange (Signal) → Pin 9\n\n**RGB LED (Common VCC)**\n  - Common Cathode → GND\n  - Red pin → Pin 5 (with 220Ω resistor)\n  - Blue pin → Pin 7 (with 220Ω resistor)\n\n**Buzzer:**\n  - Positive (+) → Pin 8\n  - Negative (-) → GND\n\n**Simple Fan (2-wire with NPN Transistor):**\nRequired Components:\n  - 1x NPN Transistor (2N2222, BC547, or similar)\n  - 1x 1kΩ Resistor\n  - 1x Diode 1N4007 (for protection)\n\nArduino Pin 4 → 1kΩ Resistor → Transistor Base (middle pin)\nTransistor Emitter (left/right pin) → Arduino GND\nTransistor Collector (left/right pin) → Fan GND (-)\nFan VCC (+) → Arduino 5V\nDiode (1N4007): Cathode to Arduino 5V, Anode to Fan GND","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#aaaaaa","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"19","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[2064.4334126412746,472.14364510045516],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"d332df42-6ca0-4992-9d92-c982e107f43a","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"1000","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[1337.5,612.5],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"96269a28-ca9a-4d81-b0ce-f5da10a7f5a0","orientation":"left","circleData":[[1337.5,665],[1337.5,590]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1337.8018270000002,733.3322825],"typeId":"10d13646-c889-4b39-93c7-eebbfe2262dd","componentVersion":1,"instanceId":"f740428d-a39d-448f-ac5a-24b4e88ade74","orientation":"down","circleData":[[1352.5,695],[1337.5,695],[1322.5,695]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-152.72128","left":"333.85321","width":"2076.93494","height":"1467.20987","x":"333.85321","y":"-152.72128"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-pos\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_4\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"887.5000000000_380.0000000000\\\",\\\"887.5000000000_410.0000000000\\\",\\\"677.5000000000_410.0000000000\\\",\\\"677.5000000000_470.0000000000\\\",\\\"692.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-neg\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_5\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_62_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.5000000000_380.0000000000\\\",\\\"902.5000000000_425.0000000000\\\",\\\"670.0000000000_425.0000000000\\\",\\\"670.0000000000_485.0000000000\\\",\\\"692.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62_3\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"692.5000000000_680.0000000000\\\",\\\"670.0000000000_680.0000000000\\\",\\\"670.0000000000_515.0000000000\\\",\\\"715.0000000000_515.0000000000\\\",\\\"715.0000000000_470.0000000000\\\",\\\"707.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62\",\"endPinId\":\"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_62_4\",\"rawEndPinId\":\"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"692.5000000000_695.0000000000\\\",\\\"692.5000000000_702.5000000000\\\",\\\"655.0000000000_702.5000000000\\\",\\\"655.0000000000_852.5000000000\\\",\\\"452.5000000000_852.5000000000\\\",\\\"452.5000000000_785.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59_3\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_61_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"737.5000000000_680.0000000000\\\",\\\"730.0000000000_680.0000000000\\\",\\\"730.0000000000_612.5000000000\\\",\\\"700.0000000000_612.5000000000\\\",\\\"700.0000000000_485.0000000000\\\",\\\"707.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59\",\"endPinId\":\"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_3\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_59_4\",\"rawEndPinId\":\"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"737.5000000000_695.0000000000\\\",\\\"737.5000000000_717.5000000000\\\",\\\"677.5000000000_717.5000000000\\\",\\\"677.5000000000_807.5000000000\\\",\\\"497.4984445000_807.5000000000\\\",\\\"497.4984445000_784.9937495000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61\",\"endPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_19\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61_3\",\"rawEndPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_19\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"707.5000000000_680.0000000000\\\",\\\"700.0000000000_680.0000000000\\\",\\\"700.0000000000_627.5000000000\\\",\\\"317.5000000000_627.5000000000\\\",\\\"317.5000000000_65.0000000000\\\",\\\"848.5000000000_65.0000000000\\\",\\\"848.5000000000_95.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61\",\"endPinId\":\"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_61_4\",\"rawEndPinId\":\"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"707.5000000000_695.0000000000\\\",\\\"707.5000000000_710.0000000000\\\",\\\"670.0000000000_710.0000000000\\\",\\\"670.0000000000_837.5000000000\\\",\\\"467.4992245000_837.5000000000\\\",\\\"467.4992245000_785.0000000000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60\",\"endPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_20\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60_3\",\"rawEndPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_20\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"722.5000000000_680.0000000000\\\",\\\"722.5000000000_687.5000000000\\\",\\\"655.0000000000_687.5000000000\\\",\\\"655.0000000000_642.5000000000\\\",\\\"295.0000000000_642.5000000000\\\",\\\"295.0000000000_50.0000000000\\\",\\\"863.5000000000_50.0000000000\\\",\\\"863.5000000000_95.0000000000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60\",\"endPinId\":\"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_60_4\",\"rawEndPinId\":\"pin-type-component_36f0ce75-1dbd-4c59-b727-b45890b5209b_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"722.5000000000_695.0000000000\\\",\\\"715.0000000000_695.0000000000\\\",\\\"715.0000000000_822.5000000000\\\",\\\"482.4999985000_822.5000000000\\\",\\\"482.4999985000_784.9953095000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56_2\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"782.5000000000_560.0000000000\\\",\\\"775.0000000000_560.0000000000\\\",\\\"775.0000000000_515.0000000000\\\",\\\"730.0000000000_515.0000000000\\\",\\\"730.0000000000_470.0000000000\\\",\\\"722.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56\",\"endPinId\":\"pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_56_3\",\"rawEndPinId\":\"pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"782.5000000000_575.0000000000\\\",\\\"775.0000000000_575.0000000000\\\",\\\"775.0000000000_1205.0000000000\\\",\\\"595.9510000000_1205.0000000000\\\",\\\"595.9510000000_1160.2400000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55_2\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_60_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_560.0000000000\\\",\\\"790.0000000000_560.0000000000\\\",\\\"790.0000000000_500.0000000000\\\",\\\"722.5000000000_500.0000000000\\\",\\\"722.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55\",\"endPinId\":\"pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_55_3\",\"rawEndPinId\":\"pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_575.0000000000\\\",\\\"790.0000000000_575.0000000000\\\",\\\"790.0000000000_1227.5000000000\\\",\\\"557.5000000000_1227.5000000000\\\",\\\"557.5000000000_1160.0000000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_29\",\"endPinId\":\"pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_1\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_29\",\"rawEndPinId\":\"pin-type-component_b730a454-d8cc-489a-b7a2-ef95453cd4ac_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1007.5000000000_95.0000000000\\\",\\\"1007.5000000000_20.0000000000\\\",\\\"272.5000000000_20.0000000000\\\",\\\"272.5000000000_1205.0000000000\\\",\\\"575.4655000000_1205.0000000000\\\",\\\"575.4655000000_1160.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53_3\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"827.5000000000_680.0000000000\\\",\\\"820.0000000000_680.0000000000\\\",\\\"820.0000000000_470.0000000000\\\",\\\"827.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53\",\"endPinId\":\"pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_53_4\",\"rawEndPinId\":\"pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"827.5000000000_695.0000000000\\\",\\\"820.0000000000_695.0000000000\\\",\\\"820.0000000000_1197.5000000000\\\",\\\"947.5000000000_1197.5000000000\\\",\\\"947.5000000000_1130.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52_3\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_53_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_680.0000000000\\\",\\\"835.0000000000_680.0000000000\\\",\\\"835.0000000000_485.0000000000\\\",\\\"827.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52\",\"endPinId\":\"pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_52_4\",\"rawEndPinId\":\"pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_695.0000000000\\\",\\\"835.0000000000_695.0000000000\\\",\\\"835.0000000000_1182.5000000000\\\",\\\"925.0000000000_1182.5000000000\\\",\\\"925.0000000000_1130.0000000000\\\"]}\"}","{\"color\":\"#00c7fc\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_28\",\"endPinId\":\"pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_0\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_28\",\"rawEndPinId\":\"pin-type-component_fefd5a80-67a4-4511-8644-deb5b8b182be_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5000000000_95.0000000000\\\",\\\"992.5000000000_5.0000000000\\\",\\\"250.0000000000_5.0000000000\\\",\\\"250.0000000000_1242.5000000000\\\",\\\"902.5000000000_1242.5000000000\\\",\\\"902.5000000000_1130.0000000000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8\",\"endPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_0\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_8\",\"rawEndPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"962.5000000000_380.0000000000\\\",\\\"947.5000000000_380.0000000000\\\",\\\"947.5000000000_312.5000000000\\\",\\\"1292.5000000000_312.5000000000\\\",\\\"1292.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_9\",\"endPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_1\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_9\",\"rawEndPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"977.5000000000_380.0000000000\\\",\\\"970.0000000000_380.0000000000\\\",\\\"970.0000000000_320.0000000000\\\",\\\"1304.0213890000_320.0000000000\\\",\\\"1304.0213890000_305.1630365000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_10\",\"endPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_2\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_10\",\"rawEndPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5000000000_380.0000000000\\\",\\\"985.0000000000_380.0000000000\\\",\\\"985.0000000000_327.5000000000\\\",\\\"1316.4649255000_327.5000000000\\\",\\\"1316.4649255000_305.1630365000\\\"]}\"}","{\"color\":\"#00AE7E\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_11\",\"endPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_3\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_11\",\"rawEndPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1007.5000000000_380.0000000000\\\",\\\"1000.0000000000_380.0000000000\\\",\\\"1000.0000000000_335.0000000000\\\",\\\"1329.1045000000_335.0000000000\\\",\\\"1329.1045000000_304.9239635000\\\"]}\"}","{\"color\":\"#C28C9F\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_21\",\"endPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_4\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_21\",\"rawEndPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"878.5000000000_95.0000000000\\\",\\\"878.5000000000_-152.5000000000\\\",\\\"1502.5000000000_-152.5000000000\\\",\\\"1502.5000000000_335.0000000000\\\",\\\"1341.7010365000_335.0000000000\\\",\\\"1341.7010365000_305.5090730000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_12\",\"endPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_5\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_12\",\"rawEndPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_380.0000000000\\\",\\\"1022.5000000000_417.5000000000\\\",\\\"1353.4094635000_417.5000000000\\\",\\\"1353.4094635000_305.5090730000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_13\",\"endPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_6\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_13\",\"rawEndPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1037.5000000000_380.0000000000\\\",\\\"1037.5000000000_402.5000000000\\\",\\\"1365.5069635000_402.5000000000\\\",\\\"1365.5069635000_305.6160365000\\\"]}\"}","{\"color\":\"#FF029D\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_18\",\"endPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_7\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_18\",\"rawEndPinId\":\"pin-type-component_f43f5baf-10b5-4113-931c-ffae3f691543_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"833.5000000000_95.0000000000\\\",\\\"833.5000000000_-182.5000000000\\\",\\\"1525.0000000000_-182.5000000000\\\",\\\"1525.0000000000_320.0000000000\\\",\\\"1377.5697220000_320.0000000000\\\",\\\"1377.5697220000_305.5428290000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42_3\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_51_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5000000000_680.0000000000\\\",\\\"992.5000000000_672.5000000000\\\",\\\"850.0000000000_672.5000000000\\\",\\\"850.0000000000_470.0000000000\\\",\\\"857.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42\",\"endPinId\":\"pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_42_4\",\"rawEndPinId\":\"pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5000000000_695.0000000000\\\",\\\"992.5000000000_800.0000000000\\\",\\\"1138.7500000000_800.0000000000\\\",\\\"1138.7500000000_830.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41_3\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_50_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1007.5000000000_680.0000000000\\\",\\\"1007.5000000000_657.5000000000\\\",\\\"865.0000000000_657.5000000000\\\",\\\"865.0000000000_485.0000000000\\\",\\\"872.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41\",\"endPinId\":\"pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_41_4\",\"rawEndPinId\":\"pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1007.5000000000_695.0000000000\\\",\\\"1000.0000000000_695.0000000000\\\",\\\"1000.0000000000_785.0000000000\\\",\\\"1120.0000000000_785.0000000000\\\",\\\"1120.0000000000_830.0000000000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_22\",\"endPinId\":\"pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_0\",\"rawStartPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_22\",\"rawEndPinId\":\"pin-type-component_9a09bf79-7cf3-4d76-9410-f7a4311d8644_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"893.5000000000_95.0000000000\\\",\\\"893.5000000000_-205.0000000000\\\",\\\"1690.0000000000_-205.0000000000\\\",\\\"1690.0000000000_815.0000000000\\\",\\\"1157.5000000000_815.0000000000\\\",\\\"1157.5000000000_830.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_1\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-pos\",\"rawStartPinId\":\"pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_1\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_49_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_965.0000000000\\\",\\\"1262.5000000000_1010.0000000000\\\",\\\"1180.0000000000_1010.0000000000\\\",\\\"1180.0000000000_710.0000000000\\\",\\\"1015.0000000000_710.0000000000\\\",\\\"1015.0000000000_620.0000000000\\\",\\\"895.0000000000_620.0000000000\\\",\\\"895.0000000000_470.0000000000\\\",\\\"887.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29\",\"endPinId\":\"pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_29_4\",\"rawEndPinId\":\"pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1187.5000000000_695.0000000000\\\",\\\"1195.0000000000_695.0000000000\\\",\\\"1195.0000000000_980.0000000000\\\",\\\"1247.5000000000_980.0000000000\\\",\\\"1247.5000000000_965.0000000000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32\",\"endPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_26\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_32_2\",\"rawEndPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_26\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5000000000_665.0000000000\\\",\\\"1135.0000000000_665.0000000000\\\",\\\"1135.0000000000_50.0000000000\\\",\\\"962.5000000000_50.0000000000\\\",\\\"962.5000000000_95.0000000000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28\",\"endPinId\":\"pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_3\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_28_4\",\"rawEndPinId\":\"pin-type-component_d2d6d00d-6536-449d-854e-7729bcc5cce8_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1202.5000000000_695.0000000000\\\",\\\"1210.0000000000_695.0000000000\\\",\\\"1210.0000000000_995.0000000000\\\",\\\"1292.5000000000_995.0000000000\\\",\\\"1292.5000000000_965.0000000000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25\",\"endPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_24\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_25_2\",\"rawEndPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_24\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1247.5000000000_665.0000000000\\\",\\\"1247.5000000000_657.5000000000\\\",\\\"1157.5000000000_657.5000000000\\\",\\\"1157.5000000000_35.0000000000\\\",\\\"932.5000000000_35.0000000000\\\",\\\"932.5000000000_95.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_0\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_44_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"962.5000000000_530.0000000000\\\",\\\"970.0000000000_530.0000000000\\\",\\\"970.0000000000_485.0000000000\\\",\\\"962.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45\",\"endPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_23\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_45_0\",\"rawEndPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_23\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"947.5000000000_530.0000000000\\\",\\\"940.0000000000_530.0000000000\\\",\\\"940.0000000000_447.5000000000\\\",\\\"1120.0000000000_447.5000000000\\\",\\\"1120.0000000000_65.0000000000\\\",\\\"908.5000000000_65.0000000000\\\",\\\"908.5000000000_95.0000000000\\\"]}\"}","{\"color\":\"#7544B1\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19\",\"endPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_19_3\",\"rawEndPinId\":\"pin-type-component_27375bda-91ae-44fd-a8b5-a4fede174c00_27\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1337.5000000000_575.0000000000\\\",\\\"1337.5000000000_567.5000000000\\\",\\\"1180.0000000000_567.5000000000\\\",\\\"1180.0000000000_140.0000000000\\\",\\\"985.0000000000_140.0000000000\\\",\\\"985.0000000000_95.0000000000\\\",\\\"977.5000000000_95.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_18_3\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_18_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1352.5000000000_680.0000000000\\\",\\\"1360.0000000000_680.0000000000\\\",\\\"1360.0000000000_485.0000000000\\\",\\\"1352.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#aaaaaa\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20\",\"endPinId\":\"pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_1_20_3\",\"rawEndPinId\":\"pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1322.5000000000_680.0000000000\\\",\\\"1315.0000000000_680.0000000000\\\",\\\"1315.0000000000_1100.0000000000\\\",\\\"1547.5000000000_1100.0000000000\\\",\\\"1547.5000000000_1040.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_1\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-pos\",\"rawStartPinId\":\"pin-type-component_977f2642-028e-48b9-a72a-d1c123fab533_1\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_16_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1536.6004420000_1040.0606180000\\\",\\\"1536.6004420000_1085.0000000000\\\",\\\"1667.5000000000_1085.0000000000\\\",\\\"1667.5000000000_440.0000000000\\\",\\\"1382.5000000000_440.0000000000\\\",\\\"1382.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20\",\"endPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_1\",\"rawEndPinId\":\"pin-type-power-rail_720e8feb-7c9f-4b8c-bf81-569d7ef1c5bd_0_20_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1322.5000000000_545.0000000000\\\",\\\"1322.5000000000_470.0000000000\\\"]}\"}"],"projectDescription":""}PK
     $s�[               jsons/PK
     $s�[����H  �H     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino UNO","category":["User Defined"],"userDefined":true,"id":"b269da49-8c00-4ebb-bd25-5859ea0c7cad","subtypeDescription":"","subtypePic":"e30496d1-6e1c-40fa-a66f-2add70ecdc94.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"a7fde0f7-2836-4f0c-aad0-66dcccec46ff.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":9,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"HC-SR04 Ultrasonic Sensor","category":["User Defined"],"userDefined":true,"id":"f7a95729-a811-496b-83f5-7789de376adf","subtypeDescription":"","subtypePic":"5a738b76-89aa-4728-b8e5-f09c859dbb14.png","pinInfo":{"numDisplayCols":"17.75472","numDisplayRows":"9.29339","pins":[{"uniquePinIdString":"0","positionMil":"724.31191,21.31240","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"824.30674,21.31240","isAnchorPin":false,"label":"TRIG"},{"uniquePinIdString":"2","positionMil":"924.31190,21.34367","isAnchorPin":false,"label":"ECHO"},{"uniquePinIdString":"3","positionMil":"1024.30154,21.35407","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"SEN-15569","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"SparkFun","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"ba153158-cccd-4fb1-9320-38bebad1b7f9.png","componentVersion":2,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"DHT11 Sensor Module","category":["User Defined"],"id":"8f4dc0af-d812-4c84-aad9-cfeab9e8c28a","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"fd2cb464-8539-444d-bb0b-3750bec3ea07.png","iconPic":"3024baee-4b71-48cf-83e2-7da05d24f50a.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.00000","numDisplayRows":"20.00000","pins":[{"uniquePinIdString":"0","positionMil":"377.28000,150.07000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"497.05000,150.07000","isAnchorPin":false,"label":"Data"},{"uniquePinIdString":"2","positionMil":"633.62000,148.47000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"ir sensor ","category":["User Defined"],"id":"905c0666-7ddd-4192-a785-7e454e84ab15","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"8f771a2d-db90-4bfd-8b3e-8d66edcda07a.png","iconPic":"0c7fd013-2f4e-47d0-a46e-2d19cc1fd6f6.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"18.65672","pins":[{"uniquePinIdString":"0","positionMil":"210.52632,61.78319","isAnchorPin":true,"label":"out"},{"uniquePinIdString":"1","positionMil":"360.52632,61.78319","isAnchorPin":false,"label":"gnd"},{"uniquePinIdString":"2","positionMil":"510.52632,61.78319","isAnchorPin":false,"label":"vcc"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"4x4 Keypad","category":["User Defined"],"id":"4898f56e-60f9-4315-8c2e-83ff52744e63","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"bf314729-9196-4b76-b154-4ab11fec66f9.png","iconPic":"a88da2ca-7e0d-495e-a5bf-cdc1eeca5e78.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"17.20701","numDisplayRows":"30.38685","pins":[{"uniquePinIdString":"0","positionMil":"565.86878,53.87644","isAnchorPin":true,"label":"R0"},{"uniquePinIdString":"1","positionMil":"642.67804,52.78953","isAnchorPin":false,"label":"R1"},{"uniquePinIdString":"2","positionMil":"725.63495,52.78953","isAnchorPin":false,"label":"R2"},{"uniquePinIdString":"3","positionMil":"809.89878,54.38335","isAnchorPin":false,"label":"R3"},{"uniquePinIdString":"4","positionMil":"893.87569,50.48262","isAnchorPin":false,"label":"C0"},{"uniquePinIdString":"5","positionMil":"971.93187,50.48262","isAnchorPin":false,"label":"C1"},{"uniquePinIdString":"6","positionMil":"1052.58187,49.76953","isAnchorPin":false,"label":"C2"},{"uniquePinIdString":"7","positionMil":"1133.00026,50.25758","isAnchorPin":false,"label":"C3"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Tower Pro SG90 servo","category":["Output"],"userDefined":true,"id":"507015a7-8113-03cb-aee9-f593197b129c","subtypeDescription":"","subtypePic":"879f6d20-9391-47d7-8a0d-9140b0e14aa9.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"32.91732","numDisplayRows":"12.50000","pins":[{"uniquePinIdString":"0","positionMil":"128.47478,784.02778","isAnchorPin":true,"label":"Signal"},{"uniquePinIdString":"1","positionMil":"128.47478,659.02778","isAnchorPin":false,"label":"+5V"},{"uniquePinIdString":"2","positionMil":"128.47478,534.02778","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"iconPic":"c5725ab6-c6f4-4984-98e2-b9c0e10adf5a.png","componentVersion":1,"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"RGB Light (Common Cathode)","category":["User Defined"],"userDefined":true,"id":"01cc3eef-ba83-0e3d-7920-e5931d8f1e12","subtypeDescription":"","subtypePic":"4a8a1475-7a47-485c-913d-9939fe0b1f0f.png","iconPic":"3357ace3-f4e2-44e5-8366-d3a4568261a9.png","imageLocation":"local_cache","componentVersion":4,"pinInfo":{"numDisplayCols":"3.30000","numDisplayRows":"7.58333","pins":[{"uniquePinIdString":"0","positionMil":"15.00000,15.66667","isAnchorPin":true,"label":"R"},{"uniquePinIdString":"1","positionMil":"115.00000,15.66667","isAnchorPin":false,"label":"G"},{"uniquePinIdString":"2","positionMil":"215.00000,15.66667","isAnchorPin":false,"label":"B"},{"uniquePinIdString":"3","positionMil":"315.00000,15.66667","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/acf95281-a80d-4c2c-84ba-9b0b6c51a552.svg","propertiesV2":[]},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Buzzer","category":["User Defined"],"id":"773dd385-6643-437a-99c0-a6e92849b80e","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"f093df24-6efd-4d47-a863-17c5645b3aaa.png","iconPic":"72f663bc-d85e-4d27-9085-2f4219a623d3.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.39400","numDisplayRows":"9.39400","pins":[{"uniquePinIdString":"0","positionMil":"369.64933,323.50295","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"276.84173,322.54893","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Fan","category":["User Defined"],"userDefined":true,"id":"3ce813a8-322b-4f90-a9f5-e0d3b4eaeefb","subtypeDescription":"","subtypePic":"9ce856c6-be81-4769-87b3-53be9928d02a.png","iconPic":"627fe4d2-0152-4b97-938d-4b9176d7a483.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"12.40259","numDisplayRows":"10.33548","pins":[{"uniquePinIdString":"0","positionMil":"17.51879,45.11974","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"17.11467,117.78346","isAnchorPin":false,"label":"5V"}],"pinType":"wired"},"properties":[],"componentVersion":1,"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":" A3144 Magnetic Hall Effect Sensor","category":["User Defined"],"id":"10d13646-c889-4b39-93c7-eebbfe2262dd","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6a97e33c-aa93-4e7b-a2bd-349ce97096b8.png","iconPic":"e65d6d59-bd1f-4659-a32c-fe6c1b0070ef.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"2.74401","numDisplayRows":"6.03012","pins":[{"uniquePinIdString":"0","positionMil":"39.21268,45.95745","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"139.21268,45.95745","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"239.21268,45.95745","isAnchorPin":false,"label":"OUT"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     $s�[               images/PK
     $s�[�R�W�  W�  /   images/e30496d1-6e1c-40fa-a66f-2add70ecdc94.png�PNG

   IHDR  u  v   ��:   	pHYs  �  ��+  �	IDATx��	�ם�����w�}!��l��Zhz��@?aK3�`l���-Ü1���vws�c�w������=��-,��lt��#��%K��� �ElE-Ԟ9�ݪ�����̈��ܾ�9A%��q#n�ȼ_��"!�fs]uD��$�\B�0$R+�B!��� &�t���4H�BQ�&�뿿6�m��#�B!$71��_�yd�䪰��s˚�u5��NC��-�B!���&��E��]S($7	!�B!$/�UaGQ� �7玕�%�7��t����˒i�(���F��C��B!�B��EaGQ��u[7a�����������!y�ђiF�����!�B!�&ׄE��l��emM��8If��?�J���2)K��̙3�ih�kB!�B�p䒰��s@u$��X^e�������r!�B!�&W�E�A� yD!�B!Ğ\vu`�KB!�B
�lvu)R���B!�B)H�Y�Q�R �b�4I(z4����±ȼP(6Mb���hB!���d������gL�ۧ���ή��^7n�DB}���'�;"��|���)*�Hqq��_����}�Cr%�$���';e��a6m�/J�l�V�,7D�Z�Kk�B!��Ad����������'��s/^��󘢢"Yq�d���������_:}2�D�\_(����uMN?۵u��.�-��-��77�B�w�B!��6aGQGH����6�>�-^���u��f�Κ"%�ֈ�,����3�z�����v�.��]�X���vٮ���@6	;�:B�XL��D�~w�>Ow�u]s��ڪG67�%�h|y9��1���2���ns����,��v�.�e�fڪG�G��)�R�zA��pϰ��S��]��o���ϧ��lvu��8t-}х�İqsi���u;+ݼ�(nr#�!�B�lvu��0qA��?A���B!d(�vu��(���˥�:+vU�ln�H�gB!�B�@�2�6E!9JT|��K�b�<�uk:�S����̮(U���]��v�n�+�Ѩ���z��P($�)��a�l���n.@QG�����S���������:P^^������%_n�leڞX�3S��F7��ܺa����tww�},��%2r���8d�l��]/���������%W�^M{_�pXƎ���e�l���n.@QG���z�����ܬD��Ç���9������v�T��0A*jj���Zjkk��#���m��l]�[�ym(~����EZZ�?&ҙ�ab6v�X�%����]��v����D"ERQQ�քTODQw5��(�e�l7�vs�� ����Ւ
��w�Tg��@̝?^.�=+'�~[�����bn�!�ʌ�!��%1��?�=��5^�?�W�1y�x]>n�T]3C��~���4IF��D^&�(��yw����\����Q$<�ǁ:v5�lݒNҔt&hzb�/xL��.�e�l��v�"�	�y"�v�.���l&�Άx�\B̝<|X>nj��C��Q#��j���s����i@��a)���R,��v� o��5)�6M�/�s�6w��3&���Hn�h(�(�C��Y����<1c�l��ݠ��
7R/&�l����t �Έ�n��s{�Jǁ�2�s��e�q�t:��]�q�`�.�H穓����rd�T��?�/2�����^�3���J$K�G���D��>Jy�Oz�'3��v�.����^�p!���k��Γ�(�e�l7?�O~�qŕ+W佷ޒ#��i55Rk��+��K�"�G�ʸ��"i;}J�ܺE.�志ًɄ	�8 &M�E �f�#[�xQ���=�'m^�M�]��v�n����J����a�l���uDA���.W^��\?�^�;&}==��qWq�ʱ�~"��2e�!�a�I/a�͐�#�B!$#P�%�~�{�D��'�*�����(~ �$Y_V&�엽O=%���i�K�h8�$Y�f���B!$cP�8����C`���ʩS��[Ɉ�"�|��4��?ɟ��*��B!����Y.�񆴿�[�PV*�t-�.��7������+�ň$��7��/a=K��B!�d��Y.O��_�5u�r���(nP®�Hξ���;�]'�.^���B!�BR���@���;;��Z���C�
���YR"o�h�L�9S&N�*Ğ�"��.ٕ3/�pB!���AQW����_K�'�'��Ύ����G�R��.����e��մ�B!��"uHgg�m�\S[#�?�P��;�,���W_�O�/�q�&	���e��θt�B!�d������Rc���u��Rˈ����K�2��P!Y(�B!$cP��?u�|~�ti��J���Q5���"= hj��UUr��i�&`�+�D�Hӯ������L��,P�n��J��3fL���W�]��v�n����K�������]��E�fu2��J���P���}\\/;O������ ӥ�v���r���y�g��4!�ڪG6/o�޺��E�^�g���r�5�8�L{{�tu%@�v�.�e�^���\.X���gp�8��v�nf��F(�
���pD:._�l�(Vֺ�R�% SB*+D�AC�;�Ĭ�������6�4��v�.��8��c�:�\ii���vB�v�.�M��l�����x��T��I˙3���6�غO��!��BrO��Ӻ��;���^����t��vb����g\�.�e�l�i�^�v"�q;!e�l���n6CQW`t��H��2^�`8"�R�t�!�)���$��uk6ׅB�-n?�DdĈiM�4�b��b)�5�]��vٮ�v�"�,�iND5zB��ő�]��~�� E]��z�Ttg���7l�E�p]tw&c�j��ӱ�Iww�\�xѓ����]��v�h�+P����]��v�����("��^�v`�#��pcţ�^��}A�1i\�5��#���Yа]��v�n������]��v�:BrXʊ��f�Bٺ�9�6Q� 5�$�B!YE]�Q\��<LK]J�BrSM$������+����M�B!�B�%7f����ha�����\1�r	!�BH�AQW`�"ER\^.�L�:MuN����z��7�>�5�Y)��fs�@R�1tg&�T�p,�u�|��X�j��t`�l��]?h�%o���n��׋�]����+0FL�,��[q�X_�d#�XLjg��X�B����[����ۿ��)���:t!%覊ϼxe�d��v�.��/�z�]����f#uF̈́	r�w���L����b�!���O��;(��q�JL���}�3�x;5/�D��pmb�B!��E]�1a�l��g�IyMMV�:�>c�<w���I���"y*��&	E�FCrԼ]8�g��i��p����B!$7�����m���Ei�L^�{��U��kJ++���LF������6 �:�1�~�mB�C	<cQ�톼9 �Ƙ2Kgϐ9F�׻���!�BH�������jI���U����<o�Mz����/۬u=��9g���ds&���|Ff:���[�çdE�.�ґ��M����>-�&��i#���xE���D_?(�9x>�BH!BQW�\w���jӯ�v�Ȭutݱ�|�s�B����R���2�<�z�{fLTbo�S�$W�3�g�ßW�BN8��M���E�e��?S�B!�E]+��[�T"}�Uֺ�hTb�2��[��lc��k	���n����D�]r�52��F�_j�\ �®�!;��h�{v�.P�,��}�8�K�I�/��Vgg�kt�⵪���l�

����%K�x]F�-��@�A��Jw���BH62e�k�@�-���z�{��qawǌ��#D,q�"��Ϥ�CއuNY�6|Y�ϽV���wBH*`+���&�1���
� ���P�6[�*ʔ�0�	��xcz�O^�J˳>�-/�����KnW}��e�p�X�q�k������~5h}���Xi��l|�ׁ=PjZ�����X~�l|��� ���E���1�����u_f�3����(�
X����"���[R9r��_t^��+����z捴����,%]W��Gwi�|0sQ��6��(ǧޜ��%�W��^�p4�z�N�M���G�NT�~�0yHֶ��m��#)�]z��������k�'��k=Ld1�����'�j�j�O���H��bw�R��8�lu)Ʊ�_^?ŗɽ�O ��O��BM|�=����^-00&������t�w='ZLڡ�����n1���O��y|��ϸ/���>�p6�86W&~��@���-R�~��v����𙄢����t�����d����~Uz:;?�]�4]W8"��o�F��:���v�o�-�zE��ًmw䅣�o*�n���������u���B�_k�>��>�)�ښɤг��W���	��ǰ�a��ɒ�Ƹ�$�1�!��ˣ���6_�E�_YA,�Řઉ��>�q�jf���)�t��z��p]О��Ax��%���7=̖;e�B�|?yٓv��8�����x�u�/�PlZ��|�=��z|zu��f��M7��3����7c	�m���~�}�o,)�
�������o�������Gv}}�J�����/}�+a���Rv^�����RЙ���Ϟ��o��ՙ�x��#i��%z�ݐ�A���uB[i�� �u�fr�uz��, �yjV'c�z�����gF	��L�1m0�_Y��0��x鎨,9F��1��A�d��m��7�S��w�����ǈ�hA����B���ĸW���Ό���z}���8?�+������1lN��7�74������񷖢������kk�7��]�0i�\9y*0a��^����ZXi�	;��N��!�4��������M�T� ����g_2<tC
�̮ts���~���νmZ}� k!���D�ڮ~�~0�����X�(7[���t�u7��>��
��ۆ��n�����z��A�,fk�c|`���S�l�����_��,�;�/�+�)T���3��H���.�ʊ�"��%6���#2j�t�w_T	���������ꀅ�S_]-��Y|I���&���];a秠ӄ� +�<*s�ޗ�����Dx�Y�nH���VgGܽ�C�:e�o��,c⌶!�!Lp]1��>�߫k�����/�ԡ-sL�H��7Zܩ{��)����DL�7������G�[Q�^N�16�����\@�v1Np~]/|��G�Xt�N�PI_�v���9�c:p�xy��ݍƘ�k��J������Qň��kE?$Ľ�,ۖ�E}}���7(��n�?l����q;e�\�xї�)���t�E�/���~#-t>ⷰ�X�]P횅]�����?��>$O	
L�Ryr�I�����ܐ *%f��ۧvGN���ަ�_b���ya�:L�0q�rB�bhD�.�ؿ)_Z2H8@X��DN]+�
�Mu �cU�K��Ճ��X�u��	�����"���@�^�D?\~=��y@ kwD�}���xy�hGd�wf/���OQ�Ǹ�A�-��a��Ȭ�V{�Pԑ8�c�Ȣ��[�����+R?m���?�I���tG���Iф�x�7T{��m2a�A[�~]�� ۅ��-*����t�vOO�1��(k�%p�n���S�$;h
�IM�&A��K�i�x=�18`��dj�O.Ov�Ƥ�j��Ѽy_&&���t	
s������o.��N��^�� ��NFa��^6m���!~��g��D��8�y����>��I��'�;�vPI��3u�Eb��X�ZN<(��~Jjjk�j�h��N��h,&��R���J����	�t��!�ۓ�v+�.*���%�,(7@��p���+AYhnHzb��?0Q�F�vu�3��`"�[��,�WɅI�~=Â3���A��*�@z�D����&���_�gɚl���������	���w��_���Dj��$�"ᆸ�2�X��D.��=��9����ɍ���#�D&k��5%Yjo�5�y:���2i��㔂�쎘�:k׻�y�,�B
�� �{��}�8i�Ln�YW+������w�?.��|"��쑳o�!��=RZ^.��s��q=Ʊ����װʕ�+�fϑk?�X��e�HD�r�t�K��8���}pD޾|�>���rdu1�KL�G�:����x=�/D7$�~aԓc�V��l��˥�BH栨�������'��/")ӢN���y��+r��u��Yi�l�7WTT$+n�,��1VUU%����y+��g���d�	��KW���.9�Ijc6�v��,���fx�r��nHΞk��v��Ep�q>p9��h��=�p�U�.�[
��5�t�h?\�
�)��_I6�1g�h��ٕV�F,����������,�q2����:�f��m�GTIEE�||�^�@е�uH4���Z�(�ힱo�V��mF��Ew.��+���Kn�O;�a-,R�<~�]�`�D9x��,���\�e0��ص�����$;�|��6m�<����E!��1#�K������ܦ���H�(l�;8وj�V��n������2�&d*�?��]3�^|CV�5O��x�lX|�<���B����`\��w�,���������8Yy�Lyp�̂'��oճ/I!pǌI�/Ɠ�u]�`b��{���d��7��|����g��9���A�B���ۭ�����B��v�]� qn�Ə���L��g��>,���55�"�&����Sn��+WL=N �
a���)#j��X¢Y������T�>&�:B!y���a�T�L��g�������d�xϝ_�B'�t��fA�?����X�w<�$���[��:B)0�����<����i͸��g��up3��E�aJ}���z��#��{���8)�����վ��½u��I�u���JQG!�NL���7('T�s;2����	q��!$�8p���\aÀU%(��q�J���B�/`��=a��{_�s��:x�s7Ld����e�=w%�,`��G(�)p.\h�ʲ�5��L-m���nSK̻vۤ�|p��)˥��5/�5똝�J�������������l7V��o�ض�m!�b� �N\nl�[h�P����Ҋ_n��]6{��8[���<NNCQGH��'����G"��_���M���;���.�]p>9�*�	^���t�ty�ݏ���L�k��-�J���khX���E'�@E���g�(�qR(�k�vi�O7�U?~I��_1��.��HP�ȏ��H~}�tt'/��S�ejU�oA��G_> �p�X�I�?u�W�[%�X,�p�k�����O����n_��n$q�ӧ���{떑�v�G�{��A`��(~nqY(q@�SP`]̚�GOv�"�]��B'�~���.���e�/���3��.5ur�r�ZR�����b!��F�3�BD���	����3����v���ue��'!��������/b�T�������?�ӌ��N��iWM�{l{u��B1���R��Iv�/\+\�c�z����B'H�s���Źٹ?��+�cϿ��1������E!�d *X�t����)�����+��%���.7�p�l�_s{:���맨���8b`�we�1a����@d {��	������+�qR(�q�K7$�5?)!g���B2�v}��!������z�WE��K��@�!^.YLl�v�|!���ڤ*��Z�nj�6N
�|���u�P�BH�����
��Ec�K&�����VAa�6��a�öX�0%=��b�L������m��84\�$�������)))�p
	C���3�t�d-���\O������:gwV�"R�9
���2�&��{�-�T*�L�}����M!$(겔�HD"���]6��P(�����z締C��;��a&���pE����e�C�Tbě�dm���fApB�'(겔ʲR)-��������d�7i�<�ٛ��B��%����H��!vo�O^��Y/����!�;��:��U&8��"��(겔_:#��?����.I6p��]	LB�� ~A�,�5����q1�R*���z�3o:p����!�!҈�JG!�E]����u��6N�td�Ő� �5K�u�u��%IQ ���	qg�m������r�j�Q��R��[f����p�BH!AQG!��#v�jAǯ�
��t�<:���Æ�d%(�|۷��MQG!y	E!�d��[�Mi;���f����B����T̘('.�����(��<}�qu�������8S�BH�$%��^OV�ض��
<��{��];0��Dۄ����	�
�W{��vU=X�4_C(��L���	�GL�d̮U��X̟A�nX��y�`���i?����X�q;G���m�,38�T���"�F݀�����	�VӇǅ�6��!I������ yPV3h/ȶ	!�I&��CVg�}b|�Y��`���w6�uy���0n(��^�}�qȓ�i�dJOO�yd���¯�L>q5�}@�$V7�T�h�D���"� x �3N�}Z��$Fy��W��{�V���>��3�Y��2�6!��Ȕ�B���0�x�6����7�E]� +/n2u��ȸ����y��3�Aԩ�}	�^B��%e�3X��%�����G��.�����j)��	!�E&�~Ga�H�/��bN���|����Ж8�Y��MR� _��B��{?f�a��o�b���e�B�V2%�0�ł��{(��S	����)E]�I�6��z�UΘt��͈xB�3�?>�u#�OB�q2)�0'���]�Q�Z��U���k���u�ʠw��x�+�a��l>�M��u��;'n<q���..O%o�I��m��t�
���po�>�}ń(�Br�L�+�0�p�[���y!��E]��ڌ��p9�D)�9�?�3��e����n�n"�=k�b&| ���a�����U�"D�'��KdR\��Ƃ��AY7����i<ɘ�曰���C��/1�a)�ൖH5�h�Qt�X���g��F'3�%�c��
��`���	!��
��+/1']Q�7m~71n���@5�uyN<5�W���v��TQ����e7�Nɞ�O?����,��?�_n���Cr�\3���`�Vp�<�wu�Br�D�J�՜��q��06����:Y>z�P�9�Ϊ��-���������TC��cIC��N�n�tC�NS�����RQ�����}���M��*��p�'��BH��J��-fڃ�A���aP�--� ����R��ytd�?I�!VzEƗ�%�� ƍ�B��%��q�<��a�k'֍�U�@�;�S#���?qi��K����B!$U2i1üT%�3�=j�nr��3D�.��C���������@Ow׵�����	M��e�� �7���x��͙(�%�����,���칋�օBl�B!�ȴ�L�+ю����_�f>CQ��p����8�$&l��R�
J�J�.a鸎��!�BH�i��99�O3�:B!�BI�LY�̞d�J�e����:B!�B��m1�xӮ�?|!���c�^�����ˢ��E!΅mRY>8�㔉����*�W;�.!�B��L��`�����.�X �X���7|r�U:;:$bI���t�ty�ݏ�Ӈ���.!�R(d�b�6��vj�Os��|�������V���J,I�͵ӧ��ߟd����P`2kEե|��!$����5y��bҌڱe	1>o�Bm�<,$�&��,�zbng���I�Sk���c���=o�6����Xp�Ȥh�}>�����.�4o���z���.C7��m�r��s��H&�Le�b��2������#u�(��|f�ZZ��b�*�0߸�v%2�Ց�b�f=i��b!`Y+��Q��DYqL9J$�ʛ�O7�%��˄�2&���p ��b� �͢"m`тQogm��^��˷I��K�%��1�'�wӇ�n����7�������|���%��#�B� z��Č1	Od1�d��:�HC.��v"
� �����Tn��T�G_����a����)���1���1�zhf�����?���
s&����Uj�J���y���e���&+n�)e�E�7����E�3�q*V\��������	�ځ���{+_k�Q�B!�dL��.�=n!�COJMԭ�hݢ�_eU���@(b_N\��W����O��2-�v�?�D��?&�X�Qh�� u�z[��,� ��D.�A1��Fv��Wj�J���Dyp�Ly��)ٶg��>xX�_9��0�^�tve�Z�)T<�3�J�~���4u��!ݥR~5�:,}E�i���^J��$��x���%v1fLL!d�D[��(ڃ0H���#�c׮�f7MXӴ�(�����f�mq܉b����	�K��`a,Y���Q����P,rpfLTKKg���"�'���[����a�S>�c����}���93u��!�\$��h���@��*��#3nS��l��irz�ra�t���I8�h���5��w!��;���范N�qfں�8>�
��]
{��X̠��&�ɹ��iˡ�J*17`�3[⬨�+Kn�[q��LZ��P;06��٧��x�}��1c���k�,1D�t+��%��|���� �"(1��.�]�:@QGH����Ł,:�t�Vǧެ^w�T��7�O�;s���%����٦��ٲ�J��d(��I��]0X�Rbb�Nh���c��N��ר~���cj���""�1b=D���t��\���:+����Ձ?��)�� �~��[ԙ�w�E!y���*�j�NX!�(�!~2�,��d�.�~�}C�4`1�;��D�, � �pf7Ns{U�`��=s�%�S�K$ˀ���x�G(��s�X����'��vt�?��PI>�qS5�P� MW��AŨmzz��x]:����tK�uG���巆�7�s��S���[�^o�$S�dsL�S ��A�	�f��k�N�J�'���o fk������X�%�WZVv�'��.\M�~e\HH0��rLN�� �V2A�W��+?�!�OT"c�9\9��0�5i��-�4��3����D�Xt&�t�� .�IڡV�׃�Cܟ!�e�4.�Y1���w0����O��P(T�F�4S���y���|�d9�`%��z]"�O+h#��p��7&���,%]W��2\"K��6���������^I[�9i�BR�L� K�X*�	� FH%4�ǯ�׫Zl)�K��&J��\faf=�qX��ݢ3]ډ�e邔�� Z��x"p�2Q|B*B�Jz�*��N�X��awp�_!�d���}��)oߐ��I��$n�ü���}�#!���y��Úf�P�tnu�$�W��֤,��;W����ʄE���U���#�B!���$�ʹ!Obֲ��$w��#�B!���S�}@��J�W&PV:S�ARP�B!��@�k��X]eIa@QG!�B!9E!�8S�kdʈ!�B
���˕<+|NQG!̜	�e��{���D!��B����t�sy%�&N�x5g� *++�kkk�������B�Pv<����BHA1{�(y���dճ/I�@K!y��o=�
�Z��Qd��^Z��>���Mdl���Z�A�2c���`��/�ׇC6�-/�5h�(���梴���~����ˊ�v�RG!������_�|����D/�2s��	�a�u��z��^�����,kafʹ�m��P��r�O^V�v>�y����a�;��\�k��/��lqw<��1u�B
��Br��-�-R��,� DX]E�_���[��.��D�U�A��3 �O%}2>A��! ��@`BB�xj0�ԢB!��&u�`py�����Ġ��9�BDc��uS��s��B!dx(�)0�K�x�2���->�YӇ�Ӳ�Ab��2g`L!�BHr(�)0`�j����3?|A�l�D)���0�IR�hft��Y4ڶw�l%�Rq�$�B)t(�!I��S�S�E�o�Pg�T�Ol����*�bF��g�C�X��~�B!��:B
X�҉UӂLe¼�:ٸ��x"s��d���@�S%`I��G!�R�P�R`��HY��F�(��jZ}�e��.90h_�|��S�_?eP�:��B�]:�!�B)4(�)0��R�N.�o+�t;����z;�N|�*n@�ڃ��N8B!��ᡨ#��� C]8U����+�,n��A�i�I��-v(m��%�A ��9�PG)4��ר��S���s�$�r���B�N_����`��3g�hc�^O�33�c}����#B��#� �{�W�����!�l����ֺ��z8��O	D�Y*!!վL�a>N����<�d��k�h�3q�Ԕ�������!^�>)�Q�/_�p�}t��LQ��3dh?�tv��9tR	�|�#'<~�]��;��x��WdǛ��n�^6��g��;{ze���&?}�C5>w<�L�9��cϿ��ͺ~E�.��a�-3e���������^���������}j=xl������o�_o>�m��-���F�c�1c���gʉ˭������w4,S�֯xj�:v<8�~�g��Ot����r����\x���#��?,�[�z�\	�Br��U|o�z��l����<g��=i�Ng�L�T�[���v@,&+o@��S�Je������N�Pq��G$
��FGw�t��Ji�a	�'C}�=r{�a�W0y\}�<C��H*✀I*L�1��}�<cLn!dr�eF-��O���ƾ��0�Gm3DF>Z�0� v�k�!| � �c�!n��t���H��:-r ���t�s�{����o2����Ȃ�t�Ѷy=��zX�1V���m�1b�pXf��m+�c����C��1O��Ա����|�����_���*��G�|y���~*�qS��'�U�Ͼ�\m�q\xb|��1��u�B$��%]���nҵ3��"��$e*�$�ʙ��Jg�Y˛!�7�V���]��"���y�1!���K�k�&�Xc۞�s��R�������P�-ܬ�Z��*�cb�R�Q.�X �*֐��N�=�}�;�v�Nm{��59����q�և���hA��7���v�6g��ScWO��2�;�B�_�	(�!����vJ����HQ��yդ�k�L�6|�6�EJ"���o�~��l߳O�� Ŝ�'�R}ѝ+،vc���a�^�"j�,f�����x `;/�{DY~a	6�_�,^*\�l�X��} C�����"iuK��cv���p�4o�s�;���h4$�.�wʫ��&;|�YY���ߕu~@�O�;)!~BQG!9�.9�.`2z�;����j���>c镪�	R\Z+d(�
�Z�e.0	�t�]j�Mna��f� ��{,G\�0δ��������"��e�qiE�~�&�W�yQ}�f�8�M�|#�^�m����/�c��Y�#�N?X���B뵘�k� sL��c��b�������a�1AP�عUϾ�����S��Y��[�����/�ԭ|z��{�<���xL�'�W��?|AV�2k��D�b����;��*L��:B!�Ģ}���+�XL�Q'a�3�>4&5Q5�)�-䏮o^ły�v���L%w���+Y����d�!H��}���97O3D`œ��k��XQ	D��Ԑ�Xv�!T��J��uvV+�cL�^%bf������sJ�����������X�;(���ڕ�����(��P�B����Dj믑�1I)..��2���弜9sH����ȱ3%�H��bN"��@t��CJ�m��eɜ$#[��|���D��L�������E�hK�C��	I|'X�,�#�x��x���P�B��~�)�9d}U�h��>�_Ξ��L��))*�P�uwwK��I�9�_. �	��#j�4?����g�u.��̩�3�ϚIr�qL86�����H2,����鑋W����_ƷQ.��Zs6S-�N(�!��b�r��a9{r���t�!�
'�
�u��\Ǯj�m�7wL��7gd�50)��ʤ˪]vH$��u˴�$�����Y��FKQG����B�kƎ�A���������qR?+�.�4���s��</̍d(H����eu��{}�v@p_��ms���O�Bc��3Q�OBܒ����B|e��OI��c�u��T�^���1�tV�)�/�N��d_�㪷���X�襰��'�l�S�Hh�,��9C�j"��hn��Jة���e�p�5'@��Qܛ�p�EB}_�h���Ol��qW�,�$?��#����f��핎N���>ii�Pƌ����1a}�R�@D�>xDձzͦ`s"��i�;F�8��W�Ώ,�8�g�	1����b��uA����.z�
c|�S�c��2�Ȕo�@Hn7^Ǌ{Vr회k��AĹ�����B�k*++����~�\��WN{�vb+�}��E%׀0���aiy����3���c��u� ұ�+�0I�5ˋ�(~�ъ[f�b����*&�~Ʋ�Ya}�M�˼�d�b�E!��G�d┹r��>5�[J�륻�\Tu�@�/�\� `�I�M/�w��
��ҵ�Tf�ŷ�v=LG�y����>B6B,�|��܊;��ç|Y{m,�t��C��BP�m�b����k�6�	�/�K��c�I�:B!CGJ��l��!RT*�'�$��~(}�HQ$&�e��s��~�#��v���?��{�᳷)WQ7�v�l
b�
�b��7�d�n�������(����Y-�ee�neUی>I�X�5�`Q�*N�\c`��X,���p�������z��1�����B�@�8�!�p�9�N c��㇫0��z�m5&u�AB������B|�f�Jع��Q� �����6)��H(��r��8r+X0�D�[B7`��:f�n,Rv.�$I7)
&�8���M�2���Բ���dܫ�:�K�!�&�ւ֩ �c�^&��k�����9"�za�����0���N��� �-�)<�I5�	�@���k�W�߃v3HaCQG!y�ƥ�b��-�ʾ����/�����q��?�S]����hTB�L�+U��	�`����Y3�������25at
\)!x��X��8_XU~�A�B�ќo?�,�fW*���8K/ĉ���|N��s�}2k2=zU~V6X[q�ZHa4q�1�u���P�B�3�"t����¡6);s����$*�Cm��CG�����=+�b�ܸ]B��J�X��m��l��3��):#��K��v"75�o?h*M�)�Gp5u#��7^�:klU�V�L�sŽ��ӽ.���_��K�-�ΪJ
�:B�a���wjI��WE��UX�u����".O��e�-`1D���2�� ��jw�:Lt1��&ᢅ���+��"
�6���ǞE	o����+�a�M4�f�W;p�c4[1FP3.�v�n�R�g�x�JG�BQG!�XX���=&�?��L�:Q�a��붵�I&&�n,��(�48&XQ��I,چŷ�up��c`"����'R+��U�l�
. ���ڼ��eELtTɍK��Lpq@��q�
��Vu�l���y��B$}(�!�Ȏ�<��d]*@�!q�SWL=A����|tXG���qn��̻��Ä}ת/������l�3�*"�m{����J��v"�q�C���h�����b_XplڵY[�i��-j����5A�KQG!����q"\tz�\ ����%D��	���mpզW�Κ��چ1Z��\6�G�eV�Ź�춧
�ϟ��	k� �~�H��(�#��۩�����E�N����\;�.�*��z�i�CH�ˆ����E!�bb�C��N�e�t��ǉAܠ&�Y膋qD<�W�7T��o<���Ȅ	�O�V�+��o��6P�M�uy�dXE���ƣ{�i-�0n��ֺT��%La��$��B ���
[���uK	;��cN�ݖ����	�7ե��q$
v���r�� ����|g��S�~1t/�C$c�ML)������t�/�18�����S���⌱`���
�_�?-�(�!����t�b2�	0q��C;���,��aӋ�;u��:u ��*9
�]@w�3q��"��Y�L����1��W�b y�5q
\kO�Bk8w�h%��ͮJ2K���B�N�����l�v�
�򇉦������L�� ��V���N@,jk�)�x)]x�����uA~׮õ��F쵅.���+o����C�`[;�M����ݴ��,A	;�:B!d '�s$x�u�f���|����!LSu�QL���f�<%f
0
*�]�ᒉ>�+ӣ����A��ZE�3��RM��qg�bF�~���r� �E!�2�5{�p<��{�@�͙8ʳ�)�~�R����с	�q���d�Į�5�NHc��!��_������!�c����DU�.��|-5p�gG�w�vu�B��#Q�'�n�Ŝ��&�n-^&N���k�O�פrmR��9q^�Z�`�Lep�4�\�1�"��~�� �����������gm/�񡱳���"�㧰��#�BD	���M�[;ae�n�q7��gJT�9t�?���7{�?��87Ba�1�NU��i���%y�\-�r	��9�l�����3�{�Ə�uv ��J�r���cOu| �p��CY�<�K�Q�B!b��.�t~���L�MPHۭ%�0�K?�����H�X��:�Ŏ�������~Ԯ���~Ƨ��^�J]qxk��7�J�o�!�(�!�q6�Ǥ<�0ۻ~����z&�Dpp�1O�~欏Ȋ�WY���c��d�:?���͙�,f��9D.�,���uy����BqȕN�ie
�ab���@1���M'�Gkm2;V��n�]��k@������e�;l2_��hg��SH�_�L"C2����B!q`ep.�r��8����D�l����If^�[x%�(�!���ضBE��IA�)� ]��$��ɚ�U�:���	Ɔy���u1Ib�vu�BQ�:�^��{[����&b�PDz����"��lz�Kf�Ry�vhgIv���)��m:aE�.u�Ȓ��R��B"]aGQG!�8�67��0�|ͧzS�=(��a�m�>���Hn��5a���;h��5L�e4t�7���iRM�����1XDQ���KX�En��V}!����u~�U��=�N��]��\�6�#�(�!�q6�a̙��l��W���t�yX�|�)�e��L��}��a?k���).��p�3g�D�Gs.	�Ar<�CM����F�)�C8I���~�����*q@aW�vu�B�8���7wC�]�~���&��|o��M,�k�Ǆ�N5�섃X��j燨���c�G?���,jҭ]�(%D����ڸ_:)�ˤ9[&��p٥�/�;�:B!D��.t�~T> +�V)LFw<웋i�,�}��ʱā���u07k��	���_�m��֮�&�;|uw�<`�X����B qY��Qa�����s�
X��
���iҘ�)Ydq�%s�=w��Ch��hY���<�bj�X�b�L$�Y9� !�N�:��U��J�u�<�+?�����n�[�p/�f�˂ĉ���#�B������ŕ��k^΋:�+D��`R��=w���$���[f9�>մ�p���K �:^�Y½���&�i"��?�]�_ԁU�ڻ~E\ܤS�n��#��% ���K��6�O_p�\B�`D�"�x@}N��T�E!�2���f<��UWCX�y��/sU�BD����p:i�eԜ0���MYo��y���jy
�R��1�̶W���A׮s
��Y�q���@������3o���>�᳷Ƴ�"��	RH*��B@���?��a5X����k`b�{ս��`���G�DpA3'����%��;��	IV[#�J����������@H�p�m|ة��� ��&i��u�_WV�4��W�0k������v�C������6A�/�	;�:B!d <��S/�&��8�)� ��N�3pG��	��aB��J�ɂ"�oV�򖙆�IO�-�$�A�
E��Z�g����C����)p{5Ǫ�t3kj ��\��Z���f�$��]D
��E!�bt')��!W��zr���eF	�����mϥ�?��W��q"x���T��5՜��+^����[f�6Cȸ�7��;r&�,��j��s#v ���z_���n���
ƼS���E��<�$K�#����#�BL`��$f.%A�x7�.19�0��]�F��W��o �pP�@$8.�Hq?g�(%4�\���M���&c�f����\��u�E׮�L�v1vS�/k��X���ͩ�����5x�/_w�����{�1�>���N�Q�B!6����Y�@b��քl���L4a-YѸKe#t:��a��4q��x)3xx������F�i`��Z��o�FݷT���!�.Z���2��}��k���ƳٝSa��(!�L`�:7]�~��9)��XK�����j�xVaGQG!�X��w����L�1�#&�n3]��'�zB��21�,� |`�r
�t�d&��6' �k��i<�EV?�~q��e\K�?@��K����V��S1�kdWcd��h�@F�T3�&(0�����!!��XUl�����E�!DX�{ ���T��2gC�;���4��I�Y�Q�B!68����lv8�:X}��Lpa�q�7@;X\�ʊ�.�Ļ�
a�=M�lm��6�M`�k��*� B �ƣ�\!�!�>��p�*U��N4��w�\<qcm��ƥy)�����O�-�(�!�0�[9���lv�Y��v-��>��2���u�M�r%�V��Lgu+耛x)+�������	��$���c1��)�VAg�L�v�4[�܂qk%b���m]9��_nBR��BI D�]�M20��s�$e�ʄ�!�J:Y.SqC���q����D1e�g���K�A����:��"=?���7�U�}�����֮�p�����;�[�Z����:k0n����;�҉�n�:�k��̠�>��D�mY��Ld%�E!�� X'0�vc���l��Qj�dZr����(W���\� � F�Z��Fw��TeلE�1���4����������P��3�6�86�,�Nȸ9w�h[�O�1Ch�Z�eb�ly���K�Wh����$�,������J�*17`!�cJ��e�U��u�B�0@�����*�]1��ㄏ.U8���F%rp�.]�$A&�v�[���"�S�T�)��#X_��t[���y���Eg���jz����.���ע7�[�y����bH�[(�!��$�M���-3�q�'�^&	���uN�YтΩ`.1� ���ۦ���[&���nAp�x��3�?-f��t��BQG!�$!�T�f���dq��#���aW"e��*C^:V'�[A��J؁�b�w�V�]F?�}Щ��d�ѭ�e���B3p�����s�}\��7�N	]X�P� �l�@I܁q�4�3kL`�.�$?��#�"+���ݓ�(V.�TIsU�Ģ�!�V�*�J*�5
IkW�L��:p�C���H����O��(�.9�}�hA>Lܛ�I�Y\�b�"*]k��t�F�tNX�(�`�귞\�G 1b�C!E�bW��[`�k��g�^�@&��^ƒ��0Ǻ➻���\�t�A���t��#��F��[J�.I��Q7Nr������*��#fI���ɒF�TɌ�1R_\麝�!�||����Q�Q'9���Όj3$p����px%�4iX��
��(�84k/�=����5'/�w����fe���W�|��G����K�b���"�p����핮�^)�8�~%���_><u�߀����E)-�����M#MkHi�}'?��[���^^7Y6�~M��j�B�<쳮�Lm��;X��[��m�"Cȉ�$j���Z�(M?���e�vA㶦V*`�H��@y6��L�<���k��C  >�g�z/+K���V�v�V첏zJۇ��V��O�ȑ��F=k�:��Y�l?ky'$�B,&�KS,�i6��ɴP(<��	]
�M~E!��?|A��m�l\�@	���Nz��KKd��ý�'/�t�Ģ�r���?wD��kd�\�������-쐒<l0��uֆb���9�G?0�'�.qh_gI�˞�����x�r��N=;�=��5�F�!,��xS<����fi��� ���ZJ��%��C���iYx���R��d��C����3x��a���/��,��:�0��~���D[�Xט��l���DB��ZC�N��(�!$C�������N�x%�aB,���ݷHm��4�sƏ$�^��=9�P8"��r��n�T�ǬO�����˄)s]�ǿ��Aaw�;dGò�q���̠�`�>2ǆe;z�şqS�yX��/a��
d��x\�PBB�g�z�Y����k]� .��I~?T����j��6����Y�k���bL��=�I��f1�� ��h����v�m� ���E7�?���񇷮k6~����T��l���F��E!��l�Q��~ ��	���y^P5�Z)�?d���7H�كr���R?z�2:9
Yo2&n��9����̡����6��v~��������+�]�_�j*�>Ix��:�N�uՈ=�GK$Ա�ec�#N���������}Q�����f�9NJK�d��R\Z��1hA��)���C�Pr���p����'v��.MW8�"f�f�Xhc�_������o��5EJح���#��D9� �%�^ď�ȱ3�ܩr��o���D��HIi��D(���#k!&x�f�C\�zg���N'���9����\��:7����:	���~���Y��� 2p��%&�-�[C�!�c�Z*����Xo���z�p ����UŇ%Zo����_= �P�P�w���>��?K	W���0#�,�������9a���v�:\�s��M��?~a��W��񢓜��4��Ƶ��+�5�4����-��r������j	G���弜<���Ս��Q�����i:nO�_~e��]��z��EŔã%���XL��D�~w���խ뚍o�U�ln
K����L[US�BH��0_���#@��Ek��_��ܤy��vB�z��s2f\���a�G0&���������nX|[�-R�:m{u_�ʓ`ҌI2ĂrI3&�w:�^};�b�`��u���Ч8s?�2��Å�!n���Tv�\*��J��(��\Q-q| �М,�q,��q7t}�:�g�ƏG�Z��S�ں~�w�04'ځ�����h�$���87��קt��z���Ei�x.�*����HiQ��A_��W���uV��ij��ˈ1Cc��jF�����KW�>?y����������<�hDD�U�!� �y�a�߿wt-}х�ĺf���Y���E�pS���BrX>�Z��C��MU�4�D"���c�%%�3�� �J`Ʉ��dV�l���.}P[������eV��K˦_���3kL$��Y����eW���09�v�vq|�L[�2C����u=
��?5�(�	�ڰvM���>!��YJZ`=�����8f����Ht�:��,������];wXX�̥=r���>%��Vc�� %eu���%��J���:/nw 
� ��6=-~t[�tX�vu��� �%2����e%���'r��{2f�L)-���s.��&���z]�M��ܮ�G��}Њ��a����~<�O)A%�	
�DD��:�\&?{� ��c��Z*}����Gb�Dq|v�y��n��S�����U��Bf�=ރemH���ǃ�f���\�'��;���^���k*,}ϼ��%&F��^N��\m;穨õĒJVJ?x��7���w~<�D]W_ty�NaW��憈��vu����Ee���)� ���RZ1�vQ9s�}1j�T׌�&�*��ٗ������aV�@�`�	Q��������@�ud��y�$ی���I;��~�m�|rV�� 8ஸb�a�@[oͥ���J��5?����4h��cC�S�o�|cH�����C|���a�������hF�ˏ�O�O��i��8��c�z}N8fm13����Y*��"�������S�9(��~¨��<�o�z8��GyE��Ec���7��z�������9X�𛇤)^�aF%�еu�Q	�b�<�u���)u����	%�Y �t����}i�,���>Ǡ��.f[\Z/&�(gO�+-����q�IIi�tv�I_o����O�{�;�P�N !X���R��6�[�E�%�w,�ﺯtY�������/���1�|�d�8��+%��g���h^���&Xo�R_���eþ�YdC|Zף��P뿶���X�;�h���|���}��e��rN�DKK���뤭�tuu��+��	1)���~�QY��{q�b�3ǔ[K����=�n�d����ƚ�p�7L�:B�1�J��hA��a�L�aW��i�I�)9{� �?���Ĥ��Lm���Duo���t0��|��d
��q�h=D�]�����,���'�7����\���J���f���땓�ޖ1c%ma��^�O��N��*ɬo�r�zEW_�A2��uͱ��׆B᧜~���Br<�D�8��/�K
���?�}� �1�k����늴�����΁���W!�d7(y0i�͆���!����}g�Y��j�n�����y�����$va:6�R`�\�5�x�d�b�|&�.���]�#[�8��Q�BH�J��A�Y�d��(k�����3Ӡ�mEu����D RT*�+a!���\}�n���Ⅳ�且�����y-;U��lvMkHX|\ǉ�"� ��	�w�E%{h��uu��#�GOo5�����E3�v��B��/���4�όk(!�"5#o����?_^Q+�ܤ^_�xH�B�bє����&�ıX1ǉ��.l��x�D%�%􆣍��0E!��*e�R4�'�)�47A�-}R:bp����}�iU���"Ο�Z���޾��K�IiɈ���KH1~D!�xO8ҟ�S'�rC�!ގv\��{;������W1N*�[%U ��bib*Fn����.�4������e0R&&M�E��A�#[�8q���#�"_�����@!����<2^��¡6	������{]�]�>k�+cw�;Kef�j<;�`]s��k���@e���'%b1�'��fH�Ius�:B!�B򈯿|ɲ搐�D��&�2 4Cu�B!��D:��$%B���Vq�ِ��B4u�B)h��A-��t�*�: N�?��APZq;�����7��/a=K�Rݞ��B!$�h�u�O�!�xE!������ 0�wm�z	���m��zw?kmB�(q����뺯_HrT��E�%.�[^~K�;BH�PY$��%�2`���⠬+E!���+��$��M ܏^��jj��B�B�@QG!�� D���\u8vZ蜃~C��pi�	!����e��.�yN���#�B���X &�MkP�ސ�F�`��N�BH��T@BH:ٜ��BI���ar�DX0��K&�7���z�1�-�N\�F���_8P~S���y���:�E!�Y9�^�\����*i�*�X46d۪X�TI���B!i��	�c�U�u��]v[�t<�NTq�Lԩ��-R��6x��<�|�?�bжX���2-�}�D��|�D�R��`u���ie��:X"�Ȑ �*z�X?����^aB�VB"�U�l^���u;%(��F!�<t7����?\U"�G̒v	K~�F�TɌ�1R_\麝�!�||����Q�Q'Y�tH�a�v�?�g`�N��6�_��Ab�襖�k���w�L&,B}fp8_d}����j>?��ZQI�!$�	ǔ��
Qg���u�B����zۥ�r"1�®��V*J�=�w.�|��oӇ��a�J5a����2�-|m��ji��e{~a��c�����8&}�Zܚ+��gt_�<�4>�ϛE1!�d���S�f󴮭�f�8��on�����(�!�$'�������#RV^#c'��zWϼ!��.] `�3��Q�d	S v��Ѯ��7�����.��l-`~bv�8��� ���A3Ě>��%���f�����[r;E!$�)���$��uk6ׅB�-n>JQG!FOz�3��A:6
�[�����R�/]0d��P8"��r��n�T�����;}|�L�2��>{{Z%WЖ2;+�ov�.a�]�p�2� �jVЦ��m���ǂq�q��h���$��S���猯#�d+��ܝ�غ���F7V:@QG!Y&�:)��pC$������%C✴�&�n]Ոk��r���#F� }gʥ�K���ϘE�-�t���D��oZ}���k�������D�K��)�N[��p�i~㒢��̈́%�X���W��n_��BL�n���S�BH�0����DJ���D�v�3'��d[�@���;SΝ: ��V��K��~���VKQQ�J���k���H�0�3K&b��2M]EY�u���a�� ڍ�B� KYQ_�Q�l^([�5�&J��F�i@QG!Y,m���n�=�o�*�ރ��v�H�O��P("�&͓����sU�Z�ɘqU�%�I>��tN�g�GB�}B!��&nj	@�A�E�Mn�.5u���������b��=�o�j�I$����Hoo��DJ%_��Ji�V�T����%����K�ߖ1�u�l��X���H!f���}ts�_��p���.]A(�!$�Ѯ�p��r�gd+�q�DN�|Oƌ�)��5����t ��M%�p�L[gFתõ�u��@G��g�A'OA;*qO�̖�w��#��v��U�����'��*+�-k6�$EqCg���B����zx���Kx��02)e��%�Ҋ�2aRHN�x_F��&�5c%��צpis�:'�"��ە��>�(��|LUV7[�(�]wO�ډ6���LQG�5`E�b�k�o]��nl�޺�t���Ѕ���*BQG!Y&��7!6�Ƅ>�K�F�"ŵ2a�r����r���w���VJgG�tw�KG�e�]o��I52���޽�u�g��u�F�$ ^,RwH�)�%ږɲMHv��e��Ue'k���k��5�d+n��$Y��쌦*+��dU^'��b{[2�SQI3�K6%Q )RE��w�{�y�n6�@_��sN��S�>�o������v��t%@��_n��Bz����������ņP�3}O����oeQz�~�:m[�����p��4 H*mw�l����ϳ������ηӦ�MM;r�pW�a�#�@L�~�P�͚e�=��/���
j��*��knYk]�A;3zԎ}��M�6?7c�T�֭=;�j6�T�ۛ�7�W>��t�s���_�|~ۊBzl���O�*��a,������������i�80�ʫ��7_�$S�KYz{g�=�U��ڀ�2������6m˅�n�Z��q�����P 1����j����cbjɕ,} �֨��W�Tȋb�3�����2�5;=b�G�"*g�K��c��t�c�!�/�R��r�M�����3�v���3Xd�R��9���{ k�ͫ��G����v�s/�Q��1 �$.����v�]��j�'�P 1��AA�����2����{����w#w�(��uZ��y����}MXSs��F�g�֙Ry����
��z������n��_8S!����\�.u�
�? �vu cj$�\s��qK��5��2����q�W���*��ī�L|U�������ﱗ  A"�@���-5�MN=3>�ySKl_�˞��^w��0���vk[�9����옵57Ys.�Ukzn���3�n�bm��/����{�  @eu s
n~�O8pxq��V\jޗ.��0�����/�~a   �u �R�p�W��+)e�  H>B    $�    �P    	F�   �k޴iӖU�VE� Z[[������է��   ���:    H0B    $�    �P    	F�   �#�   @��     ��ޛ���eT ���徎[��Z�j��ի;g3Y����c�T}�Sٴ�6Fg�   �W���s�����z�W֯_����ı�U�����7    ���K    H0B��L��`G�}�   B��d�[m�k�   <�:    H0B    $�    �P    Q.;��u��~�����vz�Ł��   @b(�m<9hI���ӹo	,��    �Ԯ;>d��ٺ�졲nW��2��    Ԍt媧@��u    B׵�����{��6p��\sYɷ��@��u    B��w��Ĕ���?Y��?]���9�y�;B   ���?���~���\t���t���L��m|�ƲoK�+AKK��}�n    *Rn��5g�������r�5�<��/�ۋ߷q�   @��J������7t��w?��^�2    ��k[/��_eMM����Դ���q{湷,w�m���\����N���=j�<��B�+����a�    >2Y�3���eK����q�'��С���_�;?og�L���P��׏Y63oa"�   �;~|��o�tA��+��L&��)�P�?>d�ׯY��#�r�6B   �:���ǎ��|��K3��w��(7�@'�:    H0B   ���}�G���     �u    ��ɡI���;粖t�Z[[�-��H���s�mj	�\!�   �o�k�O�wy:�d]Е�)�����;�r��(7�+w���P    �R�-�$���c����l�K�����fs�Y׺�&B   �D;�����7;r4�r��x䰅�P    	F�   �#�   @��    ����]ikϜ�F�I7���+�-�   @,��pq��[������)нv�'m������    �V��j��    �Z�� ��    �^�����    $B�� ��    $�v��;hIu��P    Q֍��Փ#�TkΜ���:    �C��Ɠ��dg��޲��X=B   �D��@��u    b���T�#�   ��zt^��P    ��9�y�;B   �X���+u�<��֏��ڍeߖP    �֜�F�>>L�   �FC�   �h���B�~�U��T<�LMM�˯�g�{+��"�   H�L����m��e���G��i;t�e��(��   @����ö~C����Q��z�2�L�0�UT��
�   @����c�mn>s��+�r�"�   @��     �u    �`�:    u��ФM�̝sYK:c��-uY��    ԅ7ߵ�'�λ<�n��.���N���\�P    �R�-�$���c'���3�pU��u    ����K8j���Ѻ(��    �P    4{��zo���V���������d�   @(�~�N�'����OX��N�uǇ\����'� �   �����^��G�x��{?�.Wo���rN��J[{�5�L��F�_X�m	u    �s�e[z
q
y�.��]���sz�Źo��z�@���������nO�   P3�C�e_����@'�:    �V��.�@'�:    �Wo�.�@'�:    ����a;n����/u�8���)��tB�   �SW��Z%���S6�wВ��
,�	�   @�/�ޟ���oS�uc'����w~i�/�@`�G�   ��S#n/��]v�9�xrВL���Վ]|} �G�   �������ꮅ��!�   M��6���	�z��e���z���-�����+Υ��@�]�喪��   @(�]r����.�i�q�t�����l�(:��D�#�   E��?�kn��+�]w|�:��)�)�����N�niPρΫ6��    N{�uo�t�.�����w]�{�����i�{��W�>�y
v3���˾-�   @���J��y��PKm]���^���U��ǚ3C�H�Ǉ	u    ����׏�C�   ��)�]C0����)�g���۔�׶^h�o�ʚ��Ǜ��i{�����soYP�*��   @�|o�F���'��K�7����[�ߦ\��ٙ�Q۲��Z[Ϗ8��v��Q�f����-D�   8��i>���-��i�KͱSo���=z�����ö~C����Q��z�2�L�0�UT��
�   @(v}�	�3�P��
���_8����r�x��*���ǎ��|��K3WT�E�   ��6W��}�G.�:�:    �Q��6��(�s�4�N�/�KW��8JG�   
ma�M�5gN
C�.�1����U9��q�    �B�(��!�O<{�������1���){��̓C�6=3w�e-錵��X��*Wu    �a��[i]�վjq(f5��1��?1t���t�]tAW�pVT�z�:    ���2�ݯv�-��B]�6����e�+�d��؉a��6\EUn!B   ��OL�x��=�Ɓ7��pԼّ����-D�   8�4�n�P�B*�@��P    p~�V�\)��a����    N�ϕS�R���חB`5��42B   �P���nh��,����F�u�:��~xf�x��]�!�Z:3o�n�m������nK�   ���i����;o�7n]f�i�����-4��n�]�ɺv
t���oO�   �5�S�/�3'
t�̡��`Wm�B   ��P��d1�zvA:!�   \����K5p���0�ނ]P�Nu    �@���O�u��G�V�,�^�]��Nu    �a�Ŷ1X�6+�����;�T��rY�   @��G	��]��(�u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#ԡ*�O��G^6ki���dldU����   ��UI��ܻGlÆW�m3#�  ��P�3gθ�qv
t'O�4�p�   ��P�@�`���iq155e�N�2   ����������1   ���-����Ӂ�_{[��tz�   ����6������V�ܴi��ޓo   5B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�5���_e���N	�~���O��mz�k;3d  ԃ�-[mt�U��:4�������\`��~z� �����w �z0ٵŒ�P��06l��S��x   �"�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:4��-i�⥭��ߦ�������   Q#ԡ!��ͮ\���6�m3    u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P��0�1;8�	��F�L   �:4�S��Gf���#�   �:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P����)e���~��Ρ   �F�k�;8>k#��@���l���u�)�� CݦM�u   �B]�8xf���ա������   ���     �u    �`�:    H0B    $�    �P�Ě�����)�d2���d�W��T*e   @#!�!�����,�ͺ���͹�u���   �PuH$���@�)����X[[�   ��P�DҐ�r.   ����9tn���   @#!�!��(����9=s---���j   @#!�!��JGG��C�W�$�  ��X
v�.�rl:c���Tp�x�   �8 �   @�����q;u��Ess�uvv   P�u��ɓ'-n�w݆   �W�:T-��N�����v   P�u��l{��u]`]�.���fl�}�   ��P���n����{-�f   �O�:    H0B    $�    �P ��ؖ�6ٵ�  ��]�-Iu ���n��  @4u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u "u���?�j��Z�lr|���W߱7G��> h<�: �Z�����T��e��Ykon2��� ���     �u    �`�: ei��#G��d0�FO���>bsss��MNN��![31S��gfglv������X�>/~�)����N<�b���-��,^�������W}��S�vf����}� �x��Pw��w���ޠ�o~���-W�u��kÀz� r�/���)[7L��>d�����uZ0�^{��_�/'���P}ڤ����]�7��`J�3��5{��]} Ш�6��(��yPw�>i-��r�PO��T ���ٮ��zkoow��袋������>|������CCCv��	�Fww�vs1
"���U�V���DC�'  ���Cݢ�����3��9rĀzSm Q������mݺ�.��[�~��.�`���y�fggmffƅ�~<x�~��_�L�D�P�
z���� ��5D�kii�իW��U@�K��O~�~�7~�� �.?p^SS��]�v���7o��o���8���ةS���^������z���� ��T(Lz}  c��0���G��m����*i浸��[յa��f�-�И��o��� r�ڗ��%��C���J��
&�y�ץ�^���v�m�ٱc�\X�>�"�'  �.D�Sǭ�����!YRss6;9i-s��8;H�:�� 
����k��~���f��׍��K�N
%���'���_1�DD*��/��.dEY���/�b������v  D�!B��h.I����5kָOÑ,����u۸q�ǩq>::z�r���� �s����	s��%�Vٴi���SQQ )��A$���!�q�O  p��ujt��4Tjݺu�a�dч jH��4I��S�+5�h�������=DԋT��QHa��+�t���ۿm===���]�A�����W���Q�  �T� ��� ��G�Gv�w�@�!���\�e~��_�����+��f�>	v  ���Sj ��+�����2�q���Y��'O�^�k���y�%�#�P�;  j�P�� �}�v��?����I�ya�@��O�ľ��o-nĝ/� B}�  �%B��J w�y��ܹӭ��\�ri��B���z���/�2� B}�
� �� ��� �T~я��D�O�  Q ԅH��k�˹��Z��A>33��V:.��}�)�xa�` @Tu!v�;��K�m���J���_C{��뮳���߯� ���g��7���q���l}>���gϞ%�#� BЀJ	 ڣOa���'n��JD.��"������kK�A$���e~���?��l};v,��  �!�huk��72\�z�n�!�Z�p~~�������̙3v�7ح��jO=�Ԓ�)�=�βo������p� �  ���� ���O�n��7���w��7ߴ���߱�^zi��`Ah��ܼy��a�'  8��9���j�җ�T�D4gR�n��u�h�����K���_�> ��u 577�=����!��a���\5,R��������4b}j~]X�	  �F����o��۷�U=�����p�|�w�}��/�l} ���B��H���h_�z[�g����`����~Gջ444d���'�����>��`�  G�Q*�r�h�m.����s�aU?�2/#�%׶m��p�F�U�BN�<iw�uW !���> @q��)���<�b�I�Z[[]��sW��A��g?�ن�U�|����ȲK���> ��u����][[���k�mRhԍ7���A|Æ�����>���B�yVP�	  �G�C(ԛ711�z����d��$���>g---�Un#�.��N�8Q��P�gU�  `y�:�J�0���\��B^�a���f����:;;�رcv�m�������oO}����  +#ԡ&�&''�'��wG�7>4�Id7��Գt���馛*
!�繪�O  �2BjJ+�jHZ{{;[#���?�qzO�h��ߐ\�nccceݞ�<W��	  VF�C�)ȍ����իݰL���*��_~9�A���ڒ����%ߎ�\��S�`�[�  �4�:DF�1�"*Iok����>粗�o��Sc����!�R�h��+�����Q�竴> @iu����t];=���!K���.���K��U@�e�֭eݎ�\Z��	  JC�C��%�%х^ȼ�"�������,���  �!�!���Ӗ4�k�R�>hа�rP��UR�  �4�:Ć��iULŵ���|�Y�����Y\%�	  JC�C��`�>v��J��i?E���y`�<�zI��>���> @iu���MMM��Q6�������cY���  �(�;�ӧ��   ���f�繯�l:�|�l8��tֺS��6�ZO*e7��Xu�%��i��   q���e����_�v�u�kj�M���Rf���u�%K  @\(�ͧ2{��=P����3ۛ�i���r�.�'�pG�Cli^�u �ѿ��oڗn�΀ �N��]����K�޳��\G�?Ͼf��OJ:6k6�ͦ��=���A��z�v���hv�n��P��Ro���K������d&>���ˇ��o���^��9��V��7�x���P��UR���/��8�\��cU����>�����Ѩ�:bK���������e��5E_�k��N|c��>�}��s������7��t���Y�]�kZ4%�NǾ��Ԧʟ�;���[�Z�9sư4�k��r��,����W/ƨ�GaN��8�\G��t~*Ѝ�gz�����3�ܽ������Lz��`G�C��f�<�B3�7==]��N곸J�^��3���3���6�����M��\G\�t����7�^�����<��u@v��s�}��������nG}.����gjL,נ ��:�Fs��3;j�<�����6Y�{������!�I�r��	ۼy��W&'�·<p�@Y��>�Vi} Pk��N��=X�r5���}�*]<�P��S��*����������]x��o���q[�v����Keݎ�\Z��	 @-iۂ3��U��s�=���J�a���_��(�h�JB�+��B}��>�ֽ��z�����z�  �mz>��ط{8{_߮T*�p�7%�!���g�yƾ�P��3��~��n���O�W��U�sA��5��_��^?b��F P��Y�~�.i�����-���P4��'O��N�^{-�挎��ᾕ��Ҽ:��W��O  j!���[|�[�s�uH���GC�^x�����mnn����uvv�O�ӊnO}�����U�g\t�nsC1�����,#�������.y��^�]�}��s��]w��n+�ձ�Cs���y�}�C�.`�����/9��W����7]m�_�t�Ǽ�g�������=N�I�<��	C|���?�W�����λ^��^瞽���Z��v���%o���}��ӹ�O�n�ۭ�^Uʹ^x��K.X�L���'�]�,=Ϟk.[|.�>� h�K-Tb11����d҄:�z<���O�=����C��z��ۦpV)��,էzYM}����h5h�&9���^�2�0G��>�#�X�ԈU S��u�.�u
{���Fr�S����]c���j��q�k�z
t����K)<N���+�qc��x�y�����U.�K.��^�R�\ra1wN(�W�*�\�?�{C�;�����������_�^�<��dm�bD[tܿo��!��:$�B]SS���������SO�G?�ц����{ϭ���c��1�>�
�>�QC�	O�#5
{C����rz��^G5Luu-�֩q�Fna#S�X5�ըu�s`}w��5�������!�u��U#</�U��u����a�ნ�PJ=�K�:��
G
T{K8G|��,(����s]���u|�{�������?�=��\�9^��J����ō�f��.�pB 7L�?��m߾�aC����
j�o��4�����>��8���,��@԰�A�5J�xv��\#:���5t��o��P���hw=u�������{
���!��{������F��:��Jy�ѹ��T������[ι�WK=�bCKWR��J&���Q�L� �뗿��k|_w�u9�Q�h�����'�ܟ�S+a~��l�`t}�� ���z;Dp��z�
�\���?�R��+�=�Oe��}T���^��R����+�Z)������T�ܳe�#�uC�B��YN�+�\_�ia�f���"�!47�yuᚚ����뿶����j��`
]
!���r��Ͽ����o���L05X\/�Ĕ���G
����<�K_5�ESw�BC�ͽ\��+��a����\,u�_���{�D��`ņ�\԰��#����W˝����A��z�^a-@���_%��������T�a��^��:$F�0C���7�\�cǎ��ի]�l}.E_�;�F@>�*�]�5���䵜��`.�R��0�{���?S�<*}/��Q�B)~�}���'&c�=j��?7x�綐��/~8b!�G�78/���,�}��s��{b��K}h�ܪ��Y�y�|�:$��Ԇ�=��Cn��64D�VgԊ�~�i���p�ҩ񪆈�����_V������]_t�g�B:�PWw�9��ł�B���o��C�<݇�~5� �I�~�(�����z+_Ƙ�S������9���ߋ
���M�u����,�}��s]��yr^h��w��4۶q��
��L��ҥO�C"dzY3�N���~���.�s=ӰH�T�����|'�2���}�j��3�O�Y��q(��!
{'\p�}�o ~�\a�ׇ8?�-(n��>�zF�CS��<��{����o���r�l���m1p����Ntn�+<�6�z �R��{Ҋ�GW���BŞ7�G�C"�|��Z���/�l�z�c��������v(��y�'�\jh�p���r�����]�6�2���0�{����[e�Rz�s�@��o���Ph�[f�e:�ԳV���Gt[d,(�Gn�\�/��R��r=���=��7�x��n�VU�g��J,����z�b�S�k�n+�xB��g����v��׻/4���l۶�n��&knn}�`~}����e�]-�s�̅�rC�)֐J��]��g>rvq;��T#x��N��a�����Vl��R�p�մ^�7cY>�-L�������W��=`~%�b���=�Z�d��]de�����:��A��Be�|b�g��C��&R�S��:Ğz�OW{��1��G>bO>�d]���n���m����裏֤L_�����π�O�}�F5DԘ��c���QH�G�׿U�m����_��b��󸫄�I�W��`�J!;.d�PJ�큘w���JC6�r��r��W:��y���CQf�
[�}�R+k�BbO��h�	ԞBH{{�}�pAdvv֒n˖-��/~������d�W>�gkk+�����n��S�������\ H��Y����v�����͙toٷ1 �O--|�y����$���^��K\ �bޗ�^R�ɡpX����߽��}-^6T?=� Ј�Y�b�rz˽��F���zvq
 �gr��'BZ�+S�����F5�,�@�(@�rMλ�v�uO��=��Xw__�z˽���E���]j�߻��VOD���'>���	�"��[�e_|ql��s�ƍ��O=���q���X�ƽ��Wc��l�<-��a���G��޾�D(A+�2�G[S��"�_���+�J�䦄:�ZRz����;���-[��U�V��>�1{���ȑ�/@���cw�q�e2���8�P̵k�&�>{,���4�o���t�?�-�}��{r{2��~�o���
wn�gd	�V��w����Ҿ\Z������(@�䚝ۣ�[�ќ�SI/��[---,�CSSSv��	��[\O�+����Ԯ�.�o��W_mo���=���G�@`bb���F}�G�c
U��������Es���[�ma_1��-?�k��ƾ.c	�`(4��L�ڤya�������j����L �t�}=���|-�U�����ޞP��R/�z?z]�p�M�6�s�=���n��Vף������~x�������g�*]F��Q��ˆkX��zs|O��S�SO!�0�燺��%�wA:���{�O�)k�O��ξ۷{�ej�t&Wfu�%ͥ��.���v:�v~��2��)*�/M��뮳W_}�~�X�P��P���!s�s��
r^��'  ��J�MM��;��Lz��a�����g���5������.G�S��52�k�f��뮻���_��4��𡡁'O��|��jP��ѐ9�ysA��#�����E.*�6�^X8C�mǍ[�����Ш�4Գ��;�r	� ,����k(��\����@'�:Ďz*��hs��to���<x�:::�s����Y��)Z���k�uy_q�v��i������˙���t��o��g�J��Ri(���K�+ĉ������^5C45oם7�ysn���B
Q
z�c�r�������������=��
7|�ֆ�Q�	 ��ԋ��o�{�k�J���}]��T<�����@e]�ɤlUkk(C\F�x�7'��nsaGC�4G��@��^�_��_wD���>��[92,����z�5�\Mժ>����ի]��^�T
X��la��k��G=X�S ��_E����_��S�{�����O.D�Ebr�ٯƩ���R�/%�ߣ(@2�-���uܷo�|*�g�����?�]���-@�:Ć��Ԟo�;�����W��Ұ��f�n^�(�|�����v�����GV�_j�G���/mr��".��R�k��"r~��[����܇ͷ|f��jU����YAY��~�z{��W���{,��Jܐȼ��n�d�2}�}�G�-Z�zs���_�>�|��[~/�׿��u�.��Pņ�Qn2�V���GV<N�r��@mh��fK�,�~��L�ؼ�/u��65omjڑ���s��2��������+��ȻvIg�FFFB_eT��رc��W������W����y�fף��ﭷ޲�G���ZR@�ܶuw�w6�~Ӳ�FU��N�էz�4�qfff񶱨϶ա��`T�S���D���W���PV��^{>��Bd�P@?ɣ׵�zM��<��p�����f{8����Ke3)�?.�mږqݖ������q��S����5���[��.����̴k��z	8�t��o�iq�zP������ r�m%����e���LOQ�*��j9�M�N=cjt����]_�=?|r�gG�R�S�~ΠGa�R���zE�U��e���LK� z.����v�]���RB"G����+>�ֽ��5�N�BH�-�QK�]k쿽�s��|�O��읉�����1k7�\�QK]vm��\}��U[��P/�B��WM
�P��ڹu�婜Z���Q���ϸ�Q�79wC.s�_ϱ^�Q�\ũ�L����~�?�"B"U/�Ns�^��K*�J�%�쳿y�9�Gh����e�Ƈj���7r7�炀��X���9�[,��E��nS�\��:\=���.|�Q�\ť�LHh�U�s � h�:DBaNC�V�.)���ؚ�v���� C�R����q,�H=�@�a���F�蹪u�~S?S��T�z���:�\nOI��M��{T{[���,ן_���'�5���^˿hL�C���{����#�F�_�R�/saÅ���!U���蹪u�~���v�EE>�y�|���U8�Y�Q����>���^g�ޤ�ʿ?��ms����x$��+}H�r�3��C�׊�"�HB��E��n�΅�W�{��&�b뙨�P3������ ����O��x^�����M̱�E%�>����C�G<���yznK��(k�)��TY*[�}�a�FLX�*DUn=WQ�����ܗ�p��^y�� TaG�K�g�;{�x��:�s����"��Q�QL�!^�W8��-�p476��k�Ø��-�*��q��u}������[����.W���?��~��^ޏ��?�A�;���zE�CM�;�b@�����`4Z}��Cr&5��/����	�f�¥6����h�o��j�y5Pܢ(���k�}�3�1)Ć��e�Q�\E�[�yQ�CZ���X��X�7nue�įt6^<o�ӽ�_�p�[�=e>䨞}o���?�¨g=W����P���|���*pz��<��P�P)�i�z�; >�'����y=F>�(x�J�qmp�aFn��\�M��Ay=�E�U#��E)���qs������~��^�b������\����z��ʵaЇN�}�=��ĉ��> ���>�C�g��.Ե��~��-H4����|�P��)�i��0��"ņ �rטPO^�q5X��X�<�c&j��b�Y-ʍ"HG�]�7�WR/s��S�>ȅ߻�7M���6�p�@�>���d!�[������Hi��Fa���繑����U����;�T-������z,n���ߋz^��P����g�[�<9��0K��[�P�b���\j�q�O��	�c�a�]~�)z�~�q?R�*�O��*�P�v�Zͮe��R��z�%��7?�i�!�a.���O�]�y�����p�?����ͽo��^a���
�ş��{]&a���ɇ��^c?3L�����ܞ�C�5�U�ר�zF��z��k����)+��9���8 ��FB�m����U4&� �'��F�_|��SQ�l��A����Qܜ�\�8�����\X^���y.����De*$�h�����sɯX���lj��U*��9F��?o|�Q>/�`L�<�d�zN����}�E���s\�%�5����Ι���{~�d͞o�u!����Ş, @p�<�\�*�@��V3��7:����A�:��[���WI�����q�XT�_ �phg��}A�勢L)܇p�,��W��
{��X�)�*��u-,7��^��*W=Xz�U=�!��Baa��Z���3Y�����#�: @"�/*��e��s��~uK?���Z�����*2o-̍�����a�����'~�<?-��/k]��� �����
�;��!��N��[/�F����P H,���Х��9ao6��?�%5N\�]�5S ����Bm�a��i��ד��	�F�~��r=Vn�b�q(��H���|Q�%�K��É��n�\ʭ7>��gB  �
����Z7��Z��HX��}��6Ȁ�XX��-E�+��綰a�/�os&�x�S���(ʌj�Z�y�6�Ν_n���s-��E����r���P H$�s�����\�j����σ��\n�Ͻ��+��޲��\�
��_�����J��T�]����.���	jq�(�\NT���-�s�틋���R6�\ʍ[�Q*tB� $�r�D�f��ׅ�"���x��v���ܼ>y�߰��9Uf�\�P�ϛWX��w[F��s=�R��"4>H���'�Q�����!�_�ޯ,�K���:w)�r��R�Nu �D����Ԟ,~>��G�c�sH�z�
;~���h��}��\��y.X�\5�t�~��9�z˂|�(�P\��_E�m�P��ԝ�!��\ʭ�ߣb�Nu  Ĝ��V�e��>�x�r��;������[#���}��|(势O?�0_�\�$�)Q�?dY_~�B��~�iX[�P.�&�r�Nu!�>uڣ��6o�L]��OOO�xܺu묵��  ,n���?o�u7��,�^����-����(S#̇J�x�\�<�2��0.|�s�2���Z�F���+:!ԅh�@�����Y�k� �M����Q������Q�r�J�
�5쵪u���C�h�W��e��\ʍ�R��   Q5�)�r��@'�: !�Y�y�k�R��L��Kg���R���oO*e7   ��@'�: �\��L�ؼ�}���9t��ж�����iG.��J�]n   H�r��R��Oe��?�{���N��=8m�7���u����R�=�;  ���$�	����/�H6��3����qc�}�;�]��i@ >�y���͵س�Vʥ\ʭ�ܨ|�חr�ܰT�!B��А�>}�&e]u�U�?oܸ�ZZZܶH��A{{������Yss0�F٬�0ה�����-H�v���Z{�@����p�i@k�N����ǼW�}��C��K�+��܇>o�����[�Q�U�!B]T�����.yִ��ի�=nvv�2�L��)Ѝ�gz��e��U��7w�o���9� �  �C��Nu!���6�z��������B�̴��^�e���u����|��^���H�  �� ��6B��ު��A��C�͡Ӑ�0{�
)ح�������3   D"�@'�VBD%c!̡+��bvܿo���b�!�AI�Rn�1�R.�_nT2���[G�!�@'�v�m[p�����*t.���9��0L�D�Kgf�mbb�����͛��ň(�r)7�r������:*7hA:��Pw�С�ܷTP������fK�̀�L�gz#} �vg��ەJ�6`�$���٭[�R�T+Ɩ�G�r)�r�/7*)^_ʭ�r�F���u@�e��}m���>v���KoJQ���?��K��[�r����K�uTn��
t��w��dR�~��~cnJT�� ��R.�Rn�����K�uTn��t��w ��*���Kg�[2iBJ�?�'O�����ߺ��@��R.�Rnr�mM���[G�+�@'�}w �*k#Z}���}#�D9���sDK�t4��
�K���\S���[G喪�Nu@�e�V�-V�����   ��U�BPc�tf�bFA3E�  D-��      �tB�jl|.~�/�{����   *E�B     �@'�:���4۶q��
��L���  �"�   @��s�b1�K�l�   �u@��2@���   �H�:��b���ۖ�X�e���U�V�t�5k(�r)7F�F��חr�ܸ!�5�2�\{ߎ3�ܽ�b�9��5���x��u���i�\ʥ܈ˍ�^_ʭ�r�PD �uA*�.�׀���͛˾][[��^�Rʥ\ʭ�ܨ�����:*7�u@R)��mg_���݃Q>�u�����ЀT�ԫ�)�R.�V_nT���Rn�g�: "mM��i�p~�ξ�T*�׀�R����z����P.�Rn��F%��K�uTnꀈ�ޗ�G9���9��^:�"�N[ss��:u�r)�rVnTҼ��[G�&��P������L|c��,Wa2�vP�l6k333�K����r������:*7	u@��S�<�}=�o�p-���L�L   �B�T�n�hJ�� �)�5g��  ��: |��{��7���r�:  @}!�1�`�^�u�}k�؃_nUʝ}]��0�+:�n�=���/{̧:˟�>4�bώwX5(�r)��r����~�ߣ��Q/Z*���oߎ�Tf��7wTsn��t���H��K�	-7*���K�uTn��v͖�Y.��<k���y�_�|;mj��Դ#w�   ���1�����w6��Y��X*3�I�`�q�lӶ\�붬�h��~   @c �	�^���nwޕ!.e   h0��inS���    
e����&ԕ!�B�pvh    �IY(�R��PW����S��3    �3���GU6��c����}�y3    GC/'�����Dط{8�{��T���     G�GY>��Lc};�hch��   Ț�Ӣ�Q>B]F�3=M��   иr���o���� �Ub���ѝ}
v���   ����.�Nu�R�3�Yw߷v�RYO   @.���Lo�C.��4�����ξ�uM�#e���   P?�r�2��曻�[���kQ�f핹    IEND�B`�PK
     $s�[$7h�!  �!  /   images/a7fde0f7-2836-4f0c-aad0-66dcccec46ff.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     $s�[��n GV GV /   images/5a738b76-89aa-4728-b8e5-f09c859dbb14.png�PNG

   IHDR  �  "   �?��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���|w���������j�dɲ,˽�v�$!q��;:� �H.wGr$��B�����s)$�@(C��;.�w˖l�����&�Ųg������gƊ�7kiFZ�|������LB                 d�]                 � �                ��@�                ��                rw                @N �                �	�                9��;                 'p                ��                ��@�                ��                rw                @N �                �	�                9��;                 'pϲ�Sgj�vړ�&���{�����4��oxL���E               ��s9l��n�ץ|�C�M���>'����"�Dc�h`$�a��	!�����"�^՗jz�PUE>�#���B��������7���aI.ۺ����_{���w($               `���/�kz�@5e���nE�/���8�?2�=8����ݎޑ��j�$��&�Mf�-5�j�-֜䲱�/��a�~v�����2��֖=�z�[;���               �Dg4�6��sj�S���ӊT�e_����0�����}ښ���h���T'���	2:�7V��tf��55;y�oWv��\Z�\��P$�W�Ն7�j����               �(�|��Ơ�5�k�2x�Y}=F��Y�E�q��7?ftvqg�6�qD��w+�A�� �~��:��Jo[P��"�r��a��Ը�]���~��~��ں�               �#ľ��\�ϩ���rٲ݅�/�,H��:u���"z~{{*�k�	�;��P���;���u�*��DU[V��i�fm;أ�lث�li�X8&                [�������u�P{�g���<�Cg/�I���~��~���T�j�y܏���]��A+�+e��gɟ0{ZQj|��yzr�A���]j뢫;               2'��҅�R����ݚL
}.]rrcjl�߭G^ح��R,��/���c?mN��&���&;�ۡ�'���e�S�!<��.m��%                ]j�
t��3���5rح�����Ƒ�=��.���}G��A��X-��R���E�J�4����+S�xB�_�ܦM{;               ���4_�9�IgͯI5��j�~�>~�<��Yz��z�]��ϊY���-�++�|B�+9U/�qD��|��t�               8^�]vv�޶`j��P�ש�٬w-��������{�'4�pO2:���y:if��-kjɌ2�j�A���f��               +�ݪ�V��{Ϙ%���*�w��w-Ѕ�g�'^�;:4UM���鲷�$��x�ϲZ,:{AM�����E�oث��~8               ��ȟ^w��z�?�h�}��W�����oT�����)p�_W�.\���A�c��v�,�����ˏ����               �����Gϙ�j���Y�\�Ee��u��g�P|
u��rw�Ӯ�ϛ�s�	�oNm������Γ[��s���              ��9}N�>q�x���q;m��s���\�{�%��T0��M��|�RUӵ�N�M;g��7U$O��               �.�æ��>G�h�1��D߾�,}���䦃��D��b�.Y٨��1Gv�E0���R�w�Y�����Ү#              ��3=X��w/Wu	ͨ��s;tӥK���L_{|��&�Ip�8�q�"�1�ZH�B�K������3;��_lU<�               ��U�uㅋ�vڄ�9gq�+���|A�#��&u��<���_���!��N�}�LU�鮇6h,<y�              �d�Xt�;��ғ�̘Q�׷>v�>���ڸ�S�ͤ�Ϫ.���[�@�KȬSfW��W�����9u�
               ���a�?\�Xg̭2�����?x����+�ū4�Lʀ��͕�ǵK�r0�A�ԗ꟯<]7��s�t@               �<�>��x��TSjd��f��_�D����ׯk��t�3�M�'/Y"��"dW���?_a�ܟ��{              ���(߭/~�Օ�e�H<�Y�<����M�'��&U���%u��ꅲZr?�>4I��;24���{b1�`4�*֙�[{��j���[��-�|��Z���k�y�������v��|�C���)��ߞՖ��              ��e4@��GNUE��\���50����	�ĎF��X<�O$�c�x_"a�U"^�t�J���mV[�Ӯ"��Y��9+�
�~�˪w��z٭V}��W'|�}�܍o�u�/P.f���Q�92���;��p�H�w]{����ښ����v���@��꒼y��y�ֽ����<E��g�              LPF���.?Me�e.:�=j���=0���ѱ_������GN��w?:��?3��:���s��`ae�י[�ݤs���f��?|I9�>)��XT�kϟ�S���]�c{����	=��}׌����Z���so�ۍ��|��*<��U���k���s�Ż�iӝ8Y7~�)�<�'               L%}�ç�T�}$M�~�g���������������|��&�{k�u�:{�՞��|���N�Q^Phɑ �;�h4��ߤ�j��O�S��,V.4-��7��ڲ����_������k��w�'��0N��k+��5O+��rز�U2:��'���<��G              ��W�s�:YU�y�~)�'��m�ݻ;�w`���Z�ӕ��кjU4���[C��?��$�w[Su��r�ש,�py��"1���-��&t�}nm�>yq�����z{�'�?�v(r׃�k��o�<_5���?8�wͫ/~oe�����w�V��{���1               w96����-+���	�_z�ȓG�F�.]�ڏW���\�=��͇/����2zi�5�]���ԙ��գ/��D3a�E>}��S'M�lo���v�����r���qw^��HrqY�uW:7��ܚ��낅�l���߫;޿R��)���              @�1��7^�Hsj�������v�����|���wk�֏_���������O�-��������;_}�|��s��k"���|�C����*�R�-��;^?��mW�~P�[]�oimM|zcՏn]�P������L���J�n�t�n���H      &0z�x�	y�q��	���.krݦ�H���O}�1+����vKBV�  8nƵ�p���蛿n�K�B�aU8&�Ƭ���,�u��"�Ԕ�      �M>k�Κ?-+���m�u�?��?�z��!M0w\s�S�ł�o>�����;Kggg���q?���^w�o���_ń��؛�_�⼌ﻳ4����w�r��VMp���;��������+=�zZK�{�.{FϚ��z����      �ƪ�
�	�b*�Ǖ���Hȗ\7�5{3] 0nF�}4j�pĢ!c�����V����&��     �-+�+���ge|��xB/�hߴ�;|�;��&�֏_�Br�r�=�����냅��ܿ�i���[��~��	k"�p��٬�f�gt��x\vtlڹ��_����jy����o����8�6�Ȣ��zK��`���ơ>���!      �>�5�wLW\~gL���#� �4ޜ}$�R�b���F,�[���7����B�      H���<}�%�p�q�?:8�򮎫?}�E��$s�G/�Akk��u?��)�+/��82v�+���Sk���{fB̨8��g��g4et�:G��Кۯ�������%�%���#7��Ss{�ϙ�����o� ��O�k`L      SY�=�2OTE��J=��2&�� ��+�|�1���Q�z�6��sԦ��z,.      ��鰩�=��se.f�ƴn�����׭��I{�筿�U7}���Λ^��9�%�L���a�թ3�_O�T��0�|�C7�Y�
Dg�˻��ٴ�{�WoXۣ)����u��xlac����L�����k����<�xb<     `�cm�7�
cxbrڸ6 �_�'Te����f�=���sԪ��'���]<"     pܮ8�EӃ�_��h����W�z���q׵�lomMT�}���V�q�2����ok�ƽ]z�`nG�'L���ՋTV��ȾFB�ĺ����_p�����[�-yҔ�y��Us����C��Jt��3��3o     `��Z��'�
�Wzc*t�  N�͒Py���1*����wa��Q�B1��      ����fŌ��o���/�?���׼w������_t�}�����U�)-�8ҽO�բ�/]�������V�������9U�WG�p���G�q�ի�i
{�9���~�w,���㴧���eok�;:t�sP      ��E	���ɋhzAT.뤝U ���'�PI�D�7qרU���7��aw     �?����/Z��EV<�Я7|���w���ۮ\��#_����/Ϭ
ҽ��"�.;�E�x|�rU��}.}��y�����#�nm[jt0Rn�|�]�{9�΅5�+�:�:���nM�`\����m�     �Detj7����EU��i�Z  ِz��K�E%!���t`ȡ�a:�     ��+�1W%��'��|�>t��Bʗ�]����jFñm�LK��V�T��lnӖ���E9p��y*�:Ӿ���z{_��?����~�g?��?��x�����O�޴N�<�H$O�G_�-     ����WCA89�r��� @.�*�*o45�	���ƀS#F��     `j�=�H�-�K�~��Q��}��rŚ�
����C��>0#�5z������ܗ�b��^�HW��+E��wO+���t漴?��M{��v�u6ߑ<0�?�k.~*q�#�N�]�|uI^Z�1�=0�
�	      �٬R�7�Ƃ�ʽ���׭�n������~v�M��^O~�� ��y5�����n�XF����y��Z�͋��pԪ}�v��w��     ��բ�]�(zN���p◯��ȧ?zѿ
ԃ�k�J-���'�>}N�)��WMi�.Z1C?xz�rM�܍i�?~�ܴ�g{[oϮ��-��n�K�z�ƛ����3L�T�O_[}�ˮ��6[_y�U     �<G\�
ê/��iͽP�Vw�\�x<�3�n9���p8�a�[,D� '��G"��cccM�����rddD�P�5����j	����mخ�}.�	     `�8Y���
Һ�p4�'_;x��csͻ�9��~����%����Θ�'7P���rI��ߵ�^��i��ގ��W�zg�y����u�%�w?�γW=�������%uz|�^�<�'     �\R슩�V]^$դ!ی�yyy���W�ϧ��2?�g�;��� �{l6[j���?�D"tJ�Ac98����Tg�l2~���ES�g̪��N�t(�\&     `��8�U�Һ�h<�������+�|S8f��>�eǯw,�Q6#]�����Y���G_Q.�ɀ��i��jN�>����zx�>���0.�]�z�힇���%���<��rUט��#oo�?|�Y     d�q�&/���Z�e�u����B��#� ��d L Ƭ!>�/5����>�������7G��z/rǵ�=�E�T����"q��     `�y�iM*���V߸�����+�|F��VK��{<�����<��4]�y��Z=��.�;�;��s2�~�I��d�����/|b��|����r�#��W4|ޚ�)���jnm�6��     @v$T�iAј���N����U\T$�ߟ��n�� L>�;�^UU��X,S����z{��ӣ��0>�I^GB�JB�����t     �GQ�[.oH�>~����7]v��q���G
���9�}_]Y�'�0r�F�۾��rE��=N�֞:3m�㉄�m9𩻮�d�pBn�j����w�>�zU��atq���O	      ����/
�ȕ� �ѡ=�����D%�ũn�  LU��Ţ@ 5���Sݾ��ݭ�.���f�ûӖм����°vt     �ĻO�)�Ö����t��qι�	���]t�{�c�z�u��rQ괖jͨة]�}�9p_��A�^g��?���3�\��.�]�oo�=2�:P���skK4��D��u	      ��Q-(	)��L���p���Le��*M�=�.� ��.���_�h��W$QWW��vv�ȑ#�F�i����3#�����~��	     L8�<�޵tz��w��6�m?�VK�ȝ�n�z�:����[:��t�7&~�M���F��[�[�:�����/��8[0M�Uћ����A�gs �mM�>.=���;     H�GL�KC��{���n�A�'GQQQ*�  ��xH���"5b�:;�q�HF��n[\KJ�4� �M=.�r     `"��9�Խ=O���_w�5�S0�'/�����~�����g���)�+UU��C�Cʶ�
��9�Z�����$^|���~xL0�]׭�����.\���t܌]�T���|�     �ٜF'�@HM��,J_V�՚
�WUV�:�j �<��~�#n�ݻ�t���T���s�8�:�|T3G#z�˭�PZz     ��i���e������CO�z���L�vp��꒡���<��V�E�h��ߤl˩��%'7���s�ۿ���Y��^��������JM��g��5���<��      �bUB́��BrX�l���Ju���s�r  ���PYYYYj�B!�wt�P[��ҶϠ'�s�iπC�t��t     ���5*���R��k0�y0�ZH�����}���n�,�}3͔�Y\���j�G#ʦ����RS���´��tp����j�������\v�Ϙ3�U�'^�H(�S�    �ɯ����2� �h�^W���< ��p�\���M���~8xP�JKWw��HCADվ�6v��ƀ㭏     ��է�n"��K��n��F�����ߚ�ȯnX<�l�ٵ]��6�F���[ٔ3��g��x�dyew���iu��\���������]��댹���K�     p��ք�B���"��|>��֦:�ӭ ��RXX���1��Qm�i���3}?.[B'���.?�;=���     䎙�~5&G:���s�-�_�U!�v�=7�}�Q�u��a��tpO��:cNUZj���c�W��!#��=���ʁ���
<f�>oIw     pܪ�ZZ2*���`{iI����U\\,  �ی������L+G�h���4}?AOL�N��^���8��;     ��jH=�&v�PȈ�?z���=��w,�}�ٵ��<�H��Q��D��Ԗ�TK{��#1�=2�>!c�N����ue�6����"Ք��@���    ���&��$��s'��X,*+-UCC����t:  �c�ZUYQ�]��ڹs����L݇͒Ђ�1��E�L�[}a��     +�բ��Ԑz���uw��E[��Y�w�C�_R�9̮}��i��u�����;�^�QȨ[�Xݺ�W��X[��3��i�c�?�m     ��(q�trpT���i5�`{Ey�f̘���< �����X%+V���v�RO��7��ΘΙ6�W�]��g�o��;     ȼ%�A�{���	E���.2�hJ}R�O�_���ڧ�T�?٤��#����=-j(3�n4W[��Ǆ��r��[�e�7�]��9��    �_dUBs���w���577+??_  `�Iݓ���رC�����6��/)S�7��z4%�     2봖�4�~e���_�v�^!�v��?���ݥ�S3�E�nͭ+զ��ʆ��W6W�n��^w�Ν�W^������?y���k���\f֝,PuI�ں�     ��8�:58��˼��~�_���TTT$  0�!��+��ѡ;wjddĴ�ިΫ�sn���:     0Eج�Tf�l�hL����⾫����?z���K̮}jK���/k�^3�Hh�ၿ�f�ZK����W�>�q�p     L�/���Q9��tm��|�5k��e��@  r��bQEE����<�7v�R86���ת�Qm�uhc�K	��     ���i���8L����[��K^��`��U����=NS;��#�}��p�Z��3̿9������/���UG�oG?�q�M�*�$y�����     �o%4�(�yEF�����6�U���jhh��j��  `�0���֪��2r߿��҉K�%V�;��;<��     �ϲ��	+����U_�amO�COn>�)8�̺U�y�,��pϰ2-����� N��������u_��=]syrϒ�3�.�^*�æp$&      ���*��s����>{�ly<  �7�á��ͪ����m����kJݠ'�s������l     H��i��}�{(�ُ��!�u|U
~���f���2ߔ:����KL�i��;�?%䄃�C�,����5]��*�ڼ�[     `j+v�tz���������2{�JJ̿f  &����X�\Ԏ;�DN��/�^��U�Z�����
     S���PC�������Z�	����-��*>S;�ϫ+�z���b�k�~����׼w��⍅��50�����-G�&O�     Lm��:�lD6�	��MKud���
  ����!j�֭���8�zV���lTgL/w�u��     �i���Ե3�	����3v����2�;�̚sk��z���-�7O�<:�_B�h]�*z��x�����̺-5�;     `��kqɘN�Z���ռ�sUTĵ  0~N�S�.T{{��nۦp8|�5��9^{\��*     �	KGC���w]s�z!gt�ޞ\�p/�w�"�S{�2)k���<xM킟z�{$�-!�t��(�05��\�Mg     �"��Ȓ�1�,<��]� �Y***T\\lZ7����|�a��ݫѨ���     ��3�:`z�C]/9�k.~�̧�G��^��u��M��{Cy��5v�|�ڵ{��2*�}�x�6�Մ���R�s������1    ���nM��QUz�'T��vk��*
�1  L]��ͽ��-��=��P�bWL�֯y51�     �zґ���<(�}��{���&3k�'��_�vP����{}:��C[��s���,��3����f֭/��k�Ļ�     ���&��bD�����4w�<9�6�   ����j��q�N����ۍ��a�zC��    ��z�*�w�Zs,U<�!�t��>�\�p/P�e-�>=h�_���'BNj���P^x��5��Ћ;	�    0�����FR]L���bь�566
   �|>�V�X��;vh߾}'T�mK��a�;�U�M      㑎��{�t�^�vH�9�C�{���ƽ1�L��%Y�W�Z/���X��m!'�FO.L�W�|    ����S�v�3~�5�^�.X����_|  S��j���f�~m޲E�h��k����o;�j!�     �ݴ�|�k���*��^{��S�Z�x�f�,-���)9����#k���gj�����;�����##�6�fy�+     0y�9�:�jD>��ۋ-\�P.�K   �PQQ�������>�:vkB�*���G���v�     L0�4d-��"/9�k`��"�0���>���@�2%+W�y.���v���r���^�lJ�6��<(���     �>{Bo;�p��i��2{v�{*  @6��|Z�b�^ݸQ]]]�]�jI���=��U!w     pґ��<#䬁����´���"yM�������Ccto�a�����Ӟ�)�7�Q�2�WV�E�DB     `�p��:�rDy�n7�F���  �
�á�K�h�Νڽg�qױZ�S�G��ݫ�sJ    ��'X�1�^,���J�Y��m��r3k�3)+w���)����;���=8�US�_cV=��"�ۡ�Ѱ     ����uvը
��n7�cK/V   @��X,jjj���Ֆ�[�8�&>6KB�ʇ���^��;     �ӊ�ݦ�����^�vH�Y�c����̬��3?���d�W��az͑Pl����G�{���B���;     ��Ӛ�Y�#�nw�\Z�t����  �ˌ�f<�^y�UE���a�JgT���C^u���     ��<���ݞ�P����:�kx�ʤ��������~!�E"�n�k�Nӫ    �LKu!�Q�����F�}�%r���B  �.%%%:i�2mx�%������a< X5������
     ��۬�������Bnk�1f4f4K:��NV�y�;�+�.!�E�	ӟ�1��"     �yƥ����*uǎk��߯�K����:  �X
�r�
��a�FFF���1Ϊ���ͫ�!w     �?|.�L�8����㻈��i]�*z�+n�ʹ�~Z��FV��!fKX�BNK(nz��ag�M     &��%c�ɋ׶eeeZ�p��V�\  `b�z�Z�|�^X�^����U#�ת�Q��ͫh���     `�r:��X��㻀��EL�;���攕��#���G����z̮�s�    ����֬�8�� �d�r�R!��/�������ө��m�W�      Ғ׍��CB�E�Fw)�Y�2ݐ:;w�CɉDB;��v
9-�v�]�I�    �	�6/�E%cǵ-�v  0�8�N��l�	�ܫ�Q-)ӋG�     ��!�����
�L�g��\V��ۦ�hBѢK�
9-;����&�    `b�;cZQ6z\�������y�� �I��/?�$��a�������̂�zǬzc����     `��X�OY&d�	9/��ͬ��c���J�=3�k&k�6�{�$�zT�Y���욑sl    0Ѹl	�^1*�u����Z0~�/�  d����ҥK�~����侴,���MGG3;u4     �-1s3�)6�
���v�f֋D3�\CV�ј�'��/��f�)w�%     �>F,}epT��������X, �  &=�áeK������踷�*�S�#z�ͧ�(��     0U���g,�6K���\���h���������i)r��j�]3�O�     �3�8�*ot��j�E�Z	h ����r�e���/(
�{{�=���G��C^�<     �T�����n#�>x�vSo���a�?'+����ob�%q��T�iv�������     H�i���������j��Ų۳r)   k��AF'�֯W$��%�����-     0����z�_b�Y�BNkmMX��ͦv<e6������#㿑��8�r!�9l��F�?�     �����V��&�����\����RK  ��(???5���_T"1��R�&X�cv��      S��u;��尙V�e����	>^a�ԙZs`d�3��,���K���BN��8�̮�74&     �ی�+�F崍/�e��Ra.����  `j+**�ܹs��k���+JG��P�F"�6�     �є���cZ=��H�i6K�4�k�d�!uV���K�������L�O$4���3     ��Z!�{c���b��B\~�_   ����448�={��{[�-����z�ͣ��    0���L��^w�u��U��BN�l+̮�?�G�GM�Y�uLrZ�ߛgf���1��㟊     dN�;�y�����بʊ
  �̚5K���:r�踷��j	����%     0ut����Ҽ�BN�Mz�Yr�9!'�sͮy�oD����{W�����V�:D�zB��Խ�o(�:Mm	��;,     ���քN	�ʪ�=�^YY���z  ���?�^X�^���x�}Į�M     `jHG��fM�.�9���nv͎�)p7�nI��"�i5K�ߍֻ�k�z퐐s���f����     �gAQH���������ܹse����<  ��a�۵x�"=�쳊D"���x�pEpL?=���    05t���v�˵T�Y��R�kf�)uV��=C��mV�������9'�k��5���    �\U⎩�?����Z�p�lV�   �y<͛7O�����%��ΘZ�!m�u	     L~����Z�9��{VQY��Ys`$������;QY���ВASk�;/��TU����{:�     r�ՒЊ�QY4��U��٩�   �˂ee���վ}�ƽ�ܢ����	     Ln{�����V��&�����M勴�XCW�Mn&���n���8a�~�"!�|��_�u�����=2      �{��U���̚�UUU	   �nVS����ԛ�a�H+����6��     L^G�GRݷ���jx��h��$WrJi��<�kN������l����'��x�sW��3��?�q�M�::�����i3     ��	8c��k����nn   ��j�j�z�g��o��wLM����9     &�D�ͦ�sk��S\��_�sNU����{�f�!u����'K(��a�ԇ�d-�#rYr��B�()�\bv͝�{O�o�s     �~K�B�����n���ϛ�Z  `�<nw�a�M��6�m���Ю���     ��v���p�(�rʧ�y���4�cv]��ɴ�ܣ����:sO���C"��S����Cl�.    ��R�Q��6������   �_UU��vv���}\�9�	-(������     9d�]r��5gV��o���i_��BN�{=�X-Sk��� 2-kw���ݦ�[j�[Z��ӂ����|?|������5%�?�%y�     ��a�$��$4�m~��O   N\������Q(4��d���w�;dެ�      �l�o~Sa�æ
��3��˄��P^x��5��V��'o6MV��R��8-������O
YWQ���f�4N�m{     r��@X>{��?�f�j������E  `�r:���Ң�_ye\��Ɩ���gm޷�     &�ޡ�u��8�Ժ�kD�='����S�
ͮ�y��G���7�9�p4.��jj��҂���{ֵ�[gov�-2����     ��#�f��:�655���
   �	��������qmW�iz^D{��     ��K���p�Q^���o<|��\���U%�����X�7�(�p7���vjic�Ժ��*[�����+/�)d�}���/+1}>�Y:Y     ���hL�q�/���Wmm�   `���fuvu)_����!�v(���;     �ы;�h�I���4��E�O'W����5am�^��u��C��ޯl�j����GL�;lV���O��.dMS��o�Qw�.�     �BgLu��O͙3G��    ��r���Q۶m�vƬ<3"��Ow     &��{�*��aGעc��>x��_y��7����U��;��f�5R�	eC���l;���3Of��\�Pv�w?:�+W_xPȸ��{�YՁ"��v��C}     �aAQH㹬SSS���/   �O]m�>�����S�[֮��tq    `�����#Z�Taj�B��Z]�wOru��sj��IG�g_oW�d=�~�oD��z�<��,��e�����&W�2�����t����CY{     ��bWL��b���N�C3  ��k�=[�=��㸯����hk/]�    ��~����wâ���Z�~ ���CBF}��Gn��̮;�j��)p7�fK��w���w������7��KȘ[�}�Җ��`:j���&     �����=��TӬYr:	K  dBaa����t�m|�VZ�T�P�.�     L6Ͼ~X�h\N��Ժ%����Zr�2!��Ԕܘ���ooO+ْw�+�U�'����
�NkMy���w	�\U�5������{���P�     @���c��F���}>_*`  �̙9s���+Ǭ;ք�
�z��%     0�]�_�Ѯ�Z̿g�xF��Z����ׯ�2���������t���k�mH��΁Qmx�C'�,7��ɳ+�k��ѕ�W^���v��2����od�/��8f�     i4'��7Ϛ�t<  �?��ri���ڵk׸���k[�S���     �l�xi_ZGI�����*!�Z�~ oYc����=8��ugSN�?ٰ/-w�æ�?H�N����<P����5�c�~��    ��+p�U�;���EEE*++   2�~�t<xP�б?�htq�Q��~�     ���Ү�:�7���kz핳*��������/���VŁ��*޴\�1�0r�ٔ3wcʃ��Q�xL�=�����o?��[/_}��6��Oण����     d_�?�c��itmojj   ��n����A۶m�v́�v8gv]     &�x"�'^ާ�5����Ms���_r�TH�۾���+�+�LG�����>e[�܍��c���#g�������[������k{�Oܬ�Y~Z��?�����     ���U�9��7:��~   {j�MӾ}�422r����qMK���?���F      �߰W�9�IN���ڳk�J�����r��� �ESM��v�w��^oWG�_CJ��	�~�����&y�濬��1�6�lr�Y0U��~Z����H:~�v�զ��     �7�0,���?FC�   �]V�UӧO�֭[ǵݜ@X���v�:     �z�B����$ga��TU��yf�vWie!��tD�!�lc����}��w��x�À�H��L0>��AY"!$��rZI�����U�uuO�TW�U�V������SM����ݳ�����y���ޏ7���)�������憛��+�i(��?���F���7��,Z��
��%����}xӅ�1>_z�ة����>��?z��@ƺ1�W���;�����Uk�a!�B!�B�:V���>�����!����B!��<�6n�޽{�J����17p,ٜ�#B!�B!��V6�u�m��4���]��r���o�s�c{��r�!|��o���]�ڬ���$�?�V���V����ۆp(@X ^}֖�&����x�[R7���?{�i�w7������!�B!�BV�-�YDTS��;v�B!�����[��SOz܎�,�B!�BHr��<~��!\�{cS��Xo�ቅ�����G�����O�Z$�<��_~�$Z����N�����+.<�)�k��v��������WN���Ǯ��+/?c�����'���9!�B!�B�ǎތ���}}��!�Bi6oތ��?�LF��nKW���"�7�͍B!�B!+�W�.ݵ�)-����O~�����ǿ��={Lu�������4�5�80�{�=�V���_��Sxݹ[mҧ6u�/<e��w����y��}I���S/9cӏ:�����/���!�B!�BV������!}����A!�BZMӰu�<��ҏQۺ�xj�i�)!�B!�BV�bN�^qFsZ�E�k������w�/����Ajb��[�:s����OZ�K�=�V�%�s)�t�^���On�k��y`d!�}l���={yw��#�ݲ�=4� ���8���B!�BH+pro6�U��靝�!�Bi=�����a��c;{2xj:��ŝB!�Bi7����q����My~����gm�6��7���\yH ���?���]�/h�k<��8z~�DK�-�v�Sx�ٛ1�k�k��st{&wۯ�×�H���n�8sS��-#��|�ʯ�>B!�B!��<�b⤞���Vh�B!��&�Hc��8|Dއ��8�l�ݗ	!�B!��r�\���~�wi�J���a���m��r����o�D����͟�|�Ʒ4�5���A�Ѳ�d&W����7���׹��u���~�����=�'V���뻞>}��P3_G��i��~B!�B!��;s��r�횪b� �B!�˖-[�-N��2�N!�B!��)_���x�Y�1��Rꡞ���]n�?�p����'@<�䗾��ל������;�}���x��,Z���[���~���m8}�@S_�glz�5߼������u�:H��M#/����i����Z߹{/�o�?,�B!�B�Zek�|{����A!�BZ���~���bffF�1�:��W�Z�!�B!��^,���¿?�?�yM}��C]�W���a�s�zͧ?��A�|��?��Ugn~��67�>��ƿ��I�"-p7L���|�W"R��Z/ߵ�������_w�K���I����u��~�I#m��n�k�N�+?�s!�B!��V!��X�)��e�fB!���gs����G�>?��X��P���EB!�B!���m��+�܄�w�6�u��;�o8�O#�~����o�7�
��_t�8s㛚��nq��l"�V�����s��O�_qZ�_��#'E��w����Co?��y�����-?]��Y�����=�d&B!�B!��VS����t������韏'�B!`���x�q�!�����B!�B!��?|�!|��F,�5�u�:����;�ڵ������s س�T���ދN]w�r��=���9�VeU(P_��i\|�zl�m�k��28��>�^���~��o��0����>|��G�[��ȏx�={�B!�Bi�t�}Æ �B!��P(���Q>rD�1~�B7�� F!�B!�����T���(>��g5��:�!�?^��:���W�?��+��Q�?��f���M'���;O۴nx9^o.�-R�2�"������õ�{"��g�7�D�����C_��������Xc�sϗc�2v��wm�l9nq`qxr���# �B!�BH�QM�������@!�BV�������9�_�B!�B!����y��Ņ��k�k�4�={��<6��C�|�=��k��_{ӻ.ݵ��=�e�t���a|&�VfU�-���u�X�
9sY^/֔ן�������k{n�e���7��ϯ��������z��5u��'�uiyÜB!�B!�gCG��g߇����@!�BV�5\4E:��~��.�wB!�B!��1M�o�� ����@��x?�����w<���������:���1վ�?��36�)�6����-���9�Vg��-�w�^��u��޸l�y�6u���M��ػ���Ц�����g�l��y;���#Z��JZ\x��$!��V��YLwT��vɏ;�*4�D<\�p�,zw�)D��;#�J~��B�z~/��Rƨ�H���J���
���T~�0̧��q"k"�3A!��6t���_B!���P�p�}��I?fCg��DE�B!�Bi_f|������D��^�z�7^����n}��ǒ��7x�a�)����{ֶ_]����|��������Up�>�Ė�l]��q��u�����������ؾ�o�����m�_\��w�����z;����O�|���@!�ԋL�pzwDAGȺ#���j ��)4E�f�����0��>��f����T�@)\���+ӥ��Y瓕W�R}�4����gߕ��fB����
�k��f,>G8����P!��B�Aՠ����o��5dMYCA*��uV@>mb6�ͤudx3B!��P�W5�;�.TU���(!�B��c��u��Q��@L�DJ!�BH;�)
zb
b!a� +� �Z�f� +�X��eW��g@-�^�뭔����gК3ET-q�j�P��3U~�0����P�-�l~�[�2Yʳ���n(Hdd�ߚU�5�2���x"!���<��8�t�c�ϯٽl���߃/>m�٧oJ���9����=��6��|wө��/8uݙ���]�H�s��7�Ar��VU�����Z?��s9:c�{���[Gw�������ѭ����g���Ǳ����ι;7u�#�,������} �B����J_\�`\A_�j&:4QE�j�Fz�L
�\�T� �(�%�_����f�5���tyV
����Z��i,/����� �(Ў����k-KJq�t�W��mk��\����f��������3��o.>W؄2��H!,�E�0�H!�15$ti]�t
�H���A7����B!��P�@D�3�
�:��B!�����G4E:��~̆��Bi)�2��}q�!a�k��������/�Ӻer.�_z.�l��2��`)���7"Y|��Oh)f����A0]��y+5z�&
6�U�ee�#f�T�0�P�P�e9���"gj�ME&��TNE"�gML%ML&�	B�Z盿|�n�%�/�|��b������F�֏^���|⪷܈U�;�|9v���/:u�]}�Qˌu������9�V��h��?q�}��;^V���r����37�fvg��o���}'����\�V{��݋���?���3#��g����~�TF�V�B�M11��o
�"@WHGT�A320s��z:��aŐz��������Ei�ƪ�����=��1.�܎�Uӂ9ט�C��ޝ�v�q�}�q���o����X~�o��m�jB�U�E�D�����2f9�'�7���A!��V6tȷ7����B!��^���q��A��;�<2!�BH3��������S�1�X1EG9(��z�t�t
��%_1��Z*���j���*K�*�n����|y(�k�p�$
��sn�Y�y=��L*Yy�Y슏���ͣ-?p�,d��,ܽ1��B�
�`���-op.�ê7���7H!��v��o݇��/-ݗ�S7��o���;&a��y�[���=�������go~�X_Gd�����1����&Ve����g����>x�9+��=���/K�s{�~��w:>��O��O�����7�~���:���!u�? R&������&�A!�=�*��c5���3�bj!33���I"�J��SjQ\RX�P��uk�D��t���qI(�;�����\y�q\>�8���w� �`��8�;+� �^5���t2��2�(?�
Z��b��n�X�_�B�!��0�u�I�Ь��d��E�Bi;�u�ܭ��	!�BV5���cVa����r~!�BV7a�q��x'���3d��a�*�JCϦ�XX(��+P�-Y��;7g�
1���
���Y����qŜ`M�B,ۚ�o�Q�U�o���\�l�2o�5:�uX�`���c&"=D���ݢu-V§�׌�i��M�ӑ�=H!�+�i_���1�ױ"��b���]����O�����˛�-̇>s������9g���c+z���b����j��}��o���:�!�]/Νf<��柏�=2�oG&�?�>�Sh>z��F;��r�H�[G{zW����о������B�������jAp�	�Ur����$���ֺ�Y����%��P��s��֪�ν[���<��׸�h�b�c��`�m�)\��c�\�����¼�h%r7���������x��Z%�kC�D�+�H�j8��ł��������!!��DTQ����tw#��B!��^���
͜�e�����p'�B����`c���.�/b n��s:�T*U8OɪPf�����~"�c�2,�W(
��=��.�
�ʔb��nEYw}v-�r�ߝk�ݢ���ߙ�q(��!���=@4G$ڑ�MFN� i�0��pl������ҢL̥��ޅ�/��;^��������_v�=�ؾ�><�����+�`����8{պ�����ypg̺ Za�Y,_��ꀻ�o{�
������a5���uh8��>���S~�����N���o?��������M'G��{7�t��i�ևC+��2F�b�o�}?�z�0!���a'��� �CYD���M!��G:���Q��T�V�-�^��6g��j^6��f�lmw	���cѱ�\ðO�)��X4v���Ea��̱m�j�c�$06���`��^2�!��5_��p,�bߌ��\��B!�1�!{���vB!��Տ�i�����c�c9�_�V#!�B���l��R1ҥ` j�S�6��&��X���Ղ�f�E~�t)�WI�_��/��c�oh�w���Ex�����7t�Wy�h�o(����YR������[�i`g��X<�XgW�>m�0�a"�60�a��BV�����_��杗r�+�XGx������_v�3{�L�<=�������>޹�˱m���h_��N�v�?x�Pkv�������_��W#m�:]��� 	��قV�+V^�s�t�ħ�9�������{hb6}�����?~�l#_��|w�P\������8�}ڦ������]Xװ�t����o�BH�a�O[��Fv}V��������\!Įd�TzYPR-����z��]78�kp;v���u��v�)H��-��Ƞ�3��5�p�{߅��c�@�mξ�ލEa�~O%aZ�������X�@�3R��p'�`<�bߴ���	!��F0�I�k�!�B��gp` X�=N�BY+��	as03G��B&�D*�(�s���R칠�X~�!<J��ʰ||� �X���ߚ,n��hͯKt����c	��*�B�w(�&�f�����Jw��7�#뀡ő4#8��p`���9^�B�r��I|�_�§�y	"��������s]oo~{G��������g_�I�6����'�z�Í|���!r�X�-����_��y�����x$�Z�],���V���"�n]���w(�[%�^�jO_��sy��r�4�����dO̦����s��Sɔ�h��)9�X�B���O�緎X����n�Vԑp8<�ARUm[wG�̮h����躑�x�@W�e>�!�
�]�����{_ !���%���>��N]�,¹$��y$�I@W��C��E��b/m�av�M���ã��)<�hw����cѱ�\-�Xx�Sn�E+T�S�9�@�h���O�����^��Җ�Zߍ9(��P~m0d :/�����S���a6�:?�J!��#�a%5����B!���	��E��5���-��B!�Fƺ5l�Q07Сd��)��g�Ng�.�@BAjџ�t�*/Q�3���R,�P:�� ��k��\?�ЎlIV-�a��X�w�0;$�C7�P7��w�M��k�s�C��;�F:�DS�̘84k@7�BH����?��_���Hk�W�{���vr~hmW���s��ɹ�љD�d:�H:�}.��'̜q"m�Љ��#_��ԟ~��C�Hh$�P6�5e �����l���uD�\p+c�ۭ��DZ�Ъi����ՠ���<��To�hZ+8���o��Ck;Wt��?�(�����}�A���} ���tGU�P1�Y��L�3�@ƀ�U�Q�-
��.8��.��k��#��l�{����kα̱�|��;��	�;�A�,�h�J P��9�81?��OCˏG��CQ�����H��X��ϰɁB��/o�r�V�ݺ~$�B!�����B!�rr�C1Gmc7B!k��'�����) �@ra.�CM�P�
�6O�d�W��~�X���h!�'z���A���q;����z����Z�� �wi߰�M���Kw�N&a&߰'|�1*�:eFp<�s�:����͖BZ�����t������Z�����ߺO�����o����oi�̮����}���-�Jq���>��G������
��d�:>y�����@!����Ul�+�ٻ��������T��U��H$�`��PNAJp\d�m^����~c�9���8�X�6'��WCCа{#��}-c/+ж(J	��ǆ# �����'���0�]0�]��E�xa�-�B�n�$3� �B!큥m���c||\�1��B!-��ʾ�?�>�!�̒����L��;;[����
��ʰD��L9V#|D��לh�7�5�9�?4%<*/��y�h���Q~�W��7\�����x0?71�Y*ǚ΅px����\�ޝ�B����)�ٗ�ħ��b�wEAV���<��}ý��n;Ж�ӗ~�O.�_qB*/<V��d��ƣ�&@!��Xa�S�4�F���H-X�LAM��0{rQD*��W�݂�vAJ2Ю
�-dB�ݽ�d���E�ns�&h��~,+X5#�$��6_��yA��jl?�1�N��\�C4�=��2B��z�'�<;i��\{\�B!�����p'�Bi+�0	�Ũ�B!�D)�>�!j$���A:��:��P�av���(��vg����Z�e���ߜ�Xt�7�܂��n/�z�A|C�p��7���B��r,s�%�p�j{�f9!����Ӹ�ڟ�Sx���?��E����n���V[�-nyp&�R���}):ca�����<>�ջp(�'�R�bb[�қ���Zfr�Ш��)�.����X,^`�
���U�vQ�]-Vy�#N�"P5"��*J'lk�Y��'@�0�;S�V5o�1������d�)�\=�w{K{�p��O����3�����x��R���d�7��򶅄Bڗ��\Hɺ����!�Bi��@�G��B!+�h���*�#���X�����0��.5��b1�B,�2,������9�2�N�	����փ���k���m��G��7t�c�ܯ����P'���xvR����	!�ɱ����_`��_��NY>�<��?~߾�9�mp����cxߵ?���~!��!�¯�>�O�x�YB	��U!f�c~z�n@�ѐ��P� �_��)H�lo�8�'P5F�*|��[Zp��ƕ_���Ae�����).��5gؽ�xI���ī� !�ZĪz+_�E�r������}���`L`(?���DGg�xf���Qx�BB!m�l�������B!��=��]�/TU"��i&R:uB!���U��!��@R0Rs����:�!����߿C�����w�=��z<D���eB(uY[Zw�����*��[a��cY~��Z-��Ҿ�`���aw�oXC)Vi���͟?����9!��r��ځC!<9�C*BY�X����+w�^��w�� �g6��_�p��ڑ��[<1��_{;>��sq�� ������;��o}�pH!D��!l�3Ы$���F*��VhUА(QjQh��{�=�)��%VY4C�*�����$���Ħ��űR��l�9kns���a#L<�Z�2�sf����̥y����岗�jia�Z���֜B�0�.���[6���:��ޠ�ԡ���XP:�oN�S�Y��BY�����ވ\Qoo/!�BH{��*:::��� ������ɶ�	!��eeK�{��P
Jf��@F�2�")�ó�OT�%Q�%p���7t�#Z��+|��;ז\��R�X��+�2�:#�U%Y���X���p,(�rY��+t���~���"��^�U�oX*�͏Ǻ���>��.Le#xvJ��&�	!k�0q��?��L�CW��X�EI�������_��T�ʚP�����7��=goƟ����C�`��$����o^!�o6�j8u�D��Bva�D
ꔊ�b(=��"�@��0����#<5��=P��x��/�
�b]fw�P��zU�]�IKU�AEH]�KM���y�LM���e�tQ��ۃ�n�w�9���iz�a��5�\3Zj�K�T�}�|�X�:�o��)���F]��v��}Hk�8��c9d�cBYt�h�ܹ=�� �B!�GoOO��{�wB!�^,q�@�}UKC/x��;</�w�H��;��C�����_�ݹf?.�����[���K�*�����EEY�	;uW�;b�",ۼ�,{�+� �;�P�+�j�w(��b���+�y�s��ǻ��B�{?���U��x�4!d-��Gb�|�m�c��>��a�e~��{�ٜ\i�jeM�M�>�O�������o���B�DSLl�^�J��	d3Yh�V�]+�H�XLf����#N���P\p��u�r�(�s�y�u��5{�])����|�u׹��ŧ�Ƭ�">G�n.-���Ax����ι��{�~I��U	Y�q=A�~P���ǂ�{�897�?��P~���^�H���1ު�BHk�ѥ����!�Bi?���G�H��5A!�y4E����!�g'��d�N��@���9�٥�C�^���z��^/����v���/>��_��/�U�<��}-e��|F�c��8�.�z�a�k���B���/��E>a�k��l�o'G��CR���!<5�C�y��Ҏ���U����T��?�Z�>!�15��gnz �<sk�5p���м������N��_~
�!�Z2R��B����� �����0N���e�ca���mZ��*p)��l���R2A�z�,*�C�Ő�G�� P�C�g-�����B����&?9.�����#�k�9��!�5�6�7����5W��e�|�
�/>�,b-�ŮF�1x�=� !��c���N�Ø�-�/�����
�`�\O�@gk!���/"��`]?1�N!�Ҟt����!IB!d-b�b�:��]f��	d
�Xb���=B�A|��5�[�z�c�B,�",_ѧ0��R,�1��Eٵ�ؽ=��Zʱ����{e��7�n�	]�l~a��z<CO�P�7��m������I��Bx츎���;!�����'�������`�0�\�{��õ�<����)�^sw��n��?4�x��􊳱k� �k�
!��1ءb׈��P
����$0a5��д�a�*��)L9ũ �� A��*{ �z�,49��kp�+��z�}���5�q�׼��������qNuнJԪ8�<_|w��ͪ���U%j���P�[��|������k�42ip�
�/�Ǝ��H�rΥ������ul��XON���D�B�J�%p�F��k�0!�BH����l����	!��Z�ܫ���bC{bz��eR��/��������n�bE^��G���>�Ǹ�3��W{��u�|C[Hݻ��x�9���P�	z�y{�e߯xP9��/N��Aw���
��л�Oq��������+4%���ݠ�0�xu�Wh5�?~���&�����{>�3���O��]v
B* e9<�����C�	�5�d��ľ�������ڀ���K0���γ��q�S�ˆB�*��;���6ųP3Ә���:c�]`�U`w�KRA��T^�v�|Yh�X�Mh���"��x��J��s��c����W�U� 8^���V�9���A�KbW�\Y|*	Q�/�9��*�+��� �h+=�Q�hd4��%\U�6�D�������9��\�50��QL!dy�
ɽ�ttPC!�BiW"�4U�n�]FT��e�ӄB�.*v�J�&�L$�Ni�R,U����=DE�����
������%�rNX�e�+��j�����Bqٕ3�.w\9W9_�&>�6�����
�� Ǖk���⋉}B�\E���:K��J��B�~�w����X˰ܼ���Fb���x��^!!�m�du|��O�����j.۽ĝt���o�|߸�idrk�}`M�-�����g��헝��\�Ѱ�ĉ�$�������_��"�����C!�ܫ#n�bnjX�_D$�"R�%�^�ك�"��C���dE*�P;��$C�KBՒ�T����}�k�^t���׸�c���s�GD+� �����|I4�r�
��E�ҾB���_�D����{U��?�^�`U�pe�D"�s���\٩���u\5�52�\�/΅�رt��1!������w'�B!m���utvbnnN�1�!��5B!k��
�2�����R,)U[,Ŋ�U��l����7��s+����v��l>�T!�(��]�%���z��Kߓ�� �Nm�X����q����U����p���R,Q��'t��Ω�����%zy���d%���Ӱ�B]#�0"}8��c9dX�NY�<1����{�ғ��������%����<| _��1��Ma-���%��w�/��8n�ճ��ғ���@���ff!��|7��ܚ�!dmb������vf��sЭ[jZ��H*��f�%�^�HU!N���Łw��Q�&
�/���Seؽx�x��<�s�sn�n������Տ3�.��jw�,q��z�+ /ދD��^�w���w�<6cQd�	��d��^�Uզ�Us��<��Y���6��Ąى��I�BH#�1M.�g��B!�����$�n}Pr*B!���ҧ��!]�,�'af�&5V)V4Z� 5M�˯K&�^O9V��Q���5T̋����?(�Ek��Z����)�p1VsB�2�X~Y�X�`՜�V�%��
�aw/�P�����	��2t��GCW� �n<vB����	!��{�9���=�Kw�ǻ^����������y����'�ܑiܫ�Idp��?��޽o�d'^w�VtD�֏i|6���z߿�y�2LB��*�U0�. 1}zRG:�n�+lX��$��JcUN�r���<Ghw�{�ճ��778ϩ^�>��w#��n؛j=�9_ٞP��fV�S9�
�{�Tr�����K��xe��o����F����RM�.BVb�"�1\1�5<�t�ON���D�BH�X��^����	!�Bښx<���0��!��V����rK���40�!���B�$�B%��������p{ �j�sNT�%������j����2�~��>�������潎k�y��by����/(S���\
��۳��X�oX�u��)(�N7u���j� �'��͑��4'��"����!���a���M�򒓱m�5�����;�?�o��4��Ybm%�`��?��G�՟=��>�x�v��V֧>n��s��#�3��u��Z�1���~��榧�N�A����T�]��D��F5�WRj��f�|D)���6.��T�0�S����v��Z��=W�f��������߽,��.f�"R�߽�~�l�]J�4��5��]���C�K��QY��t�B��˿ot��[#!�BY��@c'�Bڄ���������G&�.����q�7��^�P����;��}=CQ�]^�	�׶�����m.��r��)��+}��W�5�`�h�~�����=C�B,�&.�*yx��XA��A�n���;�e�0&��_;�;ABV'V��և�㶇���x��;q�����n�YHeq˃���ñ�H5��0��M��_>��|g�4\�_|�z������H��'�rxp�qBH;V��ׅ�)�@f�2�4�I)u񶁚V)Jل(-�H4�.'J	��a�B����E*g(�)L��J㒈�?W�&�w�����YrN��݃��e�dB��q���h�t��D,	���Ʌ�����+��%
��r�����>}#8�w��:2�B�&����b �B!�K<��^\��@!d���Wîa]��&��(H�E/0s	��q��F�ܫ�C�2,A����h��ʗ`y���(ƪ���y���y!�8Y_0����݂���{�Y��d��
C��z��B7�0�_�V��8g�	:j�NЄ�Չ�W�}�+l��37��݊���)^z��4~p����#���@�a�]�B�
�[�`w��ސ�6b���U�)�l���p?� �~�(��BښH����6w���9��BɤVhi�B9%Jl��Tv����Cx�;o��T�t��m��I�W�L�c�9�9��ZƵ�:��F!#f��ڝǵ�+*��{�л��%��HUja���D,�<o�ۛnw[��Z�EA���5=��(.� �7c�����̦i:B�&�ʷnZ%�B!�K$��^�wB!�E1�k$���Y��H&�	IMC$���P����B�OP�K�K���b=�X�>�!��(f_�p{=~bа{#B�~�bP�Pf/xt�op���b�*��:6�������wQ	�K�]�͕��=|Ɔ.��A<3��v'��>�&��/?{_��)��s��׵ʩ;��/��|�?z��ٵ�D������Kᦻ����8.>m=���:k�0b���B�?{�<s�<}i��	!�K,��v���EHN���#�ZlY��
�va����.ѼPk���ցN1�~�ڃꮡv�M��&H��굼�n�ZE�Z�%�n�OȒ�d����㠂�нz�v��W����ұ|нV���X�]E+]tl'f&5�񲘁��$"���0��[�B)�T�B�Њ]B!���!�:?�R_ ���h��3�4l�B�'
��t���bq�",��k�ӳ�]���-����b-��⠻��Y�b��
��6*��H�,H�=h�=�_�<�u,�����B����y�~�X�A���v/o�*�������tF�6��v�Ơ���(9�� ��!d��������G[�{*��1�����v�a��������80�{�)~���	�u2>��w����C*vo�[��{� N�4�xde~�V���}xt�	<��	<wd�p!E!�J<��uj!Ԟ�<c�(�,X�O8�nZp��۽B��!w[��j��&Q�]u����X�Z�*[��B�[��*H��Ya�Z��+���c	 �N�=侜��hι&'\Ʌ��,�ycQ��WF�q���.b�,GkC��z	ZU��v�%�^�怹��ѵ�v蘂�s:!��]��ܕ��	!�Bڟp8��(�	!�� �b⌱0�u���G*�F:]y�g��������9���"��j��ay{�~>��S���m܌@����M�e��A�B�|3��Z��Aw�?(�����r,g��t_Zw����g��j��
�-;q#��7��ƑL�=�C��]%��0ٜ���:R�,6uᬓ��{s1��R�w+���)<���x?�%���b��y����f�����y��F{�}]_a�~�c}�0|#H���Z��sx��la�>�qxr���tET�t��e�'�YB�Z(�HIp���{�۽�)�US��.Fم(�XdW=Z��T��TK�]r��]�w,s\�+.���J�p{�d���������A�P|���f�Es�8�^)f�D,�he~{#�Sв�9T�5�R�{���oC�Gнj\�l�&���g�:.�2��P?8�`|�awBYk�49�"0�D!�BV���Ȇ�bZQoqQ�!��e�j��G&�F**x�V���;��A��@ޡ_)� ��ӳ�����z��Av� {-�ߜ�8�Zй���IhY�����?��fz�A�B��{�r,Q�������s�a--�n�a���ŽU"�m�x�`�R�������BZ�'�����P8�a�X/N�oV^���Zy���Ɣ7Y��'f�8<1��[��<���N#��'��M���\
��쑃�y�w�;���8z:��?<t���G���R���h�,�Kf
�LV�\*�م4fL��Ǧ�1!��%,Q���al�/6�O����HYd*�QU��8e��ك
U"TU��.<�ϭ��	O� ��ze��W��"�>�Z-c�qa�� �=�V��pCZ��E�r�G.��+X���_<�tY3������U�w��X�����97{˻g�]$^��*E���g�]6��K.�Cї���B���P��4��B�Z@�u3�wB!������"�������U��BȊ`��箏`sləcГ:ҙP�g����ޡ�Xk!V�R,a��Q����^[1��g�,�o�����m��V<^T��b�]���kz.�x_�����;�ޘr,�gh���6��ݱVtX���:�n=�������8>�?הӏ	!d%��K���=V1��0�ׁ��z:"�툢+F<Z�PwD��Lgr��F��`>��L"S���&��Mb|&Y�������o}���!�����A~ƘVhZ��Cv!�d�x�@�d��L�P�W��k*TI��]D)�0�� UZ�Zs�������mέm�w^�V���F@��{��%p��=�ͪ)����Jv/���W�w7��&b�ir�γ�W�M����SsЌi\���ً����Bڙ����6OB!���X�}�w��ƀ;!���eǠ�����Ez>�D���b�@�X��w([���.��]K��a��yR>����oݯK����	�{�؋�U��^�Ң���z�9�{�������������
»y����B/O�o�o�+�9�?ق,�]�EEY%�*�����@�9���+���zh���(��so�"�;��x�h6��-�aB� ����㳅���HBiY,Q��~��1$���
���
U�*�2�^��`�\�\�,����
�����(���9�X��{��[���B,r���y	\vAH0/z.�����լ����K��W!`���M�}�F�@[����0;��^ӧ"�?Z�-�d�S�"���BU�4U����B!kK��VP�x�H!��la�@Zb���'��v�?��;t�E�`M�v��t��+Ū�+x�=Hx���{��8)7�5�&��s~�2jG������J����)Ò���A<C�sd�����s��dU������b�*�0X�]f=P9�c��8�����c1(��xx"��r �B��BZ�����I����r�!�(%���{	UKk�bT�%�;ŨF��D)�F	R5ڋ�c��TS��-��p_\��d�[!�����ye)�M�����B���p��"��9�V�W4�L�*	J� ���aq���
�;[ݭ�u[®\o�C���<=N�B�U��G	t"�B!���w�LB!AY׭�Q��)�MO�C�T�%��[���!�B�Qx�+����<���X��s����K'+������^>���c|���as�kz>��'�?��ceʰ�ޠ�M�kI��^k�
���2����X
�W��;A��>�X΂�z��@~��>��?f� N6r8k}7�C�暴c�:!��F;!��'�7�pc��,f'�C�P�)����@�� Uoc�S�*�-1Gu�+�[
���T�[�����%H��~Ⓦ UK���@�St	N"��)z�͋ϭ�V�v�"����y�g{�Z"1Kz�[~�w���~���
Y�Zjog��+���K{�hUo�]Z�ͅ���HO�V=��ū���H�^��Z�$/�4�	!�B�A��4u�il�BZ�Ψ��֫�3�0;=LhHi��x�=J��Qޡ�oh��˱ľa3J�*���{��Z�Uw�����e�+��LY��9N��k������f�Esr�aP�Х$�����c-�_((�ҍ0��4��~�����6�	���&�Y���B�wB!+Ʈ�N�M#3}���(�
)QȽѡ�ʦ�@{EÂH�rIբT��
V�-j�)D��Pu��+�6��$�rZE��KdQʿ6��$��� K�xQ0�3��<�	�;���,���}��Jf,�� ތ��E�kȽ ^�x��~�m��wWUs�������!3{q��rԮ!dU!۸�ɓB!��N7�C�z�B���O�I!9yƔ��J��Y�;���EX���7���C�2ޡA�E�Y2k��A��~��<���9)���C�-ê�c���0뼴�`�e�J�dʰDs�����ߧϾ��XA���EX�aw�b,{�=h���gX����Uw���FD��+zT��G�b��濏���BY)p'�����T�t=Н=���Y�&�����ea�qJV�Z�J"�(��#R	D���vQ3�E�P{�w�qq��x�%@9%/�IF|�<%���3���&�M�*=����K�x�s+E��H#�;C�N��X(f	ּ�+���w���л�^!8�����"�3�^KSC�s�x^bv
�	�a8�{O���d�BZM2��0�N!��&zݧ1�N!�Fƺ5�7�#�p�DɩP�ۋD"�eXn>b�@����+PS{�R�꠻ES����.ǁ
��u?�P6�n���3��F��~�[_�=XQ���Y����Uޠ���A�t��g��Xr��`A� a��V���-��K��Ɖ����pź.�Cxp\���BHp'��t4����������Q(S*ҋ�v��v{Ƚ$>9(/A�O���D*qۂ]���WTn���U�
ԮP<p�&��Ϛ����4",=L�Y�Z	x��s����b���ʊ^�w����,vy�.������Dw7˹oD��y,v�U���W5��45�v݅c����<�����ԇ�� ~u��B�f7!��*��9��!�BY��0K�$�Bd����ׇ�>\��I9��?�
�{b�|���K���:�����9����W��Ƌǵ�k�m/U:
pn�*dh�W����~�l��z����}+�r����cA�}��cy���=�V�*��t�~�g���+�
��B�@�m��p�)vcB��wB!McK��s����Cv!�D�jZ���+�)�`{��5,D�%1�[���d���E3�����`,j�M"��Kp�
��E!E�Z�����J��Ur�v��T�O��	Ż�S���b��Jl�
���i��6J�jdؽR�2<����%�Z�rXU��R[C#�e��zy!�L@���e�
:6��Ssx�X�BZ���h?���	!�BH����i'�"ÎA/��!7s��,��?\�`���U���;~��/��}��ڽB����縟+��y����}�{z�~�wн��ޡLA��?�r��.7*�^�7�˫�=�.��Z���tw��3��xU��h�������	!��À;!������1y�z���>{�(ғE�)j�-8)Q��!Hɶ���U� ��(U�*Ũ�}��$
���-�p/��s��*��� ���,��x�9���V����7��ڊ��U)B��Ĭ�k�V!�6����pwWT^!�+W
X>�U��/��K�r�V��P(T�&�bC~��B��]������
��2 S�i0�N!��&z�g0�N!ąΨ�K6(�L�ca~��P�۳�څ�v�b�Z�����^�%�!z��[�K2��^j/?s��������~^XU����eY2���<:��,�f`�PQ|��`>aб�_������VwY��t��V~�3��;����#ؤ�p��>L���&�Y�΄B*a��BHC��p�:��1�����h4Z�dC�v�I&�.��C�Ά��H����dw��6��Ū�|\�/ι�P�S�Av?A�/�.+5>�n��~��H���D���J?/w�M,���.�|��c}�����`,�7�s�$�.+X��J⑟��r/W�-�.hk(�[ZdCg��!^Y����.�V��c31<=��B�JbH�]�|E!�B�pיG!��`�@gd��>}*��B4��{�ڝ��A<Ċ5E�������;<;<�z��V���;����<(7_�-��`������]��ׇd'`�<O� ��tԋ=��\鑐��ʌ�����C�>~aɇ�)Ʋ���	�;ׄ�"�Pv/̇�J&�����u�	!�T��;!���Q����&���T����m�@�W�H������r�}�i�l��}��XtA�p{�gԘ�{a_<�
�{�M�(�,'<y�N�b�L������g�������[X�o��d�Y�\�������)rn�V����A�u����/`���e��)`�ޥ�*A����](^-�4l�sص����~�~)jW����������wB!�����o�@�>��BH{	naT����r[{4�*�
z�g��vg���7��ٽ��ܘb,�F�K���t�]�#V���U̕G.�kb�I&�����Z�e<?ْ,�c-ޡ[����U���w�7X���.w��pWUk_�_�����rн��|����
��tq-D��B��	!��/���Lt��#�0�D*�H$�f�im�	�ˉS���8�liث������W��!��av7�?�4�^k�}����$h��� 'A~���k�BU�yq�J�r
W�9W�'�^��p��w668E,���]��hxw�ݗ����{�!w{��+�^��Vwun����_���G�&��N!�v�� �	!�B�F@�L7V��F!��l���,����L�-��J�d�����|C�B,�b,wqJ�dC�>~bc}�ʵ�^��kʲ���V�������0|��skg��;tΕ~�}B,O9V#
���� �a��ݯ˴a��	Z�'|h�_��0B=���x�~!!��Qp'�"ͩ�!��I`~��)Gۂ�0�Ӹ\�r�P��
B�b��0U�(T���B�W��O���{�O�
�7ShZK"V#~��� B� ��P������A���fq�K�r�J{��{i_o�]�� ��\���{i�5��U���л]�
��-���8:^�m�3}��p&�kh�:!�T�K���ks!�B����}��N!kMQp�z�p���G��,���X��/t�e<C��h���m�b�P.�^z���b�b�+����y���%Z,��׎c�ʲd6b0x ^�#,�U��nw����"�z�����z����*��z=C�b,��
�!w���.�"�0=y��^�m��~ܵ?��W!d���;!�O,a��M�kS���@bJC8^�B���v7�JV��;C��R��`Ws�P��],JY42��/��E�T�|�������yy��]�r�H��Ĥ��~%:y����	�~�Z��	Z�߃k�C��}Ѐ�ۚ��%���W��+��.�� -�^��-�[rv
��q\����QܾHf�\BH3�%/	ҙ!�BH��	x�g��:!��֠'���M
"s��^H#��J���J�Dޠl��������ڽ}Cg���ؖ(�jH����{�^�E�<�V�W�Z�[�%�Z~�_�c��;\���	������?εJP�����R�%*�r��aw�B,/�01;�}���߄�ᎃ*�S�	!��a��B��NK�ڠ�3u��$��@�x����R2��^b�(��lmwګ��m�BTu���M���Jc�x<؎j��[p�MA�4Bj�����f|����e����z���{#Rq��x1�n�<��X<�tN-���w���p�lg0�D�JQʴ	V�	W^awQ��K�*�4d-S=�"^ѫ ڿ�>��Y6BH#��;�M��B!m���n��=i�wBiw��p�`ɉ���	]��˔b����fw��v�v��>{o�V���!����j;.IΉ�ۋFy]+�����ѥY+Q�����]|��kP9�^�U�K�K�z��=Cw����S�U�ݟ����^lu�'������t{OdA!�=a��BH�{5�;�Cf� �)YK���7&�nkd(�P�x�J��	����)�@�ŉ�����
Q�"���P�h�h�g5H�NПaPA��f��i��l�T���:�,�Ɔ�~��Z�+籼xe���X�r���~��2�Uy��\���a�D�q�a<���o�0�N!� �˽�gp'�Bi{��`!���@g�"!��-g�aG|s�Ǒ����9�w�G���J��C�2���$ˢV?ѾV�Ń&{�K�ιz����w���֊�؈_g�!�Fd�[�U�O�<��8X9V����q�й.�	�<Cw�P�˫���@{����#ؑߟ�m��~�u �����[Bi'p'�R� Lu�c��Q�'�BS8$L�����.X{�&:��^"�P����nXO��|^qЀ`{�k���r��k>V[��Z�,���(QJ��j�=�%������/�Q,jW��]��ڣZ�
"\��5�	W^��"�J,bم+�`��p
���Sˍc��^L����}:�4�	!�fd7�����!�Bi?��t��u^BH�)�x����1$��Ȅ�D�
�/�`)~�a0�P��"��X�+Z��Z�ܝ�J)V+z}����K��khdAV�ʱd�K&��5WU�UK�=�W(�s[��	��CgA�o9�O1V-���f�������	\����QܾH�0$����wBYÄU��-��Ǳ07W�*n#(�B�����[\�م��]��R�	��V�y�~���fo���V�Z�ZF���<��8%�J����!��_���aq�+f��n���ܗD��vww��?��'^�-2�v_�$X9���|&�@$�<^?A�s=n?,���!�%����=#�!�BH{��]�Ò�BZ��.��0fB�֑����54���>>�"nk�mm��-��S+^�UK�}%K�����F�Y�s=��Fd5�����y��� ���2��2Aw���Wh˄�E>ae�U���Fc���z���G�/�=*��q��0��1�N!��	!d�Q���
"s���J#�����b��@Z\�%��u;A�G������	��	V���@��
�W�_��_���;̾��+!,�F1KD�d��d����{��{Q�Z
��ķ;�ޥE����	�{�ޅ���@�@��VÂ{.�i����>\�	�6o�]G#8:��B�� ��T:̀;!�BH�J���wBY��:��y�OEn�n�~�X2�v��v7�P����u�g�Zi\�+�1�.p�d�K�X��:�٭DA�j,�*=u=��Z��^kK^a����+�����X��a1���8��B&.޾O����BBY�0�N!k����7���x��b�bh�'��lnw�j��o#轷Q��9�^�p��
���'o!j9���
E��(`-_c���ts{���_�h����m
{{��K�j|�=�he�t��e@�+E,?�JZ�r��C�!w�}�4��8��4];�၉�0�!�o���L&���!�BiO��{A`��BV/g�aG|s�Ǒ���D����vY�P����n��o��b,���Zq�R�:���h��Z)Q���Y��ˍ���3�n���+%j��Q�dz���qgq��m�_�5]⿪��E_�=���.}Ӟ�N���b7q;v��E��$J	�  ���3�w�ޙ;��|���w@B0x�����x�}��p�
����u���w�=�KU�e����Aw�kKs�`��3WO���靻� `�@�  � ���S۴�x�����^�B�B�h P�	�+ũB�+0�����ٝ�!bQ���i�Vq�&q�a}|�Z�EL~N�Ǐ��%N�	��BV�<c�Ƕ�͏)����ʦ��Y�]&`���>�J�lo/��uZ�����*��]"^9���=�Ӥg����G����  @E���kx     ���Ɔ��Zw  &
�}�B��P��W���]l�;>a�P7�^�x�A����]��^�{�}G�#����;J�Ϊ�w^ܹi�sTH�$�FA��r��y6˱��^�{��.�����W����0�f1�q�����ame��4����ct��_ߪ��g|� ����;  �0=P�'��h}�.mV��QQ��"�B�
����xT��@�	�A��e(H�P~1�}<H|�܍;6���sl�Թ���-jP^���63�|�:���Z7��=_o�(b��v����c�'`��������V1�t��:�TA�����umu��7�ӣ�;�կft  ?�u����     #M�Z5or-	  `p�
9z�b��n�Qm�J[�"�۷��;�l/��}C��!�S���
ǈd��y�}Pb�9q�%u��?�-l�e�>�
���U�.�

���B��eeX]ϰ3Y�������+@�n��mA��n�KtB��w�Y���:j,�_�;D˥����&�w  @FA�  F�''��pw)An\(��%�L�
�z��^�]ּ o[��l�-��t)1���ڶ�U�*��$�eߛM�I����{�#L�OK�
%��;��K�_	�{�js��U���A���UAw1�n;��R� �J��pU]���%��ţ4G'�׷Z�2��  i­�;�w�<��.��    `��6��7
   �,����D��Y�Zڢ�bg�g�;�B�wh^�lW��lhO��ݽ�=�Οݿ����@�(b��a�?��ų�U��c�r,��s�����>�J�B�����V�(�6���|C�,x�ۛ������S�i����M�$�  s �  #�g&�4��V+�=K	��)�(ſ�jW�=bT�(�p�	Rq�)�jW6�+�)�Ͼ��c��)ہvS�b��I�L� b%�=�	����ΕD+C��x"V?�8�}��]lfh��;�����y��{��agG������}�R���R�f[�����p%��=o��N����si�t�~9��� {��;��9:X
�!�    0�l��Tom&T�L  Y��x��?�CͥjVv}���p7-���ll�)Ʋ���Gt���V��B�l<�HR�Y�?�0de���8�+t��
��,�.���q3�p�������+��,�b,��
dpw�� -�c�_�h�>�T��GDG��+w��$   � w  ����}�<b�N��$Ԯ���BC�+P��RњLE*&H����P{2:���40�{�$�ϙMQJ�|Q�)ռ�Ĭ8�w�u���kOؽ���лJ������PO�r�)7���k	WRъ�gv�!wӀ�+\5D�J"Z:�������h���;  �;��q����:    F���u��6�u$  �����/�ݡ��m/�8!�����o�K��b��G��IR؍|D������!�R��b���h�g���rAV�>a�83������{��.�<Ü���<C��s����,KA��b,~�i�y�Z��b�r,a%�F�&}i��Ν���.��&� `� �  C�l[�ե�l�6.��S|?A��
S}��8N7�.����1�n��bwǑ�C���~���Yl`Ⱥp5��J���lSa��YI��b�L��!��,E[C_�]|����֠�����6=�U���������įEA�E��?�.�����\E�  ��|����~m_[[��G�     -VWW���9��gh  ��`��5Y[-Ri��܃B�E���b��,��<Ġ�{X�]�Cdb�����
��B)
��0�m�{QH�{TAVZ>�jlt����~W��� ��	�߀v�=�3�����,����
�?�.�e�Xn��q1�`C�w(	�oVnї�s4vAw  4� �l��}�~qJ�u�'L��Rg\�$F����ıLX�J�R����C�s/@��7,"О��$��a��&�sE8KR�
�o*h���6�/�Un3�j���A%\Q��՝k(^�	W�vwؽ���=�*�mj���f@�]�����;┧�]����n���g�Sm����5�[ ��und��]]E�    `Y3����  `�����e��v��r`���]/�./���,�����2�I>ԎR,s�8GÔ���8A��d�
���M�B=+AG��ߣ{_�������7�r�������лS�%�|�����/��[zk�6=w�h��Yzu�D�U�  �6� ����ǖh�l[<�T�r�z���=H����D�(B�
Q}�f�=\�JW�t�=�8�:O�3.6�l�Ra�~�)h�mZ�2N��%��vw����$\��X�����n�Q���Ղ�/��C�`o�B�,X5i��w�Vw퀻0�#`����;ݨ�)�q��sAw ��byK?��b|     Á�u��V�   ������M�Z���b��>�����C���a�3Tb�<Ĩ�Xq������XL�3Ho�X{��*kY�V����y�6���vUa�n�>��*t�_P���wz��a1V�k�����B�����fe���G4v���e�����
  �� ���](����2m��e�TX[�l)�>q�n�SrA*<�֬����Ѹ�F�=�@{RB� ��������MB��=o��-A+����qQ�v����b�]G�����L�R���;����~�muϻ���"^�P�����b�]lg(�o���wό�Jy�~y�ul���  �K���U�    F�L���n4giw  H1ؾ�ۋ]_PY��hm��kb��bp�ݼ�]+��ON�}Reyuy����3��Q)��K�X��1��V���0긨^a��Ӽ/�+V�]�o��v}��r,y!V�#l�o*=�N�{��|��fw�Pluw���G�Aw  H�  �|�t�ۿD�K�,��UAv�8%�Kĩ>a*X�R�R�!w�O����v�P�y˂���AV�c�̉3/�s��`C|R��(v�4[L�'x������&��A|,_�]%bQ�x%�u+w[z�U�x��:"UG�r�+���ٗntW��VY�]�׷��\���=@�3���z��L��%  �Z#O[��¯8���    ��`�u�ǟ�M0Y  @<���:m-�h�U�v��vo�]]�^���y�q�CYѕ�Ku_r����c=ԎR,���:���H� K��Q<Bռ$|B��$�����m�m���{��>a�z!Q�_���/K�da�v�V�����\��Y:��x��+A���MY�}�hl�<��N��6�4  $�  �A<^�����Ze�j�Bp�]jkj�������(F���U�������(��R&����Qm`�!%)2���e��B���
S:�+N�d�=��%����M���c�"U.@���u�^SC�/��ks���
��l��v[޻��Fw�pp�w����{k��ڢ��}��Q�n��7��	  F������ǯ���~��     �����x��,���  Is����]ܡ�e��X	����(��x�����աv��vm�Ђ����cj�Z�=�0�^-�&��fEYq�I�c��m�QO%��>~�_(����2�0(�.�Uc��ݒ��*��G��W��5��A���[���9;w�^�U��-� �6� @�8{�H_<�IՅi�-�\.�E)� l
����L�*x�{�)aJ&>	U���P��A��m�M���%Zŝ������_��T�9l�S&��ld�#`������9��+�64�
V���������/`��{��v;�O�r�"t�uĪ�L�R��1��:�/ыW�k��9� ���V�N��[�Tp    !���Ưn�Z��	  @B�
9z�R���ߡz�������a���j�P��n\�m��Hw~Rb���}�=Zw�bٛcs~���"q�(�4
�P�|\���0�.)����ð2,=��-Ē����^QV��]��+�W�n��M��d>�t����4�ߢ�.����m5��k  $�  �����g���봱��ry�`��h]�k\(�ۃB�wF*N�UM�J�e!�����(��I�Yx����!aJ���V\1+�U��(a��e$^���)(����V�:��kto�m���U[��os���*���sE�B��'�VW�\�B�]y���~��8�x  Y��p �*    �Q�?�/6���?   �S���K:�5K[K��[,��ؘ�7T4�������C�2,U1�Vȝ���w�h�a�P{Z�XIy��X��%�/��%�����b� +��Xi��g�J ����J�r�}�]�:�_(�{�BwL_��t��7�CW~�d5+3��cT������z7���  �@�  ȁ��p�uy�,'�K�RIj�5-D	�w��6�{*'
N*�*L����a N�>���G9Ԟ��{�96�y�Q#�sd*��=FR�j���{����zawy�O�2��U�}=�*���e{"�(\y���f�^����.���{a_���ͽ�	�_nT��W���4��$  V���"@���     `��V����e4g~w  �I.�K�_*��wis�F�B;��������?���ڃ��@��j�&�X^?д����s���B�&�kc����>�����hz�
��Z��;6ʸ$ʳ��{�a�4jtw�������c�}�p/��4�;�@����ms�	���X���� ��hP~�}��Z(��Wo�[�/�s  �
�  0 Ɗ9�ƥ֝�[����,N��A��_��)�@���֮/L��R�v����~��a��վ0���,d��.�%J�϶8��c[��9_�U��{?A�U�{1����9Ab�L���z�J�����BC���=ls��\K��.�ݫ���'�9���y�ŝ-m`�v �𱺝��f��¯X�_[[�Ç     n*������  `�g��Ra��˫Tw��E*��mm�{��~���ҳ��$�Τ�"ԞU�tl�96�&y����sg� k��c%���vW��x��{.�K�/������r,�ս�6�^������
�
��}y{k�ƫS������Iz�N�   ���;  ��ۺpls��7��r����S��v�h�i^��Q���aJK�j?���)��� C�iVI��3�����9lD}��nf�)N��7�l�IG��.��D��}� �/L��*��\��73��+��R�).C��-G��M���T��b�,��aϭ�Y��x�9:w�~:���^�  �D�i�p��5z�RA�    `Xl]י�����6�  ��O��EZ[Z��R�il���~�|�R�V��.�2.��'C�*�D";�!�#̚?8��Xix{�_�[�e� k�ʱ�'F)�
:v�y��>���zz����W�v��c�W�V����X|�������F�g�Q����2�x���v�>Z@�  L@�  R��%zd��//S��XN0D�
���z�#H	+X)���X��.FyC�Ο��*���!M���ci�c2�tl��q�%}�ax\�
P~L~V��β8%?�U�񠰻)�����U�h�
��,�x%of�	W�x�w����6����h��F�{|�U�šѠFe���D������O7� �n���߿��^�B     `x����w�f�ɮ|  �g�P��tz��Ӵ�,Ҿ}�����=�=D_V��,Ԯ
�{���X���ۃ
�\F�?�9&�q�ؘ���F�(Ϗ���Y.���	Uc�P�/쾫�/'�/��>��:~��/��ʱ�ޡw�f�+�Ӥ�|��S���ͦ�g(��*ϰ�p��k��t��@O\=C�U��&  w  H�����ܩ�-�t�)�u!��u�]���_JP�q����	k^�Ѷ��(��*�qQ�G�cs~���
6~���f�T�y����2�nS�ҝ$^��'����zc���,YK�(Z�3���m���� kgؕ�V��{-�Aw�ͽ����ѽ�t�Y�pj��}W/0
  ���&KF[Zc���h�^�r�D     `8�k�zݬM��&��  
�9�����X�A�9*����b1V�՞������d�C�՞�Y��8�;�d���(��γ}�,?^�*��}.���:�H�˶���Wv�^1�*�����%�9��k���b��ap9֮�G����KZݻ�Y|,�
��0�3l4
T]��O���&/����Suk�_k   Ip ��8�?O_;פ���T[�S�����He#���� ۽-���q!Rk;?	*q�dm���ڇ[��;7���$��ɖ����n�=������DmZ��%�J<O�����D+OP='oi��X�&Y�=�c*�����V��v7���,Ch������xI#C��~���N�����S�z�͠� �a�Z�m;�z}˯�tvb�     �p2w����M،  `B!���^����mj,֩P(z}C��XZ�={V}�y�F�=�=D�kk�Z�=p��X(����,Ȋ~O�'���x��7��vw}@�����G�e�a�׽r,�{�O�b7����cyW�nݛ��Q�F��w�*��/n-ޢ�-�Ɓs��7Z�4  H��  �)�^���}k�[�M*�K�0�J�r/f�E*Y�BP�]���\��%N�!	���T�T�%o�5Q*�@{RBԠ����I�J�{������63�|�16L|��%�*�ٿyK�R9�h����d�Tp�]�����+7��ig�6�Wn��7�p��
�����"=�_�g:G?�]��� �c���~o�H���V��?7��;    �3??o4����y4� �6Ϝ+���}�X^��b��ڮ�[�ի={}�0�0Jk;��u
���C���5�P��1I��;'μ��3l���vq���h� +j�=���F��?n�Y����@����u7��0ms��cy}����+@{��n��^����<C�ݽr��t��w� �͟��nah  ���;  X�+��@c�6�6i�X���1�p��P�6*�S=�J-D�B���s�hI��+L���ݯ��D�#P��-@��v�M�'�R�1}�L�$�)��q�)��6�'�1��T���m
Xz�7���N�{N�����	Y&��NWp��"�.S���x�5}��v�����fw^�p�2K�,R��9z��5v  2�ݪA�}~���     ����5�V�Fs�m�W�  ̃'J���eZ[���b����IWyWz�	���P]�%��ʱ��ʱ�	�nw���Ϣ��q�c�g����:� ��sE��ldE��,�������{L����E���\S{�G�zC�U�U+@˂�U�U�a7̮���momё�5z�����1�xAw  pA�  ,p�x��9�LkKTwĩ1O��/P�.��܋eU�=�u���E�\�8r����$�N:�T���a�C� ���FU�r�0�%J��+J�=lޠ�]�
:&{-�'�hi�U758"��L��W��|~�	���W�6����(\�{o�#ri53���Vw7��y?�{n�}�L���7�!Z ���Z�s��X~���S�N     .�ݻg<�N#  q�@��zf�����R��U�a�K����D�����;4^�|~��3�P�p�z�=k��$��(�
f���(�|��P��'4�T���x^�l���}r�WH��2�0(�������\_н}�ݛ�~a�b,�g��1�����ڬ�����eZ��7�  �  ��`9Ozq��뭋ͼ#N�[ڃ���KJ��`%��u�)�@ej�-L��-D��(X�=��L�ƙccn��</6E)���le�1>�F�$�4�+W�j�X���1ꦆ�h�+okjenhP�ܽA�f�ɽ�iro:��w:"Tgi��p����/��U���w�շ��H��x��V9L�Wt ��z�V[�ᒞ�>;;��;    �2{����*,F  �Q�}�j���7����b%��m�OX����J�0�?���j��U~a��H4�����c�u|�9I�c��K��_��|���b9V�^���_��7Z���x���@�{���;{�;J�p�skR���y��W(~�hhc�.}i�5�����ֹv��e  �P�   ��.�p�H����ؠR�$�dK�D)پn�F�=L���S��vY���s�?�����/F%���*��(��γ}�ax̸�lp�����T��gY�
;�䱰��������
L��$�T*�*H�
oh�od���K��+'��iuw���~�{l�r����'���Uk�����H�.T������m5��5	 0Zpp���m��sss���     ����2U�U�9+�y�6�  ��g��Rn�6*Uʳ78���.�Uav{�a��h����p;���kkO�#���2О��wn�eL��,de�'�g���$�%ƙ#�����$~!u����bI�B��u<��{�Q��9i�]������r�G����ϰ��
�-�L�_�?H����u ��G  0�ON����Z[Z��R�ʝ�1�n�����"U�`�q�]7�N*a*,��&�԰�ړ����:���A�7���y������
Z&b�^����Α헷4���Wъ�_�bqjW��.ޏto73t*W��������~���ze��}j?-�'�i�� ǝZ�����������s     ���;w���`/ ��ġ}����O�v�䴶���y�bs���n!خ�!��/���ů�$�Ο��{��a���y<���a2�tl��Q�$q�,>VZ�(��}^�(Ȋb�;6ʸ$ʳlx�6<�x~����G���x�<������{��A��_�#c9^a�7T�bɼC�R,޷��A��8+@�j�0ͮ�3 �-�@ �&G���O/ԩ6�j�BwIA����*W���{�T�68ОD�=�0�� ��=��{�sm�1g:6����:ϰ>>cC��c�s�<~a*h��*��%-P�O��A�_�\�X�\{�+RyD+�pUp���V��<���7;�UG�������p���t�W�m{{��kS������1�Z�h H��Z�����rA�avvw    �!�?�޽w�x���   *r��+9�/MSm)Gc�����m���a_����c
+>Sp�]ԇ���x���H���1�m�1g:6�s�<�����K�=V�aМ8�⠼°�s��e����D��w�#����������0�нt�z���_X��&�f'����,�������A������S�
=3y�~<M�� �G@�  B(�.l�z9O�o�f�A�r9r�=�y���B�^a�_��lW.%nwft�o����6��2Ԟ�`���8s�8G���~��Ay�Ǐ#L��7�d��MbL����9���{����{W`���|�U<�Jv��3������ �J����/����zhg��|�<�d�Hխ�y] d��+)ݬ���z-�J�677i߾}     ��������&��9Z��  �u��X���YڪlR^����~�Prw�A����w�P��o��u���[�O���ˠ�ä���9&�qQ�ǝ��y���Q�Y���s�U�e+�n3Ȯgc���4���M�}�<>�W�������:�.z��q�*Ў7�ms��݃ݍ��+@�+L�k��r �>� @ O�)҃������z�,yZ�*�J#���������.'(��ۥ���B�,�ޙB$]>О05*�TZ���8ӱQ�ۚ�乒$�H�$&ϟ���gN[�2�E�*�M!Jg�nK�?Ԟ�6���{~���ū�>�=�h��ۼ���{W�j�V����:A��"�ݬܡ����9ze�  =��S7�ί�333���     �67[�m�\_/S�/� �hs�X��=�Jk������<ĠP{��(6���u
��Z+>���!���&�����6�$=6����:gV���F�/�S��Q<B�<�X��M�OL��*�1>��/l����X�~��R�+��*�Ck���?t��V���ݝ�i�ѽ�]���t}{��4�ыWO�k����r�  `TA�  $���/6�6?M[�"���)�t��%���b��`$L��������(�+L���IZ�ګ�U㢎�:'�s�����}�	��|�q�)�s����G��&P��M��A�_|?�2�v$Z�[�h���V�foN^&Z9�M�/���	Vݠ����	�V��<v|s�^�z�^���+� �g�V�Z#G�E�뗙[�hrr�y�     ٤V�9��¿�  {�}E��w�h{�:�V�4&x���P�7+�r��!eXւ��v"��:����_��='α4��1g:6����>�0}q|�0t��!n >J�=�Oh2v^a��$�%�z���^<~�?�������{�g��	ۛ�
�'���7�;+C�aX1V�
���{me�>�_��&/�On���k"  �w  ��K
�ؾC��m*����Z��
T�օ��v����ۉT�Tz��dǙ��2���4�7��>G��X\a*���)��I�v�!^����Gb=�Q�xt�V2�J*Z���f'�����۝��f&gS��{D�B����@��
 �0�
3S-ѣG�Zܷ���޽{t��Y     �dzz�X3Z����~� ��xz�H���hs���K��b,�r,���5�����������̘6��I�?L�#L#�>H1���sl�Թ����5,��=�;�G���T�=-�P6��x������sN�VNr'
�y�����'���]������7��cicI�AO�S�ը��wN�۹��Ɲ: �(��;  t�x�@�?�BkKj��K
bT��������v_�n{�J��la*k�����(c���:'�sd�&�%��|��t�a*j��lއ]�����3�d��Oнs�v×"����OW�R��{E�fG�b�jG*\�awU�]��lk��T���_�=@���{hs $��5���3��M�    2
�}��i�� �'�����p��Ţ�;+��.��>�t�g�p�l������(�'��������o����9&�qq�ę�����ϝ�vn�a�96���qQ=G�s�=����_�<��'�3�.z�;;�^��
;�v{;{��^�W���W�չ��ɶ��D}{�h\��ON��f��bm�  `@� ��)剾~�uA�4M��\�8�h`��˖�S*aJr��d���p��?�`� �����G�ccn��6�>Q��q���sD�l��mއY��3�/39�i���rbC�VKC�P����[��{��7;�j�+Q�jݻf�D���ؤ��=49A/��G˛�  ���,��v����^c���iee��9B      [ܙ�u>�����Vp �r�]z�r�VoSm�A�������՞��MJ��}����s�����1I��Y��8nsL�cm̳5?+�����":ϕ�c����E���f�+;�T��̶_���������n�]r�ݕ��M�B�
�j��=G�K(��f�D+�
*�r�k�s�܁<m��@?��t<T  fp �i��(҃�9ڨT)/��K6�|�T�����ڷ���r�{=��*�qQ�ǝ��y��qu�+B����&�t�4ĩ��Q��Q�����_O��of����0�����w�7�s�}g'/���uG��,A(��ogP	V�h���%Z�8G?��$  �͵�2}�Ħ���7n�g�z�     @v�Ͻ�����fkE�6�  �ΕcE�ܑeZ]�Юo�gU1�y�=x�gY1VP�=�`��g��fq�cIε=�d���8sl�M�\�H���ԏ��͏�-����&x79����U�}��tw���D�Aw�Wt����ao�gO9�b�g�b,Y9V��=.ޠ��x��^;NS�X 0� � ؓ�_�?=�M����-[R0��ݸyA��^��t�T�T�@E�P�T��g����S!V16��4��Y��?�q�c�̱9?��f��?_����cfE����+d�-P�O+��?f{��w�� չ�tW	U����������u�n�{�#`���M-�JK�r� l�-/]��_>N�[9F7� Z �1�V���o�^w��߻w�֫U:x�     �lp��]����L�_v �Qf_���/�+ש��o{�
�P��=ĶW������v�R,�@{r�v�R,��A����8�;&�qQ�ǝg�Y|����ʰ���+�G6�v�]w��8����q��(s��e�)d5hw���{P9V�_���՟���>����h����ʱ6�W顝%���Ezi:G۰ C� �=�W.���-ڬ4�\.K�%!�.��6/t�TS���V�ݽO��~A*���x�L�Fw^��C߇-�I���`�}�8e2vU�q��������L���`Et������ɖl6s]!Klgh��bU�+^��Un�])Z��,Z���c�%z���������k' `��n���TKt�P]k<�f^�~�>��     _�]��2����ѝ� ����E:Ӝ���&�d������r��J����3�{��X:�a�`�^s�K�|�4�øs��dL�c���=?�sQ�(�d�c�3�G��g�+��m{��1I{�6��/�?�[���۞a/��{����O�d5]����궹oVnѷO��͝3��]�� �� �=������-L�N�D山^�=D�
�K����v�0�,0�.�ڥ"?v��Y��$X�8ns�ɸ��α9P�N
��s������{n��T�<�Av�qY������NQ�'t��	U�6��������.���Tb��ʠ�İ;�o,N�__<Bo�=�% V��N݀;3;;K�>H���     ������ϛZ+�Eӕ   ����vn��秩Q*yW|ho�/��-���p{X�]�?�`{V��$C�i��Mƙ��2>�3,�DT�O���h�A�����)��
�Ρ{~�c��#��B�O(�$����w�_�:��7����W}�ns�׷��Tc��v��ϭ2�m�  � �_�\�#�[T]l��ؾ�P�I��^����=�}Ad�m]�X�=������x:�m�1g:6�x[s�<�^����%L��f�=� �\�U��$�(�9&��j�AwjU�	�{����wX��_��	U͐Fw_�]�a�X�'Z	b�����6�����z|�"��u�:4+ @�6
��]�#��x~�q�=���     �����sZ�|铕 ���%:�}�6��`{�/,x�a��'���
�=�|���	���^)��H�P{�`�0�����8�l�9�d���8sl�O������%$��:�~7�����
Î�y,K>�lp�]~Wݩ?���ʱ�<�|~����|�X�����.msWc�x�^8Z���E��-�"  � F����:�-�'�A����Z�����8%�%N!���l�9&�6�ٚ���4Q�([�Tй��G��ƚ�O:c!`%9�fx]��Aw���n#�6~��d�UO�R�34���P�#V����B�����'V��Uo��Wf�g҇[���y�� ���r��pJ/���ܺEW�\A�;    � �w����ϛY/R��'  ���ӟ�ߦ�b�gE1V����՞mc)�C�`�M/p��C�c�u���I��I|?q�>L�o��'jx=h~o�f�]5����iK�/T��k-辻���c�x��'�����������kc����׍z��}B/>x�^���4c �� ���im��Pme�/�^*�7/����@�Rk;��T���ܳl�05�U�uǘ�3g���i�o�򜘊da��D�]5/n�]66�U�qSQ)�����s���"�x,�����KE�]uC�i;�Y�{�O�R53���f���%ݷ77�rs���H�u#O�&^; �\_-�Ƿ�@Q����?���z�     @�8�c�|i��e �Q��ã�ڨ4W|.u���u������b,R��͂�=?�I����f�#̊?��7���hc���o����u����u��Q�ŨAv��$�D[~`ǲ���[�S�C�{�A�X�_h��V|�hs-ƒ��|��4O�*��������  �w ��q�`��rj�����r��Pa�f�v_�}��$���߹7�`�����*X%1.����l�#��e�8B��-Q*�|I�m�u�R����%D��?��;u�
AwͰ�_�R����z��f�fG�
hs���V*�J<.63x� ���Y�Eߝ8H�O�{sX� `F�Ռ>^��<��=��{tee��9B      ]xE���u�y�6���Y   vN�����h�2G�A+>_�����&����!��T��s��ilf�p=�Ax��c���57�s�:�ϕ�5�6?)��d� �°�I�_��o:6�ߚ�C�y
��!���{��Ϣ���V�����g��9^_P��S���=��B�ց�)z�����w�i��6w @�@� 02�r����"\���ݶ8l/4/�	��Ĩ��8�T�°���FU�Jb���8sl�M�Y'��%�Xq����&��l|\!k�*�����kt���t����`�mso
�U���/���Ukk�բ�W��2�����~��	=4y�^���6�  |�R�ǏmQ9�=��G�>�y     ����]�i�Kho ?Nk{�Ֆ��+>b��>����J���Ty�}�����^Ϣh�I��:>�$Α��Q�@��F�1�����A�z�q�@���i��ǒ�U���u���x=D�^g2�H��{�����{�&m���a.��Z��X�����U�����@�,�ʩ��4C @v@� 0L*ЗO���R�i^(�K�p�/�Դ ]RP&P��c���@�+N�.Ȃ�D�Ez2��,	S�"J��l��26����:ϰ<������-aJ5?)q�d�	TA���w�Yн;��B��Q�����n؝H�aX��me��W��@���:�ج��<KJ���}���;g�[��y�V  =�׮��=vt[{���"����ɓ'	     �Í7hkk�x��V�fkho /g�����w��;��*خn���{�^�P�!�����ڳlϚO�5�P��1&�L�Fokn�v�<��d�cD�����mޣx���H�/��h��t��	��P��1��sꕟ�-�'���6��v�{�^�0'������r(�����6�_�;@��& ��A� 0�|�R��nRmu�ۼ���=�
�5/x��~AJ��nE��T�u�tnG!�E,�`���8slηu����fw�r�����l���T�׻m�|+3
y���e�������v~��q��ྦ�X��o�>g�q<�Ƕ_o��ƨ!�$�������� ��(Tⱸ�����W��t��%�w�vQJzw���uA�D�_�r�\�`%�7�FO[�����k�՝�N����Z���v� 0�|�\���ԩ�ӿ���'ND�     ���u�ƍHs�[����  �e���pu��+;��vU1VXV��Ϯ�(��c�o��C�/�"
���٠}&c����۞v,��6�$=��<������������>^T�0hn>�j���3&k^b�~�j�iP=���~���f�]��� ��۾�,���~��3t�c�m�__��.ҫ3(� � C˱�y���Z[�I��.�ۃ�)�8Ծ k^�	TV�)�@E$���.���Y� X�3.�8󢜇C�Z����hyyٹϦ�򶾾N�j����֜muu�9��y���t?��r�����?�9r�y���� ��C������[�>���ǝ1�;v��x��{L]�SA�M��6��q�.P����l���Αl�].d���9�N�-��ngP�Y2�*H��uD+1�rw�)�*q|�r�������q�YA3  �Z#O�����5��^�z�     @�|���/Y���]��� ��!z��R�����+>����
/Qj�c���J��H�?0�/؞�'8J�a�sm�1g:6�sm���A�gdo�7���,�u��X��9~x�Z!�6s��������5�=?>��5�~��{~|���q�x?o&D	Ǉ=�Iy��yI�ޓ
��O�K�9ǆ��/4kt繒����B�~0�Cnr�����{�TM�~��љV����N��'��On���� � @� 0�<{�Dg�����߼�ڮng�I��jkl�
��\�"
n]@�=[��a��-Z���?�q(j~~���t�������h�c�J���b��I�j���l[��|a���k��O�<I<��x�ۣG���Ç�[�?~�Μ9����Iq�)��&��l|\!+m�*��cqC�I��M���wG�L��i-C(��BU�~�p%�r���&��z��5B�+�ڣ 	������5z��J�^�L�s!w @0��9y�N���u�'׮��Ąc�    �d`�lnn.�ܷ+c4X  �i{����X�x�~�н���A�=��:�v�j����
��be1�n��tx=Ip�=�(���3=��������'�X�",��7q�f߳�b,?��s~�,���㍿f=�-�r�𼟏�/Ȟ!�[=�$o�#�g;Ȯ;�tL��z��4��c6�B�s�����=��z�F��{���H����/krov
���
�P,�<CeI�F1o��{���e��;Oo��	  �w �P������˻�Y�F;��q�]-VS�`�\��.h7/P�0.J��T̰�^�j�}����(����>n?���ݻw��u6�x���ܹC�o�v�t��
��ysŹ������Z�b֩S��ĉt��9�k�8 �x��&b�ߓ�L�B�
;�V�]gNRb���t���[�`E�̠
����knmq��2�*ߚ���['���U�e�w�������������Յ#toAw ���f���R�O�"]�5��ߧ�=�     �4[�!�z+
��ݩ  ����<}��6�n�NQ���a�������Cu�����څ-�lwoU���ۓ�	��?�{�$Ǚ��3Gg>kK\ru��}gs��n����~|�o]_���x����0 >_����£� /k�w��~�R,wc?�����<�cϐ=B�UAx� |�P5��WL;��o��%��m��6��݃猪��"4�����c�՟E߰�*���&��V�ů����'/�K�y�n  �� ���S���pq�6kT*��"T_�=��]���Z��
T���ym��T�
���FI�ʒ`e��1&㢎W��d��:��YT���u��u떳���
^�n[|Pc<��r��N ��ٳ��,p�>�d�I�SA�GM�29�t��t��{w�lBU�Gw����+q_�~�h%ib�u6�5���]���V������x����  r>X*��G��l���4�޿O�[�     �.�>��666"���v��B  ��wȅ7*����|Cي�E�+�_�Y�+�7�y�ʍ��~/�~�=Ͱ� �☍�cLƙ��2>l���ݻ����Oq`����
5|�oYO��h~.9υc����~�;}����-�ŕ�����k��aߋ�8>�jl�qA���9�z�6|D��%���&��=J����y���W������W��w����0����=CI1o[�w�;g��[���H� �w @�)找u��^�F��R�@Լ.P�� QJּ`n���i]t�=���A	V6ǘ�3���͛7���&�y}ff�	�Cp-����xs��@�-,lq�������;}������-qJ6�f�=��v����qC�Q�S��}ϥ�����%��D+�k�h%��>��|�$T���s��󸃫����g�'��hmk�  @d��:���=u|�h�{�Gǟ^it     sVVW���t��sE��� �}�;���D;��i�Y�;�uJ��0�d�goQ��K��s�p;�t?��::�2��k�Y�#�nv���qQǫ氷��u��Cd���|;ݺ��¬�����N�7��;� ��/^tJ���;���{͊|O*��+���h�X�}Ĥ���T�;$�� ����r�w�P��W��Eo��)�6�g�����2�p{s��6���K���.5w��� �d�J �4W���ZY�Ri���.	���T�@%���`�b�i^0
��\���S���+�>(a
�U8qE+^��C�lf��߸q�����M�,NT�U{�7�M�����c��}��%�z��s��Z���Ç�E�8�j�iP]gL�*�x�@�Μ8���I&c�	����"U ��'�$Z��uD���{���`���}��<m������4M���hf  x�p�L����`I��`�z���ߧ��z�     @|�s�;��ܚ���JoΏ  d���3]��3��!����o�g�K���W{v��ڃVy�n��߆�˲}�����9&�qAs��daa��9���E�#�}��<��j5�~����_�i���~��𻸱G�-�&�����8�wcl��I��h3�n:?hLп��"�
�Dҍ��������]�Ք����y�g����!~a���ze����Q���1���$  H
� ��O/h��ڨ�hll,P��o�*g�Y�]'ܮ/R�O,J�}���{��='α4��1'��8����wC켱 �K�n�v횳��)��փ>贼s����rn��\$��{*�ɱ(������ݻGq*���]J%T�[�u��^r�+Zy��v7��mm�\gS53�VA�_���Ls��r�2�4��f @��K�U�G_9S3�7{�.�>s�&Z     ��?��)���'�%Z�.  d��w�@���Q�K�COQ��7�~��.[�9�?���7�����]�f�S�o{N�c6��cc,}��}�7d?����Od����/ߡ����G�&¯ytg�71�~��	��{�P56	?��� ��cI��Q����a�t�t���w�+@�eY2�P|W��εD�x>���m�����Xk��da��|�~6��;  p d�c9�օ-Z[�Ky�T�!U�}Ik{Q*N�/+n�݀��(ۓ����"X���E��=���O>��i�d�D� *�o�����¯����裏:��'''��s�P�8Av�q�,PKb�������E+7�޾���$�_+�VA-��}ϵH>��Ag���%���v3�M���������5�V �63�E�[+�ĸ��_k?v�	'     �h,.-���t��[�ϖ�Tp- �.�����gk�V����w���l�n����S�U�j��������q\w��8����m����|�>�d�������$x{�W�}�k#���X\�u����-���$z�Wv���A��QǦ��}/&���]���
�=oP�t���}��7Ty�&�X|�F�N���������U��>  �� �L���"=R�K���n�B�#T�(P�S������rq�+L�8a*P�"��G��+NeM�ʚ05��U�q�a�C�~��#>qC;�����*D(�)�����
��������#/a����#�<�Z������v�=��x,��eHW�Ϻp��Ztw��=\���+]�*L���$����(R����o}���zf�U�^�_ߪ  0o.�o_�R���%�}���駟}�     ���?�����?,�9!w  �"O�.�d�U����CU�=,��kn/����E[�Y�!�z�n���ݒd���m�xix�Y�m�#�8n�f���\J��?��>��g��� -\/�������_��{�СC��9���X�'B���sd�+��19>�~��9�������o{?��o�s$h��5�N�=�7l6��1�0��u|����]7��)�ꌩ.�џ/���s�ν �-p d�\n��������N��cc}��[�`{Ѹ�=8خӺ�#R�n���ĩ���m�������cq�&9���b�@;���y�ZXX�,�����Y\����l�v<x�>��O;"/Y�B[�Z�#,�6��,����e26�}j�ʹG��ΐ�h���xz�n��+J)����J�
Z�����k�������}�Q��	 {���<}�R�G�l͛��Y�����     �x���$
|���J�   kr���y%�kT/��v�g��y�����`{���������C�:x��Q�'��h�x�q��.{�b��-����$ ����Z�O��\��� �r9���,ǲ�T�]g�m�0�Yۧ�7B+@wW��c��e�a{���.��=�X�m�Awɭ�#�-���۹A�&/�O5��  ₀; `��<P�N��Z�"oj�50�7�X�k^nmW�.�ǂD��%�"����)BJ�JS�JC�2�6D����w�	���`T������_���ǯ�.\�'�x�{�1G���,p��TQ���H3�WԲ)h��'j������T�D+U�]&X�m��}�zD��
�����9�hU[��o�>H��N��"� ����2F�i��g��|Ժn=r�;v�     ��K�w�܉4���^����ٔ   S�<����^���"�Je�gh���}�@uV|nߏ��}DF�CtI��`���zV=�$<D����������o�M�����x ����_��Սxc�5��ɓN{��rQ��Ą��5��g�+;��|R~���A��|d�tw���u�A�#7ݐ;_s���*߰���X^��N�*��X|NW�LӋW��/���udS  �@� 0P�9W�s�[T]mP�\V�S%�@���_��_ZP-N��v�p�,��1*q�w�Ɩ85,��A��GE��߈�e9���G�k���Q�j�
A
�Y����̌����K��0�۹��g��Gy�>����ѣG�sl��ecvOJԲ!heI��2/L�ᱲ`�J�
�\�J��]lr��=��h����s9�h��Y�G�=������^f��z������	�Q~�{����/?����     ë5~��G���\��� �,���"=�y�j+M��Ͼ�,c�P����������C4/��R�=K>a��a�s��a��]�yjj��z�-����� �;g����_w6�_[yh.�b����w�B~�pI�+;���8(�P�?��A��ecڷ�/�;�]�Y�7l��e�X�1o�{^����Y�U]Y�/\�;G�ӛwP� �� ��Pl]�}�*���5j�>$pxAG�
j`��ڋ���`q�+T�
T:Bӻ%�>�8eS8ڋ��Q����9��R����hii�  ���#��#.Y��C�T�O>�Y�>���=ֆ�eS��r,��g\1�dl����<��{�p�RT^�tB�m�J\~P��.6��r����U���U}��x��|� -m ��^�v�H7�Kt�`�h�Ӱ���٧�6z]    �k�篷�~�h0�V����  �B�H��+M�X�I��Rh1�?Ю�zC�E��vY�]�;T����]�9K!�a�	m��Q�i�_'p��]��׿���!�����_�_������C��SO=�ln������s��
Îۘk3���8(o0ʾ�1��n�]~��d+@�J��0�����o�X�m�9o��p�t�q���x�ɭ)�����^/R��^  ~p ��ġ=w|���O��O����eb��l`W��t�T��&�_�bT"Uĩ���6�4ħ����b/���o�;�C��.mllh�Z �`��������~���v||�;޶@v<!���m�Qq�'j��q�V�Vw��{��=��+Z��D+���J����{�t�./����Ã��<� ث�v~��ߠ}��U^"�ͥ��I     r����V3[1G�7�����_( d�+ǋ����QY�R���U�X���xޡx_�z�wt�0����3I{��ld�}�tǈ��/d�������۴�� M��
����+�8Áw^������}��s�z��16��6Ι��dlZ�L�������C�O�l�v�5tV�*���M����7�
�B,�/��;�W��k����r�  �� ���D��7o��z����zbTH�=�}A��.n*QJ���j�YV�	��D����~[cm�:'�9M��-/��r����^�J�B �����=������g�q������-P��hיg�����|[�vq��hŻ5��h��T|�F
�J|<qs��p՞���p���`�]�0���>U��_��／�]ٹN�'/�_C�; {���k�����3��s?�v�i���      �壏>r~)0*�WK4[�E �_�T���7h���ry��3������E���;4)ƒ�7��0�Ŗ/8ja�4���q�iyu�7�|�	������!��=��������1\�Łw�	��C��~��I�L�XV�B��Y
��橂��Vd����5��%��ۥXM�o�b��=�0�R��'��	�K��[�
е�}��N�.^�_͠ ��+ @*�r���s�X�F;Ţ|Y���es{�0�me���┩@����Vf�]�:�>�}Y�?�c�㋋������ij��o~��!F0x���������'N8aw��_����w����ε9'�~A+������}��V�k��n�VwY�=��]&\�Ʒ���҃��w!�����w�h%�U|�W�/ܠ''�G3cT��{ {��e��ޠ��Dk~��û�:� =z�     @�۷o��7"ϯ6r���> �AS�}��.m,\�|���cI��cx���v��E����[^�0x���۞��q�eϐWyf����_w<E @z��I�������6{�����f��}�st���@o(	?�Ʊ�}Ĩ~��ؤ�����
Y���	�-,��{\y�{{�[��in����]�P��ʱ�V�n��txm������S�� �� ��9�?O_?�F�J/�.6��,+(�D!���L�T5/�*y�]�xA�ʊ0�Q�D�����v�_��W�ҁ� �v ��������^z��������/~�Nk�X�~�"�nS���?�A�������J��w�6�!��kg�q���N^����b�ΐ�tﷶ��}���]��XD3 {����ӷ��i�dv�˿��ޢ��%��     {���%z���#�竱����N�  `�L*�s����괶����+���l���|D-�0g��s�� |���n��0����4�s9�� �����������˗�r��|�3N9��Ç�ー���IK�G4	�g1�n�C���A���|�S���
���{�a�����A�>��/�$��f���ţ���1�[o  ��;  Q?U��
w���E�1G��5����m]A�ؿ��Z��k^�ol��S�J�b�D�Q� X���fA�������,� 1����?v���t��!�җ�DO?�4=��s411�kK��������N��q�+bV�B��J)X�uʮy��J�r�,�`��.Ch"X���`��A���K�.�/n"��^b��������s�֧$��^^E�C�l
xV    �=
k�|]'����ݫ  �3�Jt�1C�M�(��M��D1-�P,y��'��D����O�1��9lωsL<η�����\�š���M d��{��g��輿�Oȁw.�z���r%��.i����U�����Mƴoy��;�!���6w�TY�9����6w��Ϯ_蹶�byW�z��6w�_ع_[[�Ϗ��쑋��x�  5� �ϯ橸|�;��@�X^P��=P��1aJո��]����)ه��ĩ,�س"LeQ�⥃9���;��+���.  F���������c�=�S���x�`��?�����ZI�mݳj���V�[�h�\��s>�6��҃�K��UO��r��UN4�$M��z���L��N����Q�z���^an�@�/��SǶ�箬����|�Y)%��;    � ����F�z�o�R�,�*e �A���ҷ�Qc��J�U�����a�������ü� �Pk�gwe�;�9/�F�o{N�1�8���Ρv�>��й �����������իN�;�\��V�v���4�B��6�%9�F�"R��ܥmR~gGZ�Em���^�н���]��t�y��a�X������)���K��T���� ���; �:�r��󛴾x���r�eA�ܮ#P� ����(N�"��q�T�
�*H�b��g)Ğ%aj�v��6g�x���B� {�`�+6��O��Ot��ez��睶��~�����f�=��i�)dE���Pq���ݑ�:��ab���� l�if�������y����w����[<Fwװ�  {�?,�љ�:�����B�Bx�]z��'	    `/���~��T�V��c�W�����#  ����g��h����l�lnW�����=C3�PԹt�C&kޡ�y&���?��q���+��o���y��/~AKKK mfff��������������}��_�'N8c���G4	�:��<՘0��G�dw7YA�x^�����=��)��o���,]�Y���s=���c�ze����	z��AZڈ�b `4A� `��
�ľ9�.mP�<������۽K�T��vUk����S�~�	��]�J3؞��d#����:������4==������ ����wy���t��G��;����äh���ߦp5�}��b��˾���Ű�x$�s���*�.�w+Yؽ��J�ۿN����  {��������OߺX�r~�L���m�����    ���no��&����8K�^��O��X	 0��(���;T[�SylL��cu|R�D�C�Ȅ��M��$�؜g�/�Q�۞�?v��z��W�@;{���nm��r n�u�W�~�嗝�����B,.���W�BgϞ�E�P���bV<��-�i߲7�+��[��O�
}��&m�=�p��/��cuW�_�_C�
����3\Y��[�?:Gܯ  � � ��/���i�n}w��T���=\�R�f������SY
�gI�JJ�����z�~���:������ �˽{��?����p��qG�z��gk||�cC��#j��oK��j�]ܗ�hE�%�^��_���;�]a�#^u�)��W�`�����x	^^~�;��m� 0ڬ7��ʽq�����+��u3���>o>��C    0��縷�{Z�����R�n�� �oN�*S�,�P�j���W���ڶw(jZ:�!pg�x|{)�>(�0���͛7�P�3n�  loo�k���l��OO>�$}��_v�|�;.�@��~�j��$�z���]��+��u�܃�����r�^)V�z�BUΪ/�.��s�6��v�.�L���W��c�g @(Z ��Z�yp��+�(W,�>�+Z�c
T��3�*(����/V�Mq*�`{�ι�B�w����g?sD����#� ��~���o��lG�q�ݟ{�9'�>66�KR���?�j�l��m�V<�=�c\QJ%VqSu�iTb����to��*��!/�U��&�6w�`%�V����3��7˴�2w F�{���8FOߌ4��kלא��I    E�p;�qp��*� ҧ\$��KuZ_��z�2�0�?W{�}T���w(���+>��C&-�0+~b��m�;�o?��cz����7���S�%�  q������{��y{�ᇻ��zQ��#*��8b���d���ή^���;����t�A�0�Py��ks�b���������?n���D��� �X�ѷ��h�2O�R��v}��]>0L�R],�m^�^T�ɒ85������8��+J���?����t��]�� ����B����lǎ������hיc;�v���&ъ���w��E�J&V�53�!��@�W��k��EcP��Ks��3��'��2� u�[,ѱr�.����ǟ|�Ρ�    �_�p�}nn.�y��<�:7�����   ��8���V����w�J�t���������۳��I��Ohc����s�����_v6�� ���|���������裏�/��x�:a���B�~[~���$C��8ct���� �~�f�{P�]'��^��"�j�g�5VP����]�ޅ#����4_�/���A� �+ǋ���UW6����*G�*���*�p��8%knW7/�E*&-1*+BԠE�4���n߾�R?�я�
�  M�������ߝ�ĉ�o|���~�i�=��z��Eݟ�p��P��/+��qE)�X�ii �Vv�  ��IDAT�'��A'��煦v�A�����[U�Ly�&�]�7�D� ���6�����t�M��&w~]{�G    `��ro����lno�����i��p;  ]��(��۴Qkt�C�K�:R�](�����a�ޡ��ݽl�=+a����:G�9����*ϯ��
���� ���/~���q؝�P.��ַ�E�ϟw�������uΑ�����h�Cl��Dާ��뷹������ð�{^�N2X���-��o���nЍ����9x� �Up D��tb�&mmR/�..%hԾ���Tr��w,H����$�a��j�v����g�(��o:�> ��g�L��(�{�5���	 �'>|����(��SA��G�����9�P$@Y������d���쓙��{f��_uWwUuUuuwUWu��y���j��!�]}����imm�C=��~3gΔ��g�}6����v�WN�Q��[�1/�V�뎴H���L�J�msM����|�lAw���!w��9N7�7���q8�bbo=Ο7OփR��_�^�W��g�Q��n�h�`ȝB!%�n�݂��������h���B�əs�v6a��Wc��ڮ��Y�!�������;tr;�+���Wnkoo�ڵk��/�7ޠH):�ۑ��w�u>��Haw�N�0Aڧ��r��~a�s8y�ۡv+��#_h�A=��ܕM�F>a�����/Pk˱��R���m��%�b�P�̙����K�H�wBHN�@��u~�5�����d[�]ZAe��,8����H����E*����^���0%�`͚5RS���D@!^D�n�ڵK�.��wߍ�?g�u�v;v�����\ǝ��sB �C��ҳ!v�wY�R�U�&w���rL)L%<�ĵPF;CR�ʧ�!��L��._�E�v��yS�ĎJ�|%�x��A?���W��"���o]L�-^���?�B!����������V��i�®����
��pN=�{��H��9�b�ǳ�bi}B����������[�ͼC�1/y�v������
=__֭['c�������g�7�|SZn��v�x�8��Sq�i����Z��K~�Ѹ�Aw����b{�F�����{:�.y��8�*���"�����1�R��O�_}M����u�k�h��z��͛�U�AD��R�P�"�X��sg������q�r�n&E)�H�mZA�p�^�ݯ���LE����y\�c���l\�&��[���ó�>���BH)!^�6m�$-��v�$^�q��x%ޓ��H���C���0����z$-R����(�ܵM�JqJy-��������u3q��E+����q��Qx�k"�t����r�m ���q���k@~�عS�0�/}�K|^$�B)D��[o��C�|�;+�Qg!�XL���ûn�DeeeF)��G4�[+�Jl7���;tr��ٱo!����ￏիW�g�AWW!�����J�K�妛n��e�/��^(�n��h�ioPw�Wt�C�v�g��^���/YP\�������E	�I�PO�K�+z�2�s�5����}?��WZơ%̔;!#�	!��1.�ϏnA�#��V0ש�vՔ��Tb[B��o^�
TzA�l�T�H�/L���mq�k"T������矗D�>� �R(ū3f��sϕ�$�����[�r�E��g_/R�1;E�|E,���9 y��)������ٚ�E�!�v��z������p����)3��@���dO8����¤���q ~�?�a>��Ϣ"�E/B!�/���#��E;l���	ack%!�X̟�Q���=Iy��J��}D�p{01n��۳�����u���k̎}߿��>��hhh0ܟB���RΊ+���#���B�N�6M��_h4^���H��=C9���˾��K�ŵO,]�������g�cY��f�ֽFS����n��>��F��a�tl9Hϐ�� �?%�ٱ����;�.o�nO/ZqJ-T�R�q�0e2��@_���y��Av/�Zv��9�)�D��$��;{����%K����]j�=��p�9砦�FڞK��h�T�+'�s����O�H����+��63��W_3iŪt;C6a*�%c��hӢ�0g^jb�;!�J}W�C8n|$�sttvJ�����gQ]UB!����ny��w���#�����`�R,N�DEg�w��f+�2��ޢ�Y���C�z�N��>^�c_+��/\�f^x��]�V�!	!�\ؾ}���u�]8�䓥��)��"�w�������R�՞�>�d��XT~a� K.ǒϧ��c"̞��!wq�<�Ae�ݤK�W�n���s���AB��	!��2;�Q=M��3��Z��,�^X��xZA���D)�"�aa�v�Qn�S�"B�+L8p@jj_�l��$����x-ܴi���~��8��3�`�w�q�v+�s��R���;-Z��k�;�IY� %�*E��$V)���T
V�qy�AI�RW��V�\E,�*�ш�G���� ��!�ͦ�J���c�zuww�7��g>�i�7�B!^c���x�������h��5�턐"��pA�0�Z2��u|�|�����:�vm��o�?,�whe�b���<�Xcv�ke��?��ڟ{�9����B��Z�E�L�<Y��>�l̟?_�^�_h4^�n�y�C�z��U��[�
��wU�{� K��jW���69ܞ����^w�p�Px�Շq���x�abfkBHy;!D�/�u񋂶F��T��ve��,ܮ/N�:���I�Ȑ��o^pJ�*���S�g�І���W_}UZ���Dmm-� -�\��(�����i�o�������k�;p7����/�h?��7��9��s���{�߽���駟��c�9F�D���ژo �h܋�U�������z⧾H%#�U�v�f$���V��,m�f�I낕��u/ϝ�'wՠ/�!�o�T�?�G��?�>00��o���=3f� !�B����mۆ��F[��1���j��Oq�ʠя����J���ۥP{.����XZ�0�;4���7��x�}�V���/K�����S����Ŀoq�nyW��ǭ�v����/nݿ[�]~}t���}������wn��)����#�<�G}�{�t3A�3t.��sxe�Kb.��|�6w�����BEA���n���K�����mۉ��&�U�g�;!e	$�jv=mt��Z��4ܮ����3��J�J�0���*�(��ҋx���b�On
X�8W1�W�<xPjk_�r%v�ܩ�_�[	��p�����Ŀq���n��倷S=�[���������bq7����\uu5z{{]�!@	�ެ��ߖ�;�C
�_x�8�裥m��rٷء�\��C�*D�R�k��3"[3�hqO��SXv�*����t+��u|�B��}��i�;Zp�Qx�s"�w�xH�>lh�B��)���:N���������ı��f^B!�D�ܻ�6���Ֆ������Z��	!Ea�� �c\+��=��v=��4�nnϥ��?����&����� ��B�v��F㍍�����-�Ο,qK���N�����n�	�~�n޿|�n����w����׻��>�m|���,]�_��q�H%Y���l��ʘ�=D���XMl�I�vQr����BEA����,(�����%�Ik�B���Z9��E�z.�ނ��+���%�b,B��	!*��&�!�ѝ)P�uY��n���)N)E*��9O+(���Lҭ���܉u���w�b�˩��q����{R���'�p-PJ!�����N��E�p��K��VD'�q/��>�n��.KG��wY��^_�V�Vs�*S���'���7�j"������ ���u鍃���o�]����ݻ����O}��v!�22����;7ڦ]vGEs{-�n'�8�ѓ�8&�/��*bc�=�f�˞�<����2�C=�{��Nzy�l�����,ϫV��o��Q#�-��7��[�L��Э�������oír&���Xܺ��ſy�f~v�o^~�s����wss��>���8餓p��J�wYK����e_/�ڕcv��Ny��u��D�=�#J>���mj�䰻�_6�0�B��n���}a���_���)�oc1!����'B{�o�QC�J��̈́)u�]_�Jl7��ە��l�
j/hF�BP��S�w/W��E���?��c�裏�A!$;�5tÆx뭷0m�4,^�Xju?�ä�N�Q��[,A��qN�V��XZ�)!PI[ �����Vy
B�9�D����"2�L/�P��ʢ	�+aF̉5b�̹X��!wBʍ�+#^?X%�|�U��xk[^[����'1i�DB!���{�b˖-�)��%���բ��vBH�Ҭ F�w`0�s(�H���ci�C=��)���>n�K-�ng����R�],���!��_��^���ӧ����1u�Ti{�~_.�s�n�ѩ�z>��3�
�_�hqG,]�%����_#�Ψ��,����k6��z�a�������~�;_d"����/�ab�F�5�n$NIc򔂚p�R�?z"U���B�L�����Eq�+�����'��چ[ZZ@!�>�k�0�o��6�u�]8묳p�E��c����)F岯ۡ�B�qC�R^%�䰻|;-`Ɂu�Vm�]&S�J�_B��o�5/doeP���!�q=��`�l��!�����=P��$`���BH|��n�\u�Q�K�B!v"�A�l�jk���ߏ��``��1��9g�hk@ ��s
��gx���{��b,m�ݨ���C����8'���W���b�
�K�dB)�.Y���sN>�d|�k_�g?�Yi[�~_.�k̮0|�=�\�C_�����м��ωE��5K.�X��aΩ�����A��	!�@k��/d,P�"U���`%�����b��0��RP-L�7/���d��8��0%��[�⩧��O<a�T��B������+W�s�����p�gH��v�Q�_H�]9�h冈�����!ټ ��}x8-^%�k"�л:�'XAլ _n���U�N\4o:V5�fEHY!��׷T!�c��§�mhlDGg'>u�񨪪!�B��tuu��M�l�1��xy"�B&��Do�^�B��Z�P�?��B�o(�ە�X����R�2��:���
�g�H$��_~�?�8�y��}	!�������O}J���ϖ�3K5���q���]W{���ͱ���/�z���!���ʠ�O�J�6��U�a{=CB��	�|1,�Bo�ެ�
Zm_P��+��f"�6�nl�N5���n�BS2� F1��Z�^}�U)`���S�"���o��&6l؀�K�b��Ÿ��P[[+m/DP*��\��fc^�����ar+���XFSʘG�p�|;�8Y��.\!C�R/}��p��xf�tP�"���ack%�)�>��&���v���8v�����B!�"L����uz_Η��p�`��vB������)]�m�DEEeN��LQ��]��R���!Z��B����u'�)�X�}�ϫV���C�0L!�8lڴIZ��n�/<���1~�xi[���BƼ�!�)沮��^��M�,����{�/�Τ�+���2f~V��H�����r,��U���;�<���̾��	)ap'd�R��_0�=m�����Ys{N��S�M+�c��B�2��70�nwB�rr/��f#!J=��صk!���x�&���I�Z�`.��L�2Eڞ���˾�KvWLѪPQ����Ou�]��'��A1�,65ԢR洃CC���J��o�.Xi���9y��O@Kx���bkG�Ըr¤!�t.��&�U��ۇ;�8T�?B!��KOO6�����n'M�!�k��V!�8ʌ�A�0� z��JcUh�J���?4���v�3>�5�gx�b��X��>�бl���ק���}�B�;��-�܂%K���3�ĥ�^�#�<R�Vo��1'��vx�Ny��!T���^H��b��p"쎄_9�	�y��k/m�=3������ϰ�_�4�u]�����!!�@D��W�t"�ѕnn7jp�&Pi�T���i�]n��(��v�8�Ǵ�� >9%`�y��c���X�l{�1�Q�H�"��.mmm���{���㬳��7���b�B�]����dv�B���x���*!@�1u�=��!v�d�d�]y>=�*-<i���6�w3���~SK�����?�D�^�44��R^l�@w4�/M�E�������x��������̙3A!���ScS�o�nkk��t��#�w��%<B��3)�#�{��B�F��ٌωu���d�]n�6�Q��p���P]�0Ҽ�|���\�����aThѯ�?��;$�� >��8�S�}'�p���KAw'�󚇘�zbL��^!�Q�P��:M�F��2�.�N�T0=��I�azh����[�������G���!z���"�2����h_�P�S:B��@��T��n�Bf{���v]q�`jA����
�{E��ul�Νx��ǥ?�p�BJ���~�\�O=��$\���O��ҶB���Ɗ!d�-Z�+b9�.�zj�,9�nu�A=�JtO�.T��:��<ON���h4�c�0f�,����!���� ��S�/O�Cm�� �x�x����b�1Ǡ��
�B!�m�[��]��z��뛫��!�8�	�C8|`��`�;4��9�7�˱�c������v�{�nc�q����b&Hh���q�FB�.�5���^5kp���c�8�����^�C��1����Ct"o�g�����z��XI�P���2�ҷ�o�K��u|�t94��ar������i��q_��ҁwBFGM���D��^�BrL+J
T�i����a��H���'�&���T��v�� ���� �����[��_���~�iD"B)M��/J��I'���.�H
�k��*�c^�����ldP"�Q�􃪰��\�E)`)+e���P2�:t�ԏ�D�R�+r��߈Sg���;r'�������:���^���hin�ܹsQWW'}>%�B�">kl����;̾���a^�W�����!�s�Tv5����|Ck3>����d�]Y��m�g��v�o���q�5&�w�Ԑd��\������x�������>K!�9�k��M��y�f�J�-��ŋ�2m��X���9y�Ӟ���ɞab�gy���e�p89�s,vGRK7���-��{���z��k:���j����}�8e��Bϐ����!#��MaR�}�T�B���L*�i�D*+�٧��8Ԯ�X����S�8}\>co�������_O��!��>�p��oH_��Wq�gJ� n���R����e�J-V�S�`�P��)��T�)*Aw���>aʗnf�*V%O�^�Tj��us�LC�-τo�7����jp��~�eO��P�uN���ߏc���ĉA!�"���ۇ?�ȑΈ��Aw�_�#�8�9��5mM	/0�V�ܳ��,{����nm7.Ʋ�ڮ�U�a�7�ԟ�ޡ2��-o�M��+~�<��ݍ'�x�<�����`;!��0�5���7�t�q�s�9��׿�ѣG%�^��Ӟ���i=Cm�]l�%���ɰ��Ǭ�]q6U�]Y����Ҟ���R�]�J�DPs���;O��3$�`����is��l�_پ���njOߖ��Z�*-T�C��"�f7�ZPG��
TJaJ�0��b�M^��l���{�n�:
S�R��Aw��p�����K/��+���jW�3�nv'֍�VP���b�[�5Aw����h�ܓ���zPޞ��K73����Ī��1(�Gښ���XY��C)+�}x�@5�	��I��ϐ��7c�[oa�ԩ8���PSSB!��\:::�`{gg�#������*�چB�$��aa����6�[����o(ƅfTh1��7T������=�S���>v�m����>���﵄Bʋ���q���htA�q��Iۜ��<�����5��P9��3���٢��.{���U3?�!��w�IԞar�h[͛�"�����x�	)s��!kSjo�
T��v=�J�r�ũ���B���^w�;�3�ƍ����kײ��BF�=࣏>¯�k�N"�p�B�ڢ�Aw���v㶈e�xc�F�Y�}+�úR�2"q?���5�,2%S�F�c��2���sM.}�{��n
V4U":Đ;!���C��SzQ��o|���8x� �O����<��� �B��A|�m���8p��#���Snn��֎
B��T�����֌
m�]��}�g+�>�cYmmW��V�C�Bz���c�q�1l_�b|�AǾ<F!�;����%K���c����7��ɓ'K����<������(y�g��q��(�cP�"��2ʠ{�3����B<C�7T������s'c��j�3$ī0�NH���/����m/B��a�"d>�`�H%R�����d&P�S����t*��R��<N˫��*	S������BF.MMM�����c�IA�s�=W2ќ�{I�*�����K:�.�Ti�JZK�R�r�	�ʟ|���ޒntW62 }��H%�M�S�U���	�K�K�� .�5���FO��Rn4��ԮZ|iJ�����Z���{�n)�>{�,���I��	!�R����c{}=����H�]3�Ԡ5~C!N3�ʏ�L�D��+nO��z�XٽCm�];볱g�-�n��g~�ȼ�]��Wnޡ���˗cٲehnn!���šC���O<!�b}����.m�b�]9榇X�u�ϗFlO�) ���Y�&��F�a��U�=�{S������ �тf�ó���� C�x:q��!A?�hN=m���4lm�2���4��`��@e���hzA���4)2��9n�On�Q�
�oذ��?֭[��C!�4پ};~������D+'�����cgh��9�����C��^P�v��Aw�p5��F���L��K	U>y0-bA����)D/��!�]�8{J/��G{/C�~����v� ��/~lcpp��سw/�Ν�Y�f!�e�
B!��җ�w����l���A�o�����+�b���~|aL3z�����:���w(���g}�c���skn���ڠ�@ֱ���R��u�|���\��=��n����ւB��E�E�D��q�%���/�)�n��h��Xщu+���3�%���>C�jʱ�H�w�3L��H=������g�pO�D�7�=ԅ3&ⵎ�h	;�B�wBʌ����A��--Pi�̦L�Sr��f�JG���g���� h廏ǭ]����?��;�B1cǎR����>*��?�|���K���}�Z�{���'�ԍ	�J=���F9设�3Z�t�Hn���r��@����RjX��p�<ak��p���!��p��js{%������}Sa�YD���?DCC���~�GH��	!�R�����)�YU���d�}(~Y�n{>� !��Yc�L�D�R>a�A�ݒw���YU��1��j�BM!V�w�?�`�{�N��<(��)t���B!J����t�R�}B�b]v�e�Aw;<�\Ε�>N�����ʞ�hlW�JQ��9�jʱ��X��7Ty�r�^3���3����@__Ż����Iϐ/��;!eĘJΚډpg�Z�ʳ�=%N)��	�Jhϯ�={�=S��~��NAȋ���)�}6oތ%K�`�����}I!�����K��<����
�y�������r�-�ʍ�|.��b����ˈ}���Sr�A�h���O��.߇/pGJ�ʼF�^/*N�neH�����I��cchvv�R~����Z���|b\���G"l����0��1{��esB!��"l��؈}��K�m�D\��~��"��R�Oa�o���b,y�F~az,fן���b,S�P�!3�T�ޡ[��w�\�Z[[�f�e˖I��B�"���`�ʕ�袋p��c���ڕcNy�^����!whf|V!��=CM9,� �<�fN?�g���f���o��3��(>U���3��!�0�NH�0�6�S&����G��]!V���n4��_h�G�Jl�Ƽ�]�%ʋW���zܶm�p�}���g�u�ՈBH����������K�v�Jp�%H�c^������%_�%G�hgPW��(�jdPݡ�g~�1[��Zp�E�T�]�x����/� R�G�*��z�L|D����d(���vk����}�
������A�K["'�D���q�@!�����&��8p��Ҏ������+���R�i�B���Oa���12��Y��c��l�ܮ�e�p1	��}�p�t+��iuV������l_[�b��ntvv�B�t���{�/H-^�W]uƌck��b�=E�B�ꂩL��'ƒ�v�c)=C#����ܳx�)��Z�]���#����Ĩ)��� ����RL��G@_�?մ`�ڞ5�����H��E(m�]+Z���:�V�R�ڭ
Tv
F^��&N��;v��C=$	T��B��>���J��?�y|�[��	'� m+� ee�|'�sc��+�� }$�-�FM�]���ވ�lrԁw_J"S�2h�Q�=��!ZE#�ۉ�)��� �m)Wv��8�s>9~ G������x�ۿ���;�f�����s�͂B!N"��&ާ��+"�WZ�x���lm'���f�pXo#|� B��v�+����`��l�Y����:AwA.ޡ�a�R�
������ᩧ������c�BH!:tH
�?���R1�%�\���*GC�ʱbz�v{���y���I�B�3�Y!�2H�lrO�z��r,�P��v������F1cp*������	q�	)q���o�{t���L�ʵ��,�.S0loO`��䤸eǺS�仏<v��A<��cR�]U�B�S���ذa���/��k�����q�)+�"0��X�v��c�@{b�ئ�����>ԭ�6w��Sb=)V)��uE+�f�J�J��&T�8������r%2�hs����1&��LT]]]x?�l۾3�O���F�!�B���L��с={�J��b�D)�;�k��ǝ!��j!��s�� �5����WhWs{�7L��[(Ʋ��5��x�Z�����R�#�^x�,]�MMM �B줹���r������&.\(]�8��c������g��G�Ɣ�r�]��Jݳa�3L]'����}��P�T�6��g8��'Ϛ�Ww�3$�Mp'��9����vb0K�٭TF�z���p{��y��^�����⒗,yLLu�����.Z�!�"ރ֮]+���;�<��}ƌ�6�)+��+0��Éu;.�c�����p����ԃZ�Ji`-ɓ@ne�АR��6�'���@�'^!y��x��7Q�"d����;kp�aQ?~ �95���/hhl��ѣGcڴi�?_R'�B�s���c߾}سg��pQ�{ooo6W�w��턐�r�\?�3>�cYmnW{��cY�b�c���Xwc1��s�=�{������B!v�{�n�x�X�l���J�y�O�9��>v�ԋ����h�3�:�.��1�=Cy��_��ͼBs�0���|e�\<�T�/�B2a������B��!�����*k��Ԙq�L�2��:-�y
Tv�ӽ���1��#B^+W��ZD{;!����hŊx���)���
�;֒ؤ+d�BB�F�(��]/TВ�ݒG���XZ��1m���he��u��~�ޗʸ�����Oq��ٓ�U͡�9w.�k�`EH93����Q��� >3��k��b������m۶a�I�2e
&O�,}N'�BH�Y'��)��;������Nk%���~#������M�,�C�����;Tb��۵��c���~�_����sz������n�:��oÖ-[l'�RT>��#�p�R���W_�N8A�'����Ct�+ۺݡ����Ҙ}�a:ܮ�'�f���|FAw=�Pڧ�	��;��A)>T�)A�03$M��0�n&R�n�M:B�Yk�=�"\�	�	T�$Hy=�.�5k���;�����A!�xѸ'�V�^����
�-�<�W���i��m�PAKO�I�	)ޞlk�L���[m3L�U�kE��ӂ�<(�82�1*Ɣ�&�>�фs���
V��;�"~��W�)5CR���
��"^K67K�x7n�N��)����*B!�:���hniI��;;]	�E�}x��ۺ*�@!EE����uO��]'�n)�����F�X����>g������������w(<D�	!����o�--g�u���N�%�.��O1<E/e��[L�P�/LݿOn�J��~�ǩ���ޣb<�ڄ��ƪzB�'��p���Z����70��Զ/�E���JY�*��iqJ�	.Y�/��2�)B!���������˗���/�9眓�����v�}
	�[=g!��v݉лr��X��!Mz�L�R�G���׍��>�^��L�*�T����H[Ο7OR�"dDp�7��w�b��>=1��@q��"^S;::��>���'N��	��~��>!�22D[{;�Z[�`�����f[gH
���;!�n_\7�޶}R�]p�cYnn��+ƒ��,����@�ޮ�r���J�;��y�%�~{�}���C$!���}�Y)�r��[��&M�d��S���!�qL1֋Q���&Zܡ�p�Pymh6t�ZP�����,����a�m9˷S�'��0�NH	q����4J��(e RY�������)��*�(7�\�ٽ{7|�A),�FA!�x��%��������xu�5��㎓�e���c�1^Y/D಺�Xb1Y�Q62���Z�J�v��Ku���6ܮ����}�~�ί�˷#�;��@�B�5vW`w8�O����"�����yV,����_#�O��	�e��ц_�!�Bʕ��!tuu���M
�w�o�]�!Zڛ�Cx��=Q�ۄw����Ds���gh�ޮ;۳%�P��=�Y�Sޡ�oX�wX��u���屾�>�\�w�u���A!�x���<��#x�p饗��_�:jjj,���C�3��g���{�"؎<C��'� {��kH��)�к�.=��H����{pѼiX��B���a������ATjHNaJ+RY�ZP�����*U�ݧ�2o�f���d�8���H��M!���l�ڵx��7�x�b\y啘2e�'D+7֋�Ġ�&��#�+����S��<�,ZeG�ϐB�J,CCzb����=��m���ۢm;�p�l�dȝ�Ct�'�>��Qc��?n��Aw�P�5R4�E ^+G���;cǌ�رc1j�(B!�'�]Gg�l��pqfVɆ�����Jb���"n�;�����B,�`{^�a2��K1�a{��o(֡l��*��ipz��;��>��e�=��lojj!�R
������oǪU���o�w�#3@�b7;G�x�z���S�0���ɭ�x���I{��V�t�=��Y�T�]�˔ڟ�;�����.����!e	�B
�wBJ�S���K��CYE����S���օL�*o�J'�nE�*��� �A�h��Y���z+v��B!����<���R;�W��U)�^YY�x���rib�g���xZ��i	E�{2����Ҥ^ =q��(�S_��B��\{jϭZ��*��i���X��84O)?D�}kG���C~�Dk��)�d����Q�0j�h�gm|?�@!�xd���AOw����� �F������Q�C�	!���-�A��`�7̘�9��ڬϙ�a K1�ٌ��|��v�L�ʱ�;,�w(ظq�ܼy��q�B����_���җ����j|򓟔Ƴy}V�)$�nt�z�V�5���3�}}�=C#�0��/��#M����<�wʵp�>,�7��+r'�ap'��|Y��5"J��h`�>�`����˜V�	��+��ħBαm�6����k��Fq�BHY!f#���;�������SO��R])6/d[/�(e�ob,&	S��	�J�"��)e�J�bג:���U�X��*�J�|��a�V��zp79˷3�B�Hc`ȇ�����uc�8f\�Ao4Ɋp�XZ��T�"�.�⭮�BUu���Z��/r�����BH��W�Ed���ߏ޾>�ŗ��O�.�{������a���vB����sD��9~M_a:복p��w���V�enW��3��)��ɰ���|�)�8p ��s�/_��/�B!���[oI_�:묳p�5�uh�=E7B�����������J0�������ˬҧ�~�����X�X�AoX��%��aΜ@��	��~k{���jZA�Ԃ�)��
i_(u��Iqˎ�B�S�>�����?�)�K�BH9"������ӟ���~:���:̙3�v��.��f7C�`�)���u�p|!R�53���LO=�^���
V��2���[��yӰ�! �q����ht���Ǘi��8�L�����&�(�Yg������!������Pb�o�|�VW.�>�Jߠ�UH���a�B�A(�Å�{�h�hm�m�gec�v�g�R,+3>붶k
�|I�F�Z����Q����������$!�Rz�Ϧ+V������*\r�%	�3�h7=E'C�vy��mNz���H{�iIZ|>�b�\��d��g_:]4wV4V!ʐ;!���;!�̹~)ܞ���ۍ2�4�Z�xzA�p{	
TnNn	Z�iᩧ�½�ދ�;w�B)���X�n���
\v�e����Ip�Ǌݼ�m��M�u���)��آ�R�:�9Zt��P����C�]�ʅ޶}��n�7�8� !#�7���UC8z\3k㟉K�5A|V�h�%�B��}~l;T�]���g�	!�A����EOgk�3�!ܮnn�ll������b�5��9ﰜ��Ny�bٰan��6|�� �Bʙ��6�|��x���?��ϫ
�����}��;�^�л]��2�;i�0�ص� �(�p{.�3	+�r'�	p'ă�57��ܱCՠf$R�O/�hoW�TÀ{b���<*P���U�9��}�����͛Q%���/n V4:������s��_��_YY������n���wYXw7����/�[���7p�o^���^��뭛�]6Դ�߅�������o�s�Q�V�C�V��d3C1E)���z�	�im�r=�\z��*��0�}P��>���}XĐ;!$Ns ��Q�a��(�����n�%�BF��}gO��B�@!^�*,�ٍ���W�-��^��p7�吻�Y����*��"C�)�8ҽCyl׮]��?��g�y�_x&�2b�"?��}��v~��`֬Y���͎qc�X�w�=C���Xz���oh�/Ly��s��c��;e�w���#&bծ�3$�Np'�c�3ϏXkSFS��p��@�
��M-�k�B�;xU9	Rv	Z������;���)��O����ߐ�o��n>w��C��u��uĭ�����_{ܺ7����/�/F�߼�Ϳy�z+���{(n�׈�{����o~��Y�����1{��4/����(�z�E�l�I�#�|�F��ɠ�I���he% ���D�R�d�B�D�}�~�BZ&Ta�بx�wB!�x������� �wW`_O�m��R�c��C���0�s�k�Y���C�Y�M}C���^�{q�h���~�����?����ɭ� ���M�߆����ߞ��!����n޿���w��s��r1���.^o�,gr�o^~�+h*#�o���v���R���K/�%�\�����>�c�Z/ďtr_'<C�|��Mg�2���*����Ý��`���Uː;!6;!�̹�ڶ��@����&P��N-��Yim/o�ʫb�v],"���?�	{��Um�
��"�(�틍���p7\:���.~�n�]��w'�n���Y�y��@��ߝ�_�p�k������n����_ĺu�p����+�,X��[�r2_Q�l[�x���&!b�CFm�z(�7�
V�F ��X4�A���! =~B������JL�ƬQQ�3�J?�(%�B�"���}~���t(��a�f\$�+����gd���b�Bʦ��r,#�0[1VF�]tOl�¸K���-�ϫ^�޺��r�-ضm��.�������pص��߭��Þ�Hn������^�(rӻs빋�b����^��x�q+���߼��+�d�#�o>��x\����SO�G?����/J��}f�pb�EY����5�2�|=�Kم�պ���y�;�p��V�EĽ�B�
�	�g�"�ј��	����f�
Zi`�/ 2��S��g��xY�r;�n����؈[o�����kafB!�"�%K��oHm�����Ri^Ю"p�)J�G�-1&72H[��]ĺ��KL9�mf��(e.,)�W�c��'r_|�,���	!*D���? -ۀi5��UŌ�AT���Bq�����A��	aO8��!^�BJ�P���z���+C����À{��Xf�v�w�Y��_)�ם�<�;�C
�U�B!�x���z)�~����.?���B��X)x�V�U���>����%�Վ���X�T�(�n)�	� ��	"d1�n��@��,O-�g���*;�b�O��ŷ}�-[�;���� �B�5�lق뮻N����ZL�<�s��u����d�*-ɂUb�4�`r�Rm3�פ�!��Q61Jo�\X7��ݙf��}��/u"X'��3�rSj�0�:��5����wB!�z���ā� ��F�j'��"�~�lno-0ܮ�j��j1����澡y!V�ޡS^9z���z�����_����fB!��G�X�B*����q�EI�>�������d >�3To��Z�3�B��̛�=r�&������X����R��2'DeW������A�)e!J��M+������/RNPv���書�����B!�#�V�=U43,X�@%�h�y�\������ے{@V���É��m��h��`%o7�ޏ����m/9˷��AI�W�����l�@e �)ՃR�}R� �V��B!��	�����d�]�BH���p�~��[S!�\���`��+�#,c����7t+�N�P=������o�믿B!�X�������W^yE���c�)(�.�y�#�z�Av�mj�0� K`���8��+T��S�d�m_V]4g�7U1�NH0�N���:;�����p{�Ԃ*aJ)Z��T���X�B)Rv�O������׿�U
�`!�B
c�����o~#�V?��1{�lǛr]��(e�o>���<�_B�J�++�E��`�Ijj�*X�#"����Z�\0oVՃB,30��Ξ��*�1L�a��R=�	�C�c �BF:�+`~���P{k���ka���@���EnoI�bn���cۭ��Fޡ/��;���z���p8���_Z���@!���X�n�}�]\z���w�����C�'<A�z!�3�nt;<Ch�ܕ����7L\������ʽ�6�h��9S���C1ݽ!Y`����Ҭ �5"h$PY
��/�n7�Z�����N^�
Y���o��w�!�B�e͚5ذa���*\q��u�SM��{5�^�6��2������lj�$X�MTc�w�e?X�x�Ѷ�8�l<ɐ;!$O"�>��V,25��Tc\��WI-�����8!���oȏ�:#tE�#b�?�b�Bʏt��9=�M��Pr�g3��,��=BS�P�g�`��v1�����:��~�z�t�Mhll!�B
�����s�4#�(�:餓��|���1;����b{�v��9y�����=&�A��3�e���a��=���h�T��>��3��	q�/�aTw�$*�M�zU����������1]a�R���������tHK�,�c�=B!�8�h;3����O�Su�Q7-�^jM�nK��=��_�`���`��~�k4hדc�Vr?O�3xJ���A_|	�@o 5&��C1��Q�/��z�vM�g�?���B����P"����3�O-�h�gԇ�0�_B��@�R.�BO�A�7�z��<��!�h��a���S��a�]�z+�^�av�zgg��c.[��3>B!�m�6)�~����Ø1c<S��]/f��u��3@a��*u�(�Q���h­�pѼi���Rd>7=������4�R��n�ҋ�4ܮ]��)Sz�}�X���X^z�%�r�-ػw/!��<������·��m�����/Gee��"�v�Q��<�l3���	r���Ա|ꛚ�1��PmQ�i݁����S�4	!�0����V[#��*@����z�c�m��g����U�B
g0��4�4k#C�1Ѹ>0_��?�K��uB��I��C��K��k�Ê��!��7�l7���0ܮ��Y`�y�,5�P�ꫯ��#g|&�BF|���G�|���G�җ���KY���^/V��}�0a��y��� m�y��g��:���/�7˶@���OOab_#�`fk�B�2�����J?�S������R�������m�݆g�}�4XE!�gm���_�6w!Z͟?_��	�)ۺ�T�籲My��`S��a&V��V��i~F�v�̹s�\�!��}���sB!�B��n���&�a�����XJѺo�_�%p��+��S�b�g��Z�
�B)MMM��O~��~�����1~���ci��#���~�P��{�1��sG��!//���Z�bѼX^�iW	�
��OLaZt�xMR�@��n0�H�K�=-V��� UB�v/
TN�SbY�z5n��V477�B!�"Z�����K/�D���*GE'���b�RV�ɂUz�A�
�6���,d�~a����۱�F�2���!�B!�B��º�nW5�+�C�ٞs�g܍��f�a"�.}�������_|�E�;ܳg!�R|D��#�<��k��?�!�8�U�*0�z1��J�3�b|Xnp�x�>��Ɏ/�Vk瑯��G*�Be9V�n\0���g�)!V`���"P7>����Č(���)u��3E�@���Xe%ܞ
�g��<��	*ۺhmS
�Y�&34E!������=�܃w�}?���t��ˡ�!����n�Jy_Z�Y�J��vYf(X�o�����s�~C�B!�B�H��y��q��Vh�B�vP^�%ܮ_���!ʺ���v��@��׳����`�ҥx���B!`�޽��/���>�_=&N��I��ʹJ�3��"��T=�P���5���ؖ��=fҊe��,�_�uέ;O7𚎐l0�N��L�ǿU��`t8����^�H�R�ۃ9���1��v�He%��T���*;�|����?��o����B��ٴi���.�/��r隭�����l�[��1����u��^�)��{$�	}M���s���(!�B!�229k���M�R,=�Ь +�p��;4���v��(o(�C��� �~��ޡ@���b��B!�A�W�^���~����NS]#y�#�;��x�����ɞa�i]�"�3����s,��=�0N�}'N;b.^��b,B�`���P�ǉc�1��)����@f�=hw��0����/Rv�Y�zGG��<��� �B�������ߎ�����?�9���<��`��U��N+���1�s?1�O�Q`���O��[(XB!�B!#�/���ѐlOy���(�L۝	��c	2�C��K!�n����)y����B!�E���p����O~�1c�x�#�zl����l�v?�v�3��Vy�:!w��1�M��Ġ�3�~t6��Yuxu=CB�`���]�ǩ���ۯj`40�/�-��@rQ�18n�n�G_~�v��ٍ�mذ����� B!������ޒ�ܯ��:,^�X�heE�Ү{A�2ڷ�m�VYZ��*kX���%�J!ZE"�߅����N��B!�B)|nz�5"Taɞa��K��S�	?0�G1V��v��(�ǯs��J���!!�R���U�V������~�3�x�Ҹ��v���� ��y���@zfA��+����ZL��tn��%�.���i�N��{9�3!z0�N�T���Ξډ��1�`R�2�V0cIݝ�'�ţ�n�C\*'�*�c��0��n�w�}!�BJѦ��?�7n�~�L�:�VQ��w�ڭ��H�R��c�[�@yU�j��R?����H�W������w�!wB!�B!��9~J����t��v�0q;��ݩp�<^.�v/{�����^�u�]x��08H݈B)5�����W^y%��?�555յ�������m�z4�&<�t�=f0�]!w5�׃�XƸt�Dpxd�;�l9Ȑ;!Zp'�fB������쒚��۳TF!��U�p�|�PH��\*;)���-[����MB!���<�6oތ믿��~��*�I�^��U� {�����{��V=25����t��t���M�} k�&�%<B!�B!��'GO
b��.�|~�`���=�GLy�����z�a>�v�~��v�ns�X�uz��BHy �����c�����/~��;.o�P�^�л�����Tz�Z�Pr���Y�f׊�q�pnl�&�BC+C�(a��	��=/�ۏp{k�(�jo׈U����L�=d/�p{�)+��YѺ�d�����B!�������_�_|1����a��ўlb�����ؔ��!X�"���K�,��|n����-����)ڱz�0���#�B!�BHi2�� >�߃��Xf)����u}À�?�y��k~���a4�#�<�;�}}} �BHy�u�V\{�������/�\��s�#�;֋���6������ܕ�+0��2Wl>à{bc�0r?.�c�cOg�!D�wBl�º(z�&��m�!��v�@�h�t�=!J��KZ��/ܮ�Z��p{1D'�)��޽{�����úu�L�O�B)m�P�裏J�K7�p�=�Xך���`W ފ`U�ԃZ�.ٲ�2ȏ5��1����c�=�8oj+��B�z!�B!�R6L�ǿW��`tȴ��7�C�e��_��v'|�R���;w�č7ވ��z�B)?z{{q��cӦM�����ӧ�j���sٷ�<C�}M�r�=���	�+=@Ց
�0�3Ln�D�8a�r�gBdp'�&.��(iۋPEe�H���Su�=�6��?��n��+gE��"Pɷ_y��z�hjj!�BF|����i��ˤk;7��s�׭m^�r")\	V�XJ�J$Ī���CX8;�e�U�K�B!�B!��W�ǉcZ0�Q5��b�����@@�˟Q�e9ܮ�GZ���av��^xA*���� !�B�����k�a۶m�����|Eu���G�]�gh�g����)� 2������}5������	�x��?"��;!6��#��5!2hn�,�&��ͦT�T��S��m_�m̥K����CUU!�2��
�/�}�ᇒhu��{��!��d�Vʂ���k:�} e+��`e(Z%�*e+CO�A\0o�o�1|O!�B!���S��+S:��ݗ�+4�Xf��z,�����b,˾�N�]��nw��#�n���Ӄ;��V�B8!�BFį~�+�������kQ[[k�G�]��gh��U�0>(y�6c�/��_,�1L?~��D�g�����X�{4g&#�	)��N��P#�������4��$R�X��kU>b�����V���!�BF.����G}$M?x�I'���`��U�UM��wu�ݬCA��p{j9�����ƹus�t�$�B!�BJ��χf�!�ѥjnW.b��7(�c��n/�?0�p�֭Rk���Q��!�2�~Ճ>�M�6�n��������J��ݾ��g����
�����[1�2,e�=�����pW'Q��*��>2Ra����?9����T�Qs��􂁌����`6�`��ۋ-P9-H)o�RѺ�?�	��� �B�ڵ?��q�%������4��ӢT.�C�2z�vVv��3�\���к�p%?GE�=��mo��Ś�!B!�B!��X8o=�͉p�N)������>���J��K�`1��B�z�'p�M7���B!җޮ��\w�u��׿��t���	�d7�f��v��)=CO��r7�˖��9�y���ә��� ����z��ȅwB�dƸ ���Ɛ�o:���(�����go`�;ܮ�(�v�����-�c�����?�O>�$!�B����'�����_��f�rE�2ڷ�m�llp"�n$,%��n%��J�2���E)^�~��*�Ww�������}QB!�B!�48�}�{PQQ�[�U�e�g��{�4����#�nw𽥥��z+�z�)B!�����J_~۲e~�ӟb	���v�Av��x�3T�+�%���B��f��,�/Ly������8�nVs�g2Ba���<8�ڏ��6c``H��]!PemoO�SE��U�����^�r�WL'����~�!!�B�X�n���j)�~�i��E�b��!w-�s
����6�~���T��ah^t�i�*D"�݁����e�B!�B�6_��P[#B�
��v�G����,��r�;���+��o��&n��F�޽�B!z<��3���ǯ~�+|�S�*�g脟�g�\�#�n��kו	��jhm�]{\�_��1��g���]��ȃwBr�*�Ws�����%�t*K��z!����Y��R����*�"C4��oVvww�B!�
��Iܿ��o��k���/K!Ȟ�6χ��q�t�=��{RtҊU�N�5�rQ����#���š�S�����B!�B�W��� �:��bU�x��Y�����Y1VΥX�۶�ʱCCCx�Gp�m�a`` �B!f������}|����e�]��{��f�uz���,���u3`��]}ݧ�eQ�<"������!�~��}\�	�O����r'#�	Ɂ�/����<��FPO��k`HTV���{6���v
T��zzz��=�P�vBH�"^c���v�z-> CA����GͨZi���ae~�AFq�x�H���h���G�]��{/�mۆn�ӧO/�(et�B��-X�r����Ě�n�ߖjE+�k<�K?�X3=�B�����{Éc[���$t��B!�B!���	AL�	_0`\���;�bɋ�g����c����ۋ����oGG�T��z�jB!�X����ӟ��Ѐ���7n\^�v�˞��s�_^!�gV��L���tP=��R�d�5~��F�YC��3~�r'#�	Ɂ����ڒnW�܍��u�uE*���I{�R�A��bTV���Ԅ���wظq#!��xݭ��AeUe|��^�+*+��V�ە����4���� B����_�gE�D�����'9,��M۶c��G*5�+_W����2�����M4I��F㷓�`��il@�9�9Ab���!��o���}�{R���'��(��y��=�b����ۭ�U�ǣZ��R������l�F�����W���=��^E!�B!�x���8�b/�P{���vc�PY�����e�0�R�R�;��3��e������ZX	!凔�P̰!f���X��t��\�3���@3jg�w0*�@�L��4kphC��%~[�
�c���I�9b�eBʋU�V��?����㎳��e_;<C��s�wt:�nt�1��b����)g���U>�|��qi�Qc�[�~����0���ȀwB,r�<?z[vJ�G�p{����:��n��2��:�
�C���^x�������B�7a��j��֢�v������&L�~VƷUUWI�fdF��r��xL`��	����"�p{�>~K�S�:�Gs�����c�QuR轿��}}菠��}�۽�=���	K?	!�k�.\����kp�WH׊^�̶�-X���+䞥�A{=�K݂�҂�,N��*�sd܇R�J��ub��*<�!�B!�B��j?Nӌ���~1��K�g�W���٬ˬ�����l��W,˗/��7�,��B��xm�Q��,Œ���vQ��L���m��6_vlo�G��nD�]�`� ��s0����0+"|¾~�,K�?E"�m�	�6"����@�,X�q�V
��ٶR�[E}�S�?R�v3�0t��(^�O�Њg����8)p'�'�b��!-P�U�Z���T�`ZA����z�
&�%��X%�eQ�����s�=X�t���hBH����ѣ1f�Ԍ!�T�֢������ޝmm��ݎ�8�8s.�����:���`�O��=c��q�`{F>�����3��}��Ĩ�@uu��(w�)���8F_o���{z��FO8�t���>��L�Z3:-��%[�lI�|sB�$�����'Ɇc @��l`CH�$˙d�KHv��`ccl�C�-[�uߧ�?�=�]]]=�#�)�ߏ��S]]]����zߧ��BgG�QM�ID|`A�Gy�\17������ډ�@=Ҳd�b�kZ��*־��0��f��^�?1Xe	�u����
7��{�⼅���n�AAAD*��Θ݉ޮ>�Q����)V�)t�,nW��r1_8�����Ʋ���?�0�{�9�z�h�M����'`x`Eӧcڌ�F��B ������Y�	�75cn�<�lp���^�Q��'�E�9ϴA����Nlذ�!���P��Q�0�<��^���]���E���w�%��g�0��Ӄs�s�B]Fu�:� &$p'�(,-���Y*���W)pe���
FPq�1 %���a�^&��
J%3� USS�q���o� ����/S�OCaQah*��:u�1��v�gYu�'ڳ��܉Y���򱺶k�B����]�D��O*W�Tu�n��v�Ƶ�jY(*��T:{�n�8�í�9�ww���ۘ�ԝm��n_�}�+�����z�_�˖-�{�IU7��7&��OGu��=����Y�*�# �@��Víu8���5�� � � � ��������{��#Mf�0�0�
:\�#���<��+���s����&2��k�.�u�]غu+�H�z:E�#M-
�M1{�����MF�q"���s�g�TL������=l����'�:2L�j�H4�~���Ǟ={p�m����*�B�X��Ĝ��>Rΐ����!�tqgm�?C,�0���?{�y��|!��;Z���xi	܉�	�	"�Xlݔgy�<��r�*�pmz8/d�w� �,nw�08���hq{�T~�W[�l�w��]�߿SB��L%��>�N�j�3#�1��m����x��|�#�'��������y���yv]E�#���hi5&��J�� ����'�vĀ���v�~���툡}�q.u�e�mس�Cu��]�]����YZ�M�fL��0�-6�!sy�7��P���)�"��y��˶/���Lض��+U��T�֤�z��}oll�5�\cA�v�ZG�$��D,K�z��܍��A����Z���;X%׳�S�IX��b��jlmAAAA����-�F,��a�#?�qo�M��s{,�X���&`)��1V����)?�'w��?��0�jkkA�]ۘ}���(�65,d��E"9�� v�٤b���0�b�wf���م���Щ�S�DeӦM���G�|��8�Ӓ*d�2��X�%K�I�B�џչ�pNWN�/�G�m�����?���^����-1q!�;Ax��v�Z܆���q/�Reyܹ�=zpJ��Bv98E���.c�o�[�������x�G�����|�L�ʾC��w��f�&�M�Z��=UwC웛���3�iƌ�z���Q�k
Zp�]$�vsŎ�6#xR\Z�lג�;�o��ڝ�P�d��<�v�cWu��B����5��]��"a#v��,s���\vp���cdt��������n��H��R��g�<������d�lh�T>\����[F"���y��nP_��׌{��:1�gY&�"����J�����>��k;28�9�U�9Ȧ�!��>����n
XAAAD���� F[����>�"v����y�9COs,1o����Oq{"���<��>��Sx��ǍXR&c��S*H�)X*Mr�w��G�� '���5�4�2��S,�Qn�#&�#̭�Ә�
s"���0ͶR@g{�v�Iɶٵ���C��	�Fax��9�s�X����=n��L`fY��YOf3��Il�8��,�|�wફ�W^i�W��3�3��,�����I�.�
�����v{9��y���G���k�a�7�^��ʫ�N#��ALLH�N
؏��UC�m�����s�-r�;��r�N��385���P1�࣏>�'�|2%hD���U�%31-,dg���mX�x����%]|c^�t������vE�B�csm�.�R}�I�\�v��_0�7 �ӽ���>y��]��ڎ��Z����o {���t�4��Gttvt������>l������x�	c$�o�%%%)sb�� >�+"wi���o�%|�F�'4����r=�r�����������L��ȝ � � � ��� ��j�)?�0�r�y�0`Or�19�;F|����D�c]��Յ�������;L�Y;������"��`�4��G�K)=���PR63fcFq1��^�%�=t�	�S�PP��3�W-�Iɶ���q��s+�d��u(�7���bn��mm�H�̬�e%�+��y~O0�̙2a��z��� uuu���PTT4n����D���5-��?[b��D��ײ�z,�Y�ݭ�3�#�DAw�PpA�������؜��Ђ^�Fs`�<�S���� U��R��Ǻ�СC���	�P���o�Kf�����Be��{��'���jk��bjM]�ol��k�[d��k�bM/q{�]�5��:�-/�^�i���E�\��ܖ] ��2�G�T��*{�^跌��W�T[�����r��-�hi>�CM�)u '�t��#��ۇ���cٲe	��uY:����͠�5����D�r�E����wk>��n��9��So�������]�AAAAĉ�),6bd8�!f��7t;��e����۳�|����#��eR�L��`�e������;�i�&�`v3f�4�졉�
��P�{o�D�D�a�SS�O3���F��vwv�����	ߓ1"4Ad2����iܛ���(g8�u8E��?�W.r��Et��F��2K�6��4���!��9Mh/���>2�"&$p'��0�R�����:�G^P�`��󲸝�s2Yܞ��۷cÆ���A�	�3��Y������9��Zᠹ��{�\۝�jaA����Ĺ�;�����]۝�v�k�)$�kٕ����+�O܎���k���hn�r.��hj�1-XXc������͇��Ԍ��0�Bg�H'���7���r�-8�3"o�rT��,�V��y��~��Z�^�#�<��W�JX�2+��T!z�����C�=��tM>^�Mw� � � �HyAങm���4ƒ��y(�۝BvQ��-j��S,����[�kN/��n����o��;���� �MaQ��C���3Jf:�������UF�3���C�����H"R���lٲ_��׌�ᩧ����a�e)g���M�s-	����,��T��l�9C!�444�O���o�O�=DL H�Nk��۱���w2�T�۽��5����I�nϧ>�����xTlH�{��b� &3�:�Q%����M�"�`܀K�񤺶Q�]��{��r���%nWu�[^���M�i���������暳̽��ޫ�]&���u<�]-++Ms�b�Y���M��`�7���ALV:::�`ss���+�{�x�=`e<X�kµ���Q$G��y���]8f�pq�Ԧ#���C�`��-�pFu5^�K�^AAAD<a���W����!nF��b�@��m��@0�1V &S,�9�w���3!?mi�������}� 3�X\Z��ٳ03�ʜڳs�A�B�s����a�nAkhb�A�W� �C������W_�/|����3��,�y�t���푞�Q�a��W��K��ς9/׭bĜ!o�O���:qAe>��C���ā��bZ �G��H�%��]5A������r�eׅ�C
�Yܞ� ��?��{��"&%,�T:{6J�f[�(M!�v~�Q�Rܮ��we�jܵ��\ۙ[w�I��n5/��p�R��C�c�O�vCt.��vy;^�|Yܮ��Q9����\�y��]�pIhZ�ب��ى��8x� �����L��9~�a4���k�����IX1����K��]��DsdP�sF
XY'ɕ������X���ű�5�{#Y2AAAD����im�tn�:�s�����3�&pW�b�yC�cw�p"���������������1�	f���-S�ٳȝ�H:�ww��9��`����:�d8�3�;��d���=���ߏo�����O��a�6Ɠ[L���|�ոG<F8�Μ!ˢM�����y+��� �		�	"DaN�+:���Q��#�T�<H%����/A*y�A!h%��?n��v��.n����<�_��W ���f�a��}��2)�)�زf;�k�umR�,h�צ񺶻���������e�T@�ڮ��?��:s�8�ݧ�Eum��O�v�k�k���'vV�<�N���ӧc��%FQOw7��1�{K�!�d�����׿���q��c�ܹ�@��%ӱ!=D�Z���{l��]���|����M;`�Kx����01w6��ˇ��2����&AAAA��ӫ�l݃��W�З�]toL����Y�ܡ������a��!q{�m455a���x��A�v�*-��Yef�pz�G� ����r�lZS����f�55�dlHL6�}�Y�fݺu(--�؜��z�[_���u�6	���f����eR��Fݱ��i���X���"�!�;1�aOX���Co[�Z�*FR�������T��ݿ��ʅ��w7�4e��
DeJ𪹹w�y'��׿� &:�S�P~��tV)��k�
YܮKK�VU�v�[!G�\���Q��a��mJ�E�ф�*!���<�i7��.��Usbvmw��%<�[�ԩXĦeK��{[��1��Cc�~]�u��J���z�~��[oŲe���m�o�x�#��ݸJ�j��*X���z7wY�΍�y�	�@U��d,���!�ݖ�����AAAA��e�A�u�"̎*n�ruX�vٹ=K�ǖ7�l�%���q��"n�G��߱c�!���AL�u���g�)S�bDf��Y6J9���\n9��߈�����C�BbR��k����ظq#�,Y��9C���>{k��%�U|�g�?�3��(n��C3����6��ۆ�-?Ӵ޽X4sv����DfCwb�s~����C��풘ݽ,,l8�ݢ�,O�����\��LM$q{�쑖�ڵ���W�����C��T/Y�9��hjQ�ڈ�k��[X�,�v��.��Hb�q��]�V��M���8\�M!�%׷�E=�]�8��;�������bgE�sAگpG�,s��1��N<h>xuu�ݽ�� ��FCC�����[n��g�9�U�e�,r���D�R��92DO��nl�2^��Bw��*���M���8g^>���3G� � � ����)YX܏=�S�)���{�3��g�6�r	�yC���63!q{�˘(lÆhooALd
�LAY�C�ΦS,��TD�����tک8�Ԅ�����1Qٽ{7���:�p����>��9C��'r�Ж[����q�Q���P��l-�r����:�{c�X�} �eh�;��TH�NLjN��P�oq{80)Pe��;�����p_P�0�^��@9P�Qd���,{��׍�)@EL4rrs1{n���bny��TzE͂��Esmw
�!�U����xK��Z;�k;�`��O�./����-�wtS�,�v�~�H�k�(&W�_���ݵ]�ɵ�т���x���4E_���<TU/M�8��G[�a4�գv�^���� &
�����{��e�]f�c2��#QcY'^"w�9�M��V�ۓ�ً9��)n��y�*<���ۋ4��ƹ5��nAAA١?�O�Չ��G�0E�.`��Àe�������b���y���2"��)'���`�z,���s��_��_08H)�ă��O�6'-[b�~	b2�����U������4��lj=�QgC�HGG�!r��w��K.�ĥ1�w��O��K���s�G6���{k��?ԅ�!,)�����l��3fwㅺ��1�������,�D�@=4/a{�@U �`��K���[�.�g�F�Jp\��VV�څ!Q���(n� 1Q�RT�y��7>���R��[M�\�5$͵])$��!nK�����'�N��brm���
��p8�z���>j�5��?��]ؚR����cum�����\:{�1{��ho���z��p7�6� 2���a<�����;Z���%T��Ht i,������k���<�U���)Xe��%G�p�<������j��G����h�A� � � ��˧�G���a�ۃ1��Y~P�Ypo�k�%���ڕ�X^#?G��SN0��,_��� �<�b"���U6s�S~A>�v�!q;A��:}�1-Y������C���݇��A�3������~|�[�2�s���F����c��?{߿"l�%�c����?u�0�н����)�Kd�Ed($p'&%E�YX3�	Cp�ڃ�80X�����`���^�A��9V�omtq��d�G�ǞN{����SO� 2�¢B#5��ųJ�r[��丶C!n]��]˔}�uy��?V���b|
ۍ?_����G ���~Im� �0.�v�X�k��,�k���横�u�;����j��>i�:�eF�cZu����`_]v�܅�#��D���kmm5ݧO����X���^�ږ-r_����=9X���,h���#ݟ�e�m=h��EΡc�JP9���$r'� � � �h|rA�-���*a{4q{0 ��v>Q�3s�ޣ?˂v�(K�b��+n��l�v?����ꫯ� &y�y�;�a�U2{�k�I� �0w����tdt���ذ����& �_KKn��1�#-�$���XE��,nמ7���/�e�%���=gȄ��������QD�Awb����]ރގ�1�����T�H���,�}AZ��ۅ!ҏo�瓵~2����O&����Ad*�)r�bC�M��Xf
xn�.|����н��pmR��.��ua�HZ.w��!��ro'v�P�]}<��L�k���p=ͪ���Q������%�:ˋta=sU�Q��Wy�uW?U뱾O)���+W����kOcC�|��{k1:J��ǟ��'477���FEEEF�)r�X%���Э�2V��TA+�����n���&v�PY�����S|�e���c�4���]���AAAAx��,�����|a���XcS,o����yC��a���bv�}��.ng# �[�۶mAd2��3o�a�5{���8�
�V�ߧ��ߊ�v�������� �L��:�6`����3�:�j�6������϶���t��v|��ãAv�aiI5v��DfAwb�q�B=--�����Ә���<wY�)@�r_�DA�Ӆ��8���Bܞ� �I[�~=6m���4���	�+��[��Z�'��v��]%��E��>�;�h��p��.�)�s;��Ph\��*�v���X�ǵݽY��{?uE���mW�4Kq�I����5��4g=(]��m��fwGjk��ݵ_�J��>��jj�v?}���E͢E�480���Z|�m���N�K�]s�5��}ɒ%��g�Q~�%#x�G�.���e汓]ܳ�C�����*��'/�Z�T��}���*�ŋ�S0��]'� � � ����� *�F	�an�	�CY��*W��f��M��X��!뵙/t����D2A�>��`�z,fv��"w��D�b^U���>��A��;sV�1�>��nAc�>��v���� 2�͛7�;����.,]�4�9C?m���]Ŀ�=��0���ʣ?k�|a�џ�W�9V�������j#�����X�݈�eh�;��H�NL*>Z���ûMq{����)@�}A��n�?�p�h�vU��{��;w�4>{����-���A)��la�7��ڮ�%nwmZ�����M�D��C!�v���%$W���Mu���]d�]�U����bn�wm/ѥ2�E���͸����4���|]��b��T��#�]l+7?K�/3���>���aǖmhnjAd�~���&6n܈�N:)��u���-r�
j�E��u����B���)�ٞW��ay�J��6|M�UO{έ)�ov� � � � �� pjq�z�=s�^��\��;4��bsn��s��2u�0��t��*����q�w���ĉDf��UL�^Y����<�onI�{Ǧ�����6c�}���QAd
,gx��Wǜ3d��`},��K�.�����o�?[�>k�Gfx��l9�C0Â�<!�
���ϟ�Յ
1Bw"C �;1iX83�i�{�%�������C@p_���GT���C2b	R�%($����X�mݺ��r�m�HxP�9�3���h�)��\�3�\ە��Q��x��C�'[�m�K�k�K��,�v�$��C�����n.-(���+VS{{;�|�;�mGWg'"�imm���_o��]�6�n~�e��ݹ=y��!9�_u��U��������v+`�R�S*j�AAAar~�0zۺ��v��ݕG�	�R�P=�stc�,���*�x�c%#�7���/����Z��ߏ��<D�îs����s�8rA��3���9�nj6���cxx���^�o���K|�l��d�/����{�g���U��6ms,����'�ź�\!�z��p~u>^� Ad$p'&�9Y8*�4Y J�<ە�(�Ђf`�����Q�`U�;0�zn�%m�{���-(�����Ђ �t�}�K�f��f�+*��L4��]����#\��+;�ʞ�v��
1��>;���>(���z���+8廉��&�jA�?�v�v�;��G껣�(_v>�y<� ����}0�������u.������]'Jߥ���˻z7��ǟt"�;��:���w`�@�Joo/֯_o<�q�e�������XJ�<{�;.s^E���M��W�";���(#@e;h��G�{�f�աrz%�;FAAAA���k���r 9��Qs�*��@8wP���X~M�����C4c�v��)��&Q9��l#��D���4�x�	<��#�<A�3�PV>�q{ @"4�HW�o�9e�4r��ۏ��z45��J��=������6r��A��3�I��ݙ/4J�yD�8������N��r����=���tD5���[������������Ĥ`mE?z��L���k�A1Xe/p/�Z0�
Hy��;�ܮ����|JEP��:�c��K/�� E�)�S���T��j��
F3�º�D��b]�Brg�\��^[%�p
�]�AW
�=��Z�v]�w�k;��O/q��OBr��v�L�hS)܆[����.��E��s�\���v}�V�&���/������2���vg����?q%��Q��z�a�Y����}����� ҍ���>�������m��fZ�*m�E�Z��Sts���5� "���*�"i�xpJ
PAz/���"`548����g&(^EAAALbV��{]#=��Jq��;:r������vA����ܡ��$k>�ǫ���z�!<�� �tf괩���6��|a� 2vO0A�1���������Bb�HGX���DSS���jCW��9����D�>g��X*���Q���P��jΛ���rS�.��8	&YY]�XZ� ;SҐHoH�NLx��d���	���� �/q{@b09@ɅAv\��VV����L�.�t	>����z~�ӟ��G��(�S����WV`��j̜Uj��S����n\�a�9�k���n��K�n����#�g�;wS��/C)��ݵ].��)���x���tm� ̏�w��;�k���¾)>����?_׹��O���Oe�5�����v�ל����U6�KJp��?�Ύ��`;>غ�== �t�g�A__n��c8�LX�m�$B�n��o��!W�JzPu�|u�2��O�X���Ἢix~7�� � � ��Ɍ�,,�:��`��J"�H�v{�g��=�1V$�v��nq��SHD�/Q��T��\I��>���7"������
TV/��Ad>��X�t	�Ο�C���{j���"�x����ڊu��aʔ)�y2F2\�Ǜ'�wn�k��̈́EJc,�G���q_�#?��23g�p�a�;/NG#=[�B���h̝��A݈H_(�MLhV�Ά־���AQ�.�\�)G�J�#/�e�|�����@�xF"��J�:��B6� ^� ҉¢B�*+��WA*�x�]��f<*q���) �����ׇ�k�R��
���߮F#��K�g���)X���FT��p	�!��"�ve]��]*�$lw��r��U�N!���x\�UsN%�Uյ¹#tTފ�37��ӵ]:?<��l_��A�i�g��SN��9	���a��7��;�V��W�BOOn��6et�*��r��YƯQ�u����C���#92�a��`�����Lv��.��ҝ�v����gTW�ս�0(AAA1���N?��=]C�e�>+r���k{0<�37�
�D�\��K%h]�Ŝ�#�0���d��Zv��a�_����@�Ƭ9eX�����!�۳1!�RX����}՚��߰u���pS3"����~gc�{�3f�4�7�u��E+r7s�,_h��f=��?��k!	ݝ�A�K*��/�?����}xn7�C�/$p'&,��C#��vPJ�<��f���v��rap
�Š<�qo�ma�q�_�1���u�S�������/� ����[1Ջ�pjz��q�?��nV�!��k�Y7��Nնk]U�L�_��J�,���r�NY�C®�vH墛�&W��ס�U]�{;Ϊ�|Wg����!��?wW=�a����sQ�����z�黠]�� <���Gw�qm�ͅ�	�+�0��2t=�m`��� A��W_}�8�����dt�*��,�m󺠇����<J�`��t�2��w���b��U,XfMB���w�bYi5�Ӱ�AAA�$��ݭ��	c}��d���s�����?�"l�h�%�Y��i2�����x�8p 7�|3�n�
�HX,oμr̫����� br�tGl�61�@��=�ݵC�� �t��^õ�^�{�eee���1���*�mE���l,���������򽬘/G~�-�r�QF���\���zkk���rq'��ÁaN7���� �jxA��/�T��])l�>��%hU� ��r�e�It�*Ձ�X�a����/��2"�L)*D��E���Fn^�Q���k��7����}�����Xׯ���:����06�vsYl���Ϳ�-�>��t�]�U�Nq�s\�U�w�p���q�k8ޮ��j�YO�w|����[y|�z��X쥭U=� ձ�%���*��w�S���vT}�M���?�{҉�W[���mAݞ� �T��o��o�ƍ1w�ܔ��E�!x��d���,|��$w-�������]�y��+8�%rwM�;��l6��,t��	� � � b�qlyC-{|�U9�@ `���GV��,c�5Ų̱��!���D��D2-��ZV[[��n�	�v�A�3fc������Bwg�i�AĤ���:�h�X�
�5b��8t�	�j6o�l��+++Ǖ��[/Y"w�D���2�u0�^.�zޝ3�.��{��{�-��<�V��s���A2�"�����#90��T�/$q{�����~�t���v��=U"�T�bY����peOD*)+��E˖a��2�rݧ`]7+������;છ@�vQ ,���b��sA��(�D�b}I��Aֱ
k�>~���T`k�������w;~��ȵ=r߅�9�>G��R�n�9�]�-U5ա�---x��M���mA��M�6��3VUUU)�'*x5^�
���(q.�.�n���Y�tqĠ�3@��9t��+)X580�O�����|+�FAAA��)����E��=j�P4�
�"vU�p���Ǳ���.��t��ر��744� RI0;��U�Y��fLA�����ü�
cjomÞ������#$4%R����q�5���{�ŢE�&��=тw�����}=wq�yC������_{�gu�P��a�)�/�G��`AZ��ɝH/H�NL8�/��P�n����y��tl��UkR�kxA�{����u�ReZ *��>�[o�o��6"�?6���\�b9�N���c� B��}��Q]�b��B��|sQ�Z���[��^sl��j�����;�:ŅΉsmw���G�;����]W�K�k�]�9��^:��}u�߬6V�vm�}�W��Jq����wն�����8�3p��>�w����|=�� �d��,`�D�K�.��"���'�6:��.�7w��IRq�����΃V^�`P=� u=~��ނ��U�ov� �� L����n�<����t����-|�����=����Q:����!���>�ͻ� � ��?�O+mG_���;������v���+�)�h�%������#1Qr��e���[nAss3"UL),D��X��u� �/l���N>��;�{���m;���	"ٰqX�����ի'��=��]d<"ws���P��,c�M�<F~�9Ax�ew1_(
އ��p��.�X7�d�E�$p'&s��3T?f�q!���C��CR�:��;h�z�Y�-tO|`i,��td�߿�֭�֭[A�&� Ջ�f�"���zֳn`�����f��7�����}���n������rmג��W�5�~&ҵ�YW5����;�ێ�0_�^O�c�x��;���� ��d|7�Bv�>z�]�^�w���ꃺ���C���T�q<��煮/��9��>
{w��;}�(C$���:#`u��wc͚5i%rIa���?��wV�ְ@zP����yQ�.��T~�Vb���nۋ5sb;HAd8L����_�I�+��\{ɩ�^��[~�rҷ=uJ^h�y�Ȱ�{��/���¦]� � &7��9������*�r�jq����1�����ͱ��He~1����o��a��F&�T����-���J��AD�d�dc��%�M��k�N:��H6���V��Nr��&�V�8E�F�s���;߮<�2Ĳs��s��\�"g��=m8�����HH�NL�C��S����sdLjq�-f��T.1{�v�z�=V��OA{�Y�w���7ߌ={�� �Iq�Lí}���)Sh�f�����)6�E��b��B��|���qvm7���S�\ەhH�k���ǎ��졦,soGCl��
��b.~��vU�s��~s��zv5]:���y�]^/��[�v�O"uq��.�=Q��Q��o,\��B���Flz�]�ڹ�,���p�u�)V���K K-r���]l���vq�2DzP��u�I�r�<��+�F4̡a	Lx9<2�ށ!&��9����	A������'.Kq;����C=����"�L-�ų���"��` sgNE:��݇��A�!/'�iS��G��>AaN�������A)o��/��@x�g��=�O�9Cٽ��ˇ{�ʵ����a���Y��#֯_���>D2a���h�R�,-AD<a�s�SG[�!t�W[o��	"Y��������ߎ3�<�̰b�h�e�+󅬢`����s��M�n��,�'��z�4!��o�����0�W}�����r���vu�*�s�g���i��L��S2��~�!n��444� �EɬR,]�e�ч8�Dn>�9����]ۥz��Vs�e��D�������$�b�Lخ��T~u�^<\�]
k��Bl� �%����>v��x���oG�?�vu=W��ǵ]� ƶ7�����8A��r�7�r�q��8?T�tn�rm׌o�e�,a���}��3�s>�WŻ＃�����QD����7��N�+C"E�"�Xi�F���ӭd���]re�T�,��;�;�+X���*.v���a���"����|����՟Ƽ�i����v��?���^~ã�/q������p�E�`IE�Q�x��<�[����{�������5�t����o|uM� �xS������4��휛��	��߂��u;��3QE�9�<~��q�q��4�t�[��k|�	di��O��`���������{� �T��x���9�s{0,j��oc�H��	�`����^��Tc%#/q�K/����CC�02�<؃35K��y�{�$� ҃���8���`嚣�k���ڍ�!�ɡ�����s�!3,�nc,Y�6�
���ݾ���<�w>Qe�e9��^K0�hv�&�H=$p'&ǖ�߲'������#�b^0"v�tj���ܹ���۷�h�w�	ڗ��pn��8n�=�����˵=\S^ٱ~b\���IqmWvJø]��n��v�f	��#���\۝N����w<��=|�|����vݟ�|.H;��|U�u���\�}w(�.�Aq��e��d��������q~���יQ<��uN<�d���&��λ��!X�[�w�qǸ]�p�I]��(�u���T�\ /���W/w��O��U�+COG+�V����{���|�/W:���@��=w}�l\u�q��~���܏�E�����Ū�2Gyy�4<}�e�����g^݄tᴣk��-�ή����<�t�U���'Q{�/����۾��WT"a����ع�0v�o&��=����x�p�'�������G��g���*���ጣq��V��_���W5��	�0a�>�PԊ�^&Bu;�g�$n
�v/��(�l���!�R��X�t�G�;�����^0��### �d���ՋaѲ%���AD��/��QǮ1t�{�b������h�a����/L+��H����m��Y2S$c���.���o�g�Y'��<� �2�/�a�����~/����)���Ǒ��}�����=z���|��k����#���T���|�o������"��]�����������:�ͩ�����y�+�ӥ:�C,+�U�g%��/�Z��k�����v�R}��^�vYoK�Ocpm����x	Wv�[���?q;�z�sm��bu>פ��E��y���4i�]�����:b7���pHW�]�V��H:�cqm�z@zo��E9&��w-�]),,�)�~Ǟp�mق���-z�H(�����l䀳�>;�E���r������ŝ��_m'w�#C@�Ƞ[.�^w�ɝ;2�ߏ��a����L�/�����ϒ�]dѼ�������x���b�s�'��_?��x���q�v�6����kj��͗b�te�̩�9t��?Ǉ�� �.�b��8n�<d2��9x캋q΍���~��D������D�/�u%>s�hh� ?J�O�S�.�ы�#K2��mW���W��w�A��_=���N��Q�}:�[�C������"ve���m��HA{<s����Ƴ�>�x�F�$��.\�Ջ"+�FM#br��k.]b<t���;�lCwW"�0��~��ƽ�E]��o�C�0Q�_���Bwݺ�����W1O��G�/�&p�Ŝax����[3���H)��"0��i����9�vo��� �ۃ.q{��r�da�+P�)l7zQ�H���x�O"�dmٲ��777� s`�Y�KV,Gn^���L���^���ZU"�����z*Q�؀ ��pmw����4Kծ�
'x=�X^(W�5��:��a������[E�K
!�s��um��w�&��u>w�s}򹠉���k?� �U-Z�P����wm��>o]�����q4���+y�k�q'��k�`�����EoO"���l�ڵ%r�$xO,���H.�r���ێ����`���Sl��t�.�la� �rg�{���Ŋ���!��0Q���L
���Y�)n��/֦Z�~�1�>���vά�xq㕸�'I�N�&X����ql���9˫f�o���=�"�Đ�"�t�s�'���*�Ǒs���m_@���u�:~�iB�� &='��F_K��7
yC��}�v�˯{��/�G}�̱&^�/��_��x衇H�N$���%X�r9��+OQ�� "2잣�z*Ta}v��m4�"�8��9L��\�/��Ҵ�{�:��QK���Z
��x<ͱc�F�{��BW[^��7�hID�H��AD��� zZ[� U�����]N�R��L^0��X�ڼy3n��&���8~��
?�=Y��=RE*�Ͽ+�D��l~uj/6��b����PԶb�ctd4J��TXnQ��ha���O"X�����кYf�˷���@ +����/�Gپ:W����*��έ;֮r&?�qe�dl�튦��pe�3ʎ����!5��.��-�V�s��c�}��������h�Q/�_M<��ύ=�=:��uٵ�ѧ�����st��}�L�;~�v���xpB�3��GFGB��/������y|�4i�'�Q�d�R,Z��v~����d&�o�����u�>�,`u�w��\W��H*K����%����Uve��T�1�e^n�^.�V�:��;�n�= ��!�	"��1���s�-�_|����@"w"v�P�?��,.�D�SW�/���?�"1d��=��&r����=�}�H�>�_:O�r	��� ��Q�g�S���ͱ���ͱ<��nc�(�����)z�I�p݋t�/2X<�'��~��1�A��	ۗ�Za�	� 2v/1��Ҙl����C[K+"�{�|��^q����$:��Dn�)r7J�eJwV?��{��a�w1�(�ٲy��7���d�E����~��������Xbv9@���G�J=���s���r�2cx����z��w�~�z��� //񀋾R%|c�3U�r�l���g7@�ھ����;sV)f�)CNnz���)���#�L�<���)L�PiKU4��H˭m۳�ѹ���$J��zh��t*�u]]nm�7�Gt���׹f�?�v������sn0�p�[��k��
:mvN57���w��6]�Q=M1�t��@cc�}�v��Z�>���j��v�w���]�]��<4ڊ7��ѫ�췣��A���<T>x��$�ϡ��Qt�����Σ���a�w���C~~��7ԇ�o>`�\R�[�ީr�a��{����=�������k�g>�q�"zR-N�׼����o�f~sٱc�Qte�B���:U�3�틎b Jpl�
XqW��ĂV�-qzU�TG��Μq�"<~��2J�αD��;� �2mJ���
�h.&"�|�ll�sИ�Đi"�L�s�1'��I�>>}�r<���d�o<A��@�o��fu��+�Q��	V�%n�#B���Ja�%^�"w��-ng�g+Ѣ�L�/2X��?�)~��g<`��M*He<����~:�RU�/�6���a�̙�����?����m���a��;K�~e���;;12<��޾�l?��>22����m�����[�J�N�}������$� �������v�kH�'���s]P�̩ؾ���T��c����x��=]��ݾh�%�ew)o��_�y����/s�f.P�e�%����!�1����;��,(:Fd$�9YX<��р��EG�H��*W��3@�v`H�z<D�j����2��;:��7��8�Ͽ�/50�z�����qO�O�;��=�D͒�X�b�!d��o�8�۰�݀�|Y�`֜2��)zSiX�:�RD��jn�����d]^5_����&D/S�I՟��A̫�p�Ŷ\}���y}���6��n�Kf�:��ɵݵ?R���0*j�؎�x��[��b��ja]�ٵ�%@W}nBف}�Q8m*�M�f�I����Z�Spc�ك%�,Q�Gҹ��y�Br=j������e�<�7��QM�H!l�I.3��֑����ĩ�lۆ���/F�<Y��]��}�@
�����;φd���.��D�>E�&�`2�ijw�`-oG|��#��:�+_�V<@%�1�)�]��P�F"w�HG�Б	��1S)�6/l�"��	�0q��q���3�����g^���A$�L�g����D�υ��>�����{t"���Oĝ_:�tj#"&�� =�m֨��>G}���b�0(�����\�?�v�������;LF~��rK?�����c�!��8H�rWl?S��#�d�w�}�:˙^\l�SJf�J��y�:'/5F1욗�m�z����ܜIy�#,қ��g��HY)2"Sw��H�hJ�_:�,t�Eu�"��p7:B�J�f����բ$j��o]�`#�����+_���l��э�4��Frq�m�r��]����`0���.	�{�[pւ*�~/��ɇ�DF�v� z��M����0����AZ�.� l�����ʅ����XĽ�؞���7�4�흝� �xR�x!��^���|K������̑���w?2�K�m���y�=����-�b��^� ؽ&�r����B�+mǫ��-nW�ý⮺J���7��ۅG�C$��ˌ}�e�U�ե��9=J=��!��~)>_�9C ��z=�}W
୾kR���P�� ��)nW}w�A���!���p}�=X��#��C�m�yM�X�6���^�+W`������ X@��{�5~�>���&$�$���x��}����bpc��/��]X��Eq��R�1����#8v�a��,��h��A���v����c{=��	o&�s�HU�<�������8����;�»���=���s���ƫp�m$r�C0��{��W�},���Us�1ں�l;o��Aר�YR�0�-lW�`��v3�ǅ�$n��>�C���?��?�x�>����	�X��m?�s6U�O�3X��[Lоb�*���Nڶ����x s�O���l۩�>s�RX���))�~*�}xh}��O����;P8�����T{3ޯ��;?��Ҙ���m5���E*���>k��ֱ�'C��x��G��x��ER��׼h�e;����^Bw�C���rѻ�kR:���A{ ���K��acɅ�D�qFuݭ��ӝ�ク�A�1808VQ�����)��+���T{,A�M�6��[o%q;7�w��r>��gb��eVY,�	�u�"x��J[���:8���C+�ϕ���m�I ,�����*�/oRզB��*��+��
�=l�s�@\W��Z�c��OA#�藏�x�]�k����R��q~hb�z����s�}���Ƈ��k������Ֆ.���<���v���n<5i���Sף�	o����x��;�#�(�R t���c�r�Jl۲y���O��91�`����ϸ7fN�vU�Iu *�~���G�"�����1�n�VG�E7w/76��t��ixiWj��$��yY�G��ف��4E�W��۞$�;�dza��}T͜����p��y�F�+V��*�YT>�6�?y9�|�����z���`^�Z�Lႏ�0��~au��r|����y��A�Ω�k�ܙ�{S�ܽ����Ǯ�g���9A����jЈ�@�!l��ޮ���g�F}��da�Cܮ�ٌ�̱�C����x�b�D�ۉ�Mn^.V�Y�yU ��,̞;ǘlw6���/����_�*���K�n��R��~A6�b.�����B�aV �0�\6�R�#����+s��/�����N$�E� r;k�%
�E�����2H���m�AU��^��j�/�x��A�͛7�n@kk+"̚S����iӧ���ݖ�ݿ���e�zItm�b;
�xF��{��XW�)���U�-��]MK�
vَ��\��\m��ޡ�������.w>w-�����j�N9��z����U���p=���-]%Z�<�����{��%$w�]�ﰲ�C��(?��8?T�)
��ڮE�>z���òU+���w���H�S��ą��ٽ�\�T1z$R#`����i���iJ��j�A���ܙ��� �{�H��E71`�xN���_�zA��	^x�EJ�Ι9���3'��A�EL��E��.������������0~ے�>}�e�Ȋ�q�s�?���w�ǖ=�*���u��[d
O����������9�.N�I��1D�w]��n}�D�
ʊ��ԭ��t�#��Y���>h8T}��l��W�7��\�y�P%l�m�gL(q�L<�eq���G$n'�ʔ�)X�r�#q;A�����yg��~�nڌ��D<`"wvo��/9a"w�T��3��3�}��������n��ϑ��9�5�`�5�߇s*���n�Ƀ�6"c�]��+:��^�rk�
R�V��=R� ��u�[�.��T6*��4�2���֭[q��ד������kV��d�U6�]�òXw7#	��6����>"
����Cخ�OO�v�G�J�v(��k���[�n���{�]S�E��.���<����d����Ӫ�j�1���Oa]���＼|�t��X�z�z��x��M����������kצ��B2�=X��r�5�};��,8$�2�`���۴E�b��^�D���2x
�E'!`5s`f����"U|�����5!��#*0��Kw]e�L7�N'e"uL/�3ܵc}��+�?�?����w`����Zw)>zԂ1�ÄΏ]w1θ�1����{�s럊Y�Μ���+R.r���vN�ܙ����uO�����e����m_@y�T16Ψ���	9�Q�-�`��=�s{Б+�D.q�۽G|�f�%��+��I�_2�*q�O~����?Aă��,;j%�V�׺]{@1�a�%�A���P�{/�oي��~�x���7��ϯ�⊄��3I��c,9_��K��9Ckh#ox�a�%�]9C�,<�۲�V-�kud�E$�ù�:�Z�� UPREpa0�� U�%n����rb��0q)n߾};n��F��h�T�X}��q�}�ĸ�×^�*d���&صݵ}�(W)�7�
!���{
x�y��S���S,��K,=�vc[.���?�O���յ=�~T�v�s
1��<R�����������wK���h��~�.���}1�)��Q�x�ßk;;��_O��y�MZO���0�h*�\�)w�	x��~�1V���p�=���g�yfZ���u���M¿��¯Ztw.xw��Eѻ������� Λ�-w�jpp���๽ "�\���x�;"��!w��ڌT����:��پ��f���~m��K1s���X^5��:�]}�|�/�iW�]���q�ݿ��}��b�t���'��L�����-�ണkb^��W6%���[2߼�C��&r>����'�ߨ��Ǐ�ƿ��9��=� �FŴ r;�Q�-a�Os,y�g�e��˿{;�	q�r��H��=��S�����1^�)�ңVb�E�
��w!��,�{���QQ]��;vb���1<D�ネ���/��҄���
ʓ+Z��͈�X�\�c,ކ���'s��˞Wb9\�]Y9��S��S�p��D�D�!�;��.b�ew��\u�*�C��
#�ۣ;0h^����C:Γ|�&ng��MM��&�{�s�ꕡ?�9n�3���) ���%���WJ��rgOm�K+���Gj4�vQ�X�tnõu.V�g�]��s���vR�ڮ��q�\�5Y �X�5�k��ϱ����{�:���Q�X�� ���8]��:�Ee͋�����3�q����	���?���Ac�9��_���-��'?I"��+�$�j1`�_�C�^�*�2_�XY*���!j�WG���8����`A$�>���gb��t�"���J~���xrݥ�W:��:3�����3'�]��>an�/l��p6�˾C�t���ݘ>�	L�~�]����\jY��U�:���8����&r����йq��"��͝x���0kF��u�/�w^i���o�d�g����v��� M �w�	���ߣY�X�ܵ=�)�רϼ�;wY�M�nbF��=��X� ��E�xꩧ���?��ILl�w����8z5r��2� �h�{��+W�z�B�ܶ�>�a�.�X`���c$[�az$�3�6�r	�a�y;�+���e�.c�.�G�xb������씙�x���8� 	܉�gJ���&�cR��vS�΅�{�,n���1��Q0� JO��]�ߵkn��8@	kbl����eK�?��sW@���S�ڮ��U��.�c���(���mE�;��u�rY.��\H�k�����>j�e�rx;Q]�5�W��<����|���õ]�S�Br���N�{��יl�r_�k�k۪��~���z:7�v�mM<n�`hB�xϘ;>.�WaǶ�x�OBwW7"Vp������~�� R���ɞ���Ќ%cv���@�s�A;h�P^NUx
t֢r�Է�ȝ ��g>���Ӆ1�ߘ`���R/ngl�kƙ�����9|dE����M�ó����p�&��X��-]���'�{�104�+����8��cj�9d_}�)����A�'SD����������_�-e�v�{�c|�M��앳g�^oIE)~u�U���P{&_=�Dl�ҧ|�l�͹5:z[;g�l��=�)V�Q�M1��Q���+_(�Ϳ�U�X��K�y����'q;1n��+����)E��#� Lrrs�꘣����mނ�u ����J>��q�|�%�P�з1��8���ce)^���9� r���]vr�r�R���gWO��{�A"����H{ήF[��
z�Da�������gx�D;0D#�L����L�~�uס���D��"k���/(p-�/lO�k�R���{�`����v�8�7�\�\7�MC�?V�*�v�=�������r]���vm7�";��c��O]Ѧ����'�ZW��D�*�v�8[��v�1V��5���_
�����rm�r����޸��������L�]ۭ�T��{Ͷ���X���,��o��7��W�� b����pr�����'��cB��H񜏴��ί��;�DvPR�6mA���Õ!�ҝ.�`�J���<�㧵a�4�R�� ʅ[�G�sᘜ��E��i��3����y���վ�3D���L����Sgg&~�KS[7.�����s��G�����Oo�<>y��1�qř��__x[�!�XHw�{�:��44w��c\3w����+1db"w�;1`���^y�y�� b|,+b�u����5�s�����]��QG}vc��Y��yD�����yղ^x��?��c��d&V����?0KA�)�:'��QZԄ-߄��vD�����z��^p����t��z�)rg�Ǉ������ +�1�S�.�ܭџ�������a�5�V��3`w�("Q���HkN(�FoK�ہAZ���a�{�R��^0]b!��6��ۇ�n��x%�X�1�kN8ť%�S���<�/���F��õ��u�z�׵�-���k�������k�S�<v�sޖ�<�-��}S|��z��{��K�%ӵ�%�������1�]U�e~��:�P�v�?��%lZ)���j��3�r�ǰ�c����M�����X�n���pL�<�(<��X�k�5�"m�[W��T���=R����]܍���+6�vv`m�4�v�H_8�h<���M�HGq;�	|�������&����|�[�����Q2m�����w`�o���?�:84�������ŧNX������;�$l��+ b#]E���.�x������������^����B�{��?��"w�����v.?s��A�r�0�;W�gyC/S,[�p�����G}VO���W��I�y*��/����^���8����)S��أ1��AD|�5��<�l4���w��@?"���q�=����sN���W4�:Y���smAX�ȷ�����2��]��|��34���B�Φ�ZP�>��*� H�N�-�Y(i�/a�5p�/���'�C�HT?>�;���� �X`�,?zj�,v����k����*��"Xq���W)P�M�.�]��1����f���
a���K�.W��EBre]���SW��)�v�I�Tۚ���~�Ӑ�Õby(����{i����.���������/��5g�z��q�qlT}ڒ���Y�ӵ=�-���En�:nN!��������?sHe�}
����_��)����g��+�Z�W^��6� ���ى�o��pfX�bE܂=�h��v��|�}ݓ��<`��BW���̕!,xծ�a��Y�j��KKj���Fx �x3��"?��7����^w�!��^��i�}�~�Y3
���+Gg��ߥ|�E�_�9���#�����ǿ��9�u��׿�S���Ͽ��J$�J��ܙ���?�3�[�Lܾ��@�q���8ƿ����_�W�6n���'��=1�m�y��p�G�� ��sN��[��������b���AK䞌Q���1�<_:��㙻����+$n'���.\��V�]H�B�(ؽLeM5�++���رu��B��oܸ�����'>�+?���x���c3Ɗ$t7G~s��P�=����B�nc�t����nDB��|"m���>�����T��]���],a{��)nD��ہ!�H��g"�[o�;v� A��}�Vc�Ն����ο�o&�z��,zU���F=����\݀-Z�k��O��X-�w�G!(�ۊ�w��ڽ;TN�\~����vI�5+� 
�ݮ����v�}7߹�Ϣ�PO~����ӵ��٫�ݿk����D�&��#�Q��r��9]�=�7�nWQ��nh�����k����O�;m��ֶ�����:��D��r\��/aۖ-��W�����)< �{��[n1��.\�Dw����@�S����,(v�nP�vrgx�ۙ+���]��� U�`��5�<� j���wFDt���_?o�9|w7ο����KQ1۟ӯ!2]�!r�D��o]tJL�v�??�g��·�4�h_��9������ĥ1�[���sNZ�g^�"v�������W�~�������˱���ҏ�� ���19�?��i��.S{����^�������xn����>���������y���A��5s���9��]�����}��>K�X<W��!�W .�.y����7�����o��"��+���Ea����� ����^���*����qp��_�~�z��OW>0]���cTc,�w��	Bw�����\����N��������qpp���KQD��X���Ob��~&��t{A�[�%ƈhc,1�رDA�F�*R�(W����3�3󴙝�{��7��vg�y�;�3�;��g>��/r��Y4����Gk�z��3�m���D�!�;��;(��[}<����]������#M�x��܌+��o��&���AA����&O@�JU��k{x� m�iT�vYt*��U�f��W�;"DU�tEq�{��vS�S'��t`����)��6<��3Ko���.t�6�v(�T��\��퐘k�鬔�&��YyU��ۿL[�m�m�.l]�\_�x�]�FHȵ��ݳ��,��b���l7�!]�w���~�v����E:~ŵ����د�|��P��CǍÐa���/��7���ƍq��c��0`@�N�����䞏7[�҉�M˝Nuq����w��}o�����c�@D�3{<n��r^�n����;-'�ic���S�%�<��Ex��u r� ��~��^@G�9��w�#��_�btt��$�N"��j����{yp��������^<��ۗ����v6��7�y��l��������xnX�+N�Օ���l��H�.%��p R,�ꆶ9�W�woq��	����#���d�۳I �����ۖ1ց@A�\Qa	����� "3�s�c�ƖM�-�{cC#"���V�����=Ǝ�qy*E��ZNl"w��S7���\���C�k���y'w�џ���&�|��>-��V݁H.$p'��>!�7m l1{�����=| ��*���&���T�td�(=Y��]xW_}5�.]
�BiY�0jj��>����G.�X��ڮ�s�k;08m�fS�ڮ��%��,'k]��-�C̵]��H�Y����/���W���_D�����Z�ݐ&)��!L3M��w\���"��W{l�!�w���&����1y����\��,��]����	����sg���I;n��Ǔ���VD4V�Ze%���{uuu���{'��dw��g�����*���IX	.�19qr߻c#����ɑ� �����<��0��W܏�ߙ�o�41�<�J��𒯑�=�a_u���/l�]h�M�?؆�-X����|���<H�DaN�]~�"�Da��{~s:��0,�y�����<��;?����)������'�=+��gcH�*�f�߇杭�{{W?�����v�{{&F}�T�.Y$3��?����џ��;���>#ǎvrbADfa�i����?���>짛ֈ����㷿�-n��&6,�&S�ɾ�����!�]Ï���|��~"w��.�
�ڠ�fȮ�t��}��avM+]Mrd"��Ed̩pz�.47�(..R����RT�;KL����{�	�ˁ���N�"V��9s]�����3π �0pH�%n/.QݱbumG\�k��?v���ѩ��K+ί���?T���	�u����$mw)�e�q"7]��<�S�rrf)T}[��W����M�>��m�D���
R<�45v�g�sm���ziں�+�,~�v�_��4B�X\�����ƦG��͵]Z��S��Ը�ێ�rLr?�^��.�e�sl�~}���V��.���������zp����ҥK�D��{=���C�+a%'��iz��;�`4w/�;��P�M���7�Z:�А 2Eiq!n��]��l�Մ�\z>ٸ��p៟Ƨ[�qŷf#�ɛ��o��1�����?>޸�W����L�~�����O�>:j�U�v���,�8L�~�s��G_>2m�<�������ث¹]fQ����������4s;g7=����Q>������� �Ì�B4�Xg��\$�ci̱��aaH5�*�ܨ�:�������֭�DM[�nM���}�����Љn� ��:�o�cF������[�|sn�m�Բe�\t�E����z�gb��t5�w}�������K�n��lJuC{���X���1u����nv!�	܉�b����$�Nܮs`p���v�J+n�=Q�i�hdCRJ�}y�z�X�d	"]�Ub��I���y���T���n��b,z��]�Mh����µ]GZ]�q{j]�݆Fd�I.ں�Z��<-�B1��kE��Ivmw7��Ov?_e_T�3|lhb����n��˓��������'v�Q���4h��cCwA��k; �d"n7S�F]�׺�?w�˖�uΝ��C�7��sO?�O>��ǲeˬ�����Z˝+Ӊ�L�ٽ��"ww���Vr������%r�Vm\�JrP��p0򷵥'؏���@q��\�\�����c��:��_A��Ҩ�+;��Oִ�'�����̺���3�x�۸mθr!��4�Hmi �<2�<�*�v@q����q�϶�����K���]:� ��P]^��{�[�>y���3�r��B���:�F}֑5�T=߼y3~��`��� �h���4� A�ݰ��w4�lڌ�����͔� �Y�f�%r_�`z��l�fK]�����sK���!<j��߰ȝ5���S74#uC}������l݈ne��s/�DI$�@YC��!�v�C�-h�PEA;�����ݝN>y��u��с!R���Һ뮻�׿��}G�א���e*	*��bHص�PE���zi��S+a�BaE�nǭt���.	���Ʈn]Pn�h��3K�$��݀# ��CX�n9nGB;S�N�{?K����Z�ݐfW��~��V��]�u���c�������.�3"q�X5��u��<������e���Ƶ]]W�7� �y<��د-l�	�v�S�<�?Ye	ݛ��@^�����?L�Ά�tB)�DO�c���c�qc�V�����}���7��NN�D�V��'����L!A%'�t���1��P��e?�H-�(n���۫��܃�.:��v�m��L#��+��B��D�?��c��z�r��Žۿ���p��`1��l�?�����n�%�qh-��t.+A�cf�&4�jci��^�f(�a�<j�Y7곎l�'򼮮���Z�
�;������nn!� :lԍ�_����a�G�� �X�r%.��b�p��֭��N�-uE_c,��uJ[�S��k�����;����Z�%n���k���[[Zp\�}xd�G��@w"+`����w�y��$��^�Ђ��U�A������ rǁ!�.�'���w�	��W�>?e�u7�������hFo��k{�m�|������kgֈ[���Z/���N�̉����e�:���Vl�퐦vm��k���ѵ5�.�C�/	���.W�|���D/L�vm�֋�������F�0v��7+��!��)��=f�� �D+$�C��u�)qm�n#gk:�(�+�p/���uس{7�\�:'�|UUU��l�^��QM�.�;Ye�ݳð���_YܮzP'r;3r	���#����Α�~�&|R�����@�䞧��Iq�ͪM;p���]�>�
zq�So��O�u��v���g7?�K�z=������Z`ۮF�m���v��Ȝq�a�tH�8�~�1��O��BHO��F�ƈ�jD>s��B4�oEqI��v�qo����υ��]��T#�,�9�"b�z��ЀK/�+V� A�Qٽ�5�s�U � :&E��7�R�寿E�X�/o��6���J\s�5�ԩSƅ���S�[ߠ1�Bd����o�g޵ݒOp"w����ꆼ�ݳfx���3L�7�6 A$
	܉����B4�ׅ$���h��"r���u�Ar`�|�ҥ�+���/-���.hƎ��Çjߏյ=�`=�ފ!a�vM:[����sm��wm��Iڎ=Ů��[�tN�,u��v~}LCޞ��r�յ]��1qmwo�5�6е��%��$vg�ܿFH���Ǖ���<�=V���|��Cjd W]��e[7���eC>�	s�X���%ر=wExDb��~*++q��
��Չ��.?G%a��5�]��I,�����E�vM�ud��T�ߖ�V̮iţ�)�@Db�j܋3�\��ߙ�o�4Qy��'�Ꮛ_���l�����Z���|i�(��Ó��b��:q���IY_v�˵���<�
���; �|�{�tٻm�EQG|V!�9V<�CY؞ͣ>G#�u���V̟?˖-AxQXT�1��Ð�Җ$� RKe��8d0���������_�~/�"�N0�<�%��X�)���s����t5C[����n	�պ����]/��lDeY��K�=�Ty&2N�J6 ��]#nW\�ei�A9)�� /�����_Q�9�2�-�� ��{�=\}��طoBG��}-煲N�a�c�#�L���M��ڮ���յҙ�S��.'~�vY��N���r[9N?�v���k���q�֬G������ns>����s����1Y��F�����`�ُ�8��v�����NM�6����k���o��$M3�s
��	m<�ùI!�k;߯rc���v�y��E�~���e������Ժ�%�[n����8餓2��ʤ���ا��KXy9�&�9�s�FU��{[�폃���;6��>C��r�%"1lÅ~m؆k�;���������%���_v7�� ���S��?��u��~~�Q��YG'����p������@pl�f4�<6Ɗ�����{{dZH�%�#=�C/�v�G8�ٱF}�F����7�|3�~�i�=z�Ąi�ѹ�ADn�~#}�����^{�?�
���F�����?�AJF��l�%�"�0�{���0Tc,�����}�5B� ˴����B���]7Z3�---8�_�1� �gFu�w�(..SE>	*G�n'�
݄��P��+Bw;	%%�\�d�w�JG���?��S\xᅨ��AȰc�9/5B��-l,n�,��hPvM��kD�B;,��mՋ��0Uq�:gx��Fl��.x� %v�}��#t��CS
\��vnx40M��Fb���JqM�(���>_Av��fx��vS�8�x"�;���k�C��]=���}�8�Lӣ���M����ekjL���4�6P�p+����\+��ҝ'����,"W�>m���ۇ��L�y��'}۶RҊan��Ȯ]�bڴi�gR��{&7_���M���9NL��ΰ�m��=t��C2�����G�������������>߉�f7�;�F� ��'����jވ�u�L����V�قo��;6m�� �i5�h���%���vχ�s{AD��ݣ>g�Η,���~.A�(*.��q�bȈ�q��� ����i������x�o��~*"*��s�U3��׿��H]&�ꊉcI���b�e�4�3�3_#�k���=,n?�u�(.�RݐՀ�vlƤ~C��f���Cw"�[BC�������$�Tn�AA���������ޮKT%!I�#WE�۶m��_��>�!ӧ?��D�>������ 8?�����+K�P�v��FT�Jm�\�����R��.^=��r����hp����'͵]3��$��.Ϋ���.']���x��έ���F��ڵ���p��#5N�硉=�k��=L�6�����!hc4u}k>s6�����n�/�{]R��n��r>]����������?�^y���	6���_�?��=ztƓK��MhɎ�C:r���eX�����$�=�nPv��������=�`�_;iղ�'֚xl��v#������A0��H��J�9|��˯�(O���}~vڌ�����m�Z�� �M�ʲ�Z6����1��=���uuC}�0�{{�G}Nv�|��O��nA�`B�#�MF��rA����Cѫoo���ױ���	l�g��>g�dS�0�uE[���ٵ��Y�/,������eq�m�řbEj�Q]ܹ��=�_�&���FSK�o�%����<����F�����'�d��B;!%&��\<U��v��&��T*�E�HU�����%}��G ���b��2	����M���GK���DU&��O\N$BUt*�����{��.�vy]ൎ^�=��J�N��Ĕ"�vqY�g�r$ߵ���MH����'���ihb������n�c��#i?T���i��I����*�V�i�Mb���~m�ѵ]����E��~f�6��5�.�6��q�/,,�Ga���x�n����ĒV5559�tJ�o_G�?�IX�N�^Cڂv1iŹ4pN�m'�X]��n_��zÊ�ɑ� �H.e�E "��9n0�z�(.
!�a?��~{�;yr�}����w>��Ͻ� \f�ۋ���(f�X��~�v�n��e�{ �v��%��k��T�ԓ�_:����K���,�F��)*.�������A�Iy��8*���������TK \��0w�\TVVb����f^�.��cYF��g���Y�U+��c��p}P�D����h϶)�麵{���hiiŜ�xtU�獈�@w"cݫM������so�%���۩]NT���;���v_��Ƽ�G:D2*���~X̛7���:����O�6e�ʴ�̵]'�T��d����ku~3�O��P�nq+�gXCTl���4�^+���k��rL�޵=��Aq`�v�ێ�ą��ŋ��vIvm��|�l����x�ͮ����R_[ǆ܆#p���"�,��(�caߐ��X\�}���F2�����~��{Ӛ���ǋ�΅�;s�}[l��4ͱf۽D��gajڨ󙦦/ݱyC���F�z��y?�>^^�b���ͦM���n��&TUU�=�ēM	-�|˝[��uN�;2D��#��B�;a�qqg�!�-���-�!� �e� "{�2������~���־��_��g�O���;q�5b�*� x�(D��uV�Ppo�e)�nX����������9�5�l��������+�w�^O��}0��)V�pݪ5 � 򛰛{���kؾu¦���]v�5��ȑ#�R�Γ�Z��1�S7����j��z!���L��Q���(Ϧ�1�3_/�\ܛ�o���C��gt3;��u$����P��%�Jr�(��]v`pU�DU���˽��a���D#��)�J@�}	����ǳ�>��a����b��C�?��ƵP��V�4��k�j��rm�Ϥ�[��Z�fZ,��i��fDTۢpZ�'��q����������a;�z��Wi�Z��1��%ϵ��A�凧��ڮo#n� Br;ص]8^4}����d�m���9 �p�2�e;�aM�_ &�v��-lcbE�cf�!Æb�#��k�.c�ʕ�ꪫ,����ҬL4Ų�d������pn�Vq;2���&����U�ZN���܌jM,Y� �H�:�� ��`�!��eg�Si*0����7.�>X���{���A.%��z!g�U$	��q�[���fXќ۽��M�k��HG�q�����K����&Z� ��_�;�c�YX���x��w��A0�o�nc1�{���3*f��Z"_���	9c,�nh8}�źaA�^X�&:����{,.�������Z����i�[Y�6�G[a�ց�NJ��0�!7Y�sm��W~�����;0���]~�h�"<��� ��=�0q�TTt�}���sj+
���?�y�6� ���z�`��5��b�J� X�����{	x�������v�^��˵J�����!��4Vד�Hk����"i�]p�v1�3/�sh�Eqm���nv��&����>֔��v�җ�3�/��؅�H'n�쳺����Wq�VH.k^Bri_�ɵ�	)E�����������&��u�X9S��h]
Є;��j��~�C���g�Λo� l�o����o������V�]A�����'w;a���OVX�GΕA�����5����Q=o? � �HU];� ��3aD,��l�����
L�~ӏO����p_�y{5��`1�[@���-�[ߊ�bo�vOq��n�������Y;��4��&�͑���T/��ڙ�}Æ �h�C� �`9={��/��]�;A�O?�W\q�U7���["����YK���	axG����>�uP�O�fh/�]/�k��������Q3tD�]7liه��U �X �;�v���;�P\\�80��0J�цԹ0x����줔����7a�QPA�?�������`��gب�=�P빌�&?Ln�v��+z��"r�5��e`!�03�mլc�iU\�*�U�OMԵ]I{��)n�c������ ^v�T���P����sC3���څ��<vg�;���S>y_0����Wi�{6���p޹��cP���\��(m��b�v�uyz�}�\�q�ǲ�󰦍�/���.��v����h���y��&��)'c�C��Ë-�g�X�x���p��M������X�s���WF�I����	���'��_7Q�2�ޮ��<����Xmt����	� �Օ "���/=��r_�^*��~�U|q�!	�u�o಻�����9�_!�v����ݯf�<��a�X;�cy���bzs,F*�:�%z�g�---�7o�5:A0��	� B�KeW{�|��J|���q�f!r���~�_=.��2���h�'�j�:c,�t56��{�uW3�E=|%��,
�M� �K��y���5�o��
	܉�rx�"4֭��9�ǽ�ׅ� ��B!���/�&�d�v'Q��b'���T6ٔ�Je���>��JR��O_8й��fi90�H�k{���sr3Sjc��T���V�_����R�v�vN��S{
۵Bx9&/�vS�3m��ܼ��y�rm7�MWT�l�\�5면K�k;?_$��������M���=���.�^��|e��ej�U�6
�Fخ�l/Z]���Q/�ר�Muy~}��L)�aÇ�����=�֭Y"�a���7ߌ�}�b֬Y9%fO�?��gw�92�U���a�����JT����M{vcVmw<���AD��Mw��$cj{㑫���Υ�u�
C��W_ŉ�G&�ρ�m��g�i�2��Q\��h	���~#?�$Q{ac,�v���˵C��fMܞ��]2�H���a�X�� ]�`⴩��C� ����6u�X���o��M�� ���z
}���~�m�,���d�Zy�K�1_?T�^�B�z�-~o3�a����m��R3�����Ë�⣂�8��	܉�Q2P[���v9)�9� �P����ON9mb*�$��l����[���+���$��kpđ�QTT��g���#�Dm��H��R#Ƅ���sm�*��
���ڮVUQ�:�-4��5XO������{��n��bqmW�����׳���@\�<�}AZ/����^��8_���}Í]�A�	�vV����;!%۵]����Rn^�z#��<��~�w��q��Z��i#�Y��&���� �'&n�WL�qη��7^}�~�_օ.���$��W_���jv�aJ̞���_L�#wHE�����:���î�+����c�As����-AA�0��'��Bh�O�)�nF���!�a登~u*�L�P?���;�?����A�9a���%%%��ݯ~�{�"w�+�׫n�-j��Q��G2�?���X�h�1pH-�<�:^	� "^z��Y_<��&6|�q��Z�?�r�)Y#f��|-�U!��0v;�n�U3O+����|�P#l����u�����mj���xj� �`�U�6N�5�I��(��B�D�΁�����5�톒��$l�Da���6�}Ē�
����f̝;�V��߰cm��0t���c�ۃ���E �-�Ř�����R[�4l����g��=��i|���W��!l�
�5b{h�Ŗ��(�e����Js��d��r;թ\��@r]��J� ������몾��5�h�Ь��.�ؕ�Hڷ�Ⱦ-�$��G��c53�5r��Ҿ�k; ��S�=�,+�k�܋�Y��6r<��uOӹ���s5'l��n��B폩ӧa���X��Cصs��eϞ=���Kq뭷b��Y�tJv�A�K�#������D�)
܅�F�~P����bz�f<�P� �H��]:�'L����:�H̹��W��n�/n�TZ��.:3�M��u���׮Z����QAxQ۽��ִ_O)5�"��aa�S�7�
�J�0�l0_Cd$Cl�|�&z_�t)~��߁ ���0~�D�� �H�eҌ#ѫ_K�~`��3ƚ?�e�u�Gvx1{���ͧ7�r�u4Y\ݐ��}��H�P7��j�e���Ba�g��}�z��Z�M��&�Cw"-��Tk�����E�CH���%�x'�{Ȃ7�t%���G���KP�X����H���bd
��0t��� �랬嗔�b`� ���a�⛖�Q�?�ٽ-��	��HZO�v��TC��=�h��k*57�D����ؿ�}�[���գ����O���ʳE&�޵׮c�cj�=kk@umwE�{ڗ�a���K����߷�ِe�564�M�W��5=����F��~'>]�Z]��צּ0M���D�s��0;����U���U�3|P�T���X�u�YW�ҲNڮ��ZYe���M\���G+?�ϧ���M��YF����8p� �����J�~���?A�,u�l�|+��mFqQ�FA�?ނ�cžt��[���wV�E�(�;���G��Wb�σE��ߊ� ���%���v�܉y���n@EEE\	�lJh�ۇ�}��;~���]N\y&�"�v{�A�V�����$�l�;{�P�S�k�� � �g�%/��F�ICTD:8lH<tE����vљ����}���p�Ջ�}W��îa'tى憐֭������a�h�ŋ����џ�ڡ"|w��:q{���td����?�F�ۿ�����=�,b�
AD�8����y��W�4�������+��m�݆!C�䬘=�X|�P���B�w�f�ꃦ��]�ٮ!��aj�n<�;1�!����H��D�@�
*���d�ށA�k��n��?I���ʄV�E���]w݅%K� ��d�޽���*SɶL�{2�_;|(ƌ;���'�k;;�*�wCIiI�"4�N�e��rϙ��_� �S����.�T�B;/�mX6��}�7�ك�޽�]ۃ��v���J�]�d�oݏ>5���((�՘���]9������_d���	/L�Ɔ~}tbg��4�bIl__Wg���^]-��S�)��/�bl��#ܚ9��(�����͐c��ئ��������C���؎���L�|�p���6nBE������n�m�{N�nY�2������6Kx����X\��I��`wӰ���}Vs\��KwR4\�;�n5��PVV�����0�e)��04��x��3q��ч8}��*����I�o3v�axoŻx�ɧ�^?����gɍL�ѿ���vg�e�~c���[�+�W\Uȟ.��L�!��;2��aDqd�v�MV(�*�mD���=E������"�:��Ž���[� "�`�֘�Wv.��~x�%%"�L:d ��,Tt���x������Ƅ����k��G��V�ͱ��а�><�s��X�C4�rM�x�,YԮ�*Y�ꅆv�]L��U��m߾���<\"�Xl�|^��Z��,w�	2iX���LpسOo��|����n�d�]u�X��e�k�km��;�2��Lo�L.����2�*̐^&ם��1Xk��'̌���5�F ��ٹ;c۞��z}Scfn�ϥc~��a��V���~߰ߏ�]�`��ڙ�ms�)�477c�ܹ�1ssOTp��Qk�"FDN�j-���Y茱���a�F��,cYm۬�a[[�qs���ȝ���7������xe������H9�*t�T��B,I*>A�&�D����������O&D���O~��SOY�d���2��n�Z~&�=�峡���:��(�E��X����c5TH��G�*����l_n����qS6��N����[�.����X�P!��k�5Br� V'�5�y�27��{Q��l��]#�Ո��mUq���`78�Ķ�J
�#M�־1EVH�*h��l�i�_�|�Y�)��~������w�I2~?Ҭ����\w�v�s3���`��=�]��=���~h����y��^�$���qG�Q�8Ӵ7}�/��|S\\�OT�e���i����#�%;��ISnc���k^�	� ��,��ذ�l�N���-Y9�h�=J;gy�1���w���.&��]���lʄI1�v��B�ؾ^��I��=oǐ	���駟F���q���	�t��y��G��ud��
?
\A;����+g�A3�����ĥƑ��ef״����HA��{{u�OO�x��'�w�0w��M�����/�:�e� ������W��qC�&�σ�]�_��8���B��v*KЩiL�s{s,�^�덱B��]�:���t|�TW;�IW/}$k9LTĜ3W�\�Daۖ�ۛ�23�Eii�e��X#�dj�������f�u*���G�g�^q��Ď��A�X����򙸞�w�v����3��3��m�}��]*Щsfn���3���Ϸ�oMb7t��w��R�<}dr�3S��=����2Qr�g��[6m�[�,�jxe�J���"S���]���X��2�K���u��u�]g-+��l�%��X��#����s~���ڡ�o�Ż�[�Y[{h�nئwp�k�e�{��z�&���AScސ��H),IUޜH��@IX�C�n�!u�*Q�0�'�d���|�Nt���{��L&v��R٭�=];�`Pq{�GS��&� ��풟��<���j�Zi�-�V����}Z�US�S'浻�������eA��>�~==]�u�$6��#�0e���i�5qX�N��%�E������� ��ɭ���&����:�t�{C�F������['nw�<r�r��M �k��e�x�����k|,��&����3&C�a�۵]\VP�vmD�[�ӝF$�ۛѶ��t6��Yj����]�������K��� ���I'���	(��R*�QX������k?x7w�}~�A'iIJ��q:'w>QŦ�ݱ#������@A�\s�QZ\��}iJ�y�����v+^�p�H.G���/9她/n�TZ��.>3aq�_��~{�S��A����;Z	�)Vpq�X7�넺�ew�ڡ�9#���#֚#��_�`^}�U�K�^=1y�4K�NA�O�~�u�X��˨�1�"r��^z	7�|3~�_8f���w�Z��1�>bu;c,�f���G�cq5C�^h_��uB^��F�=� [����	܉�2���cKR�%��$����5Ġ���/Dsqg$C(K�Tӓ���m�p�UW���D~2pH-�O���Im	���v��@�v�8TO0�vA���,G#�׵ݐ���SbJе�#vOq�S�]��ͥ��JJ�cS�·�Sd�$�t��5�a����(Z��h��R��NX]/����@[������~�ˎ�9���.���m"��uN�Y7eWn���gB��M�bM�;8��X>�F�,���pmW�1�x�y���Csޓ��n'�>������d�x��+�"<�ȗO?�C��ǞH�]�D���_=jjj0f̘�K@%�_,��m��g�5��p���>䄕��Ҹ��!A�nZ����'��e;��膃$�!� 8���s��R�S��}Q� w��8��w㳺= "9?a8���i(.JNq�݄2��d#e%EXx��0eTb���ث���� ���[�ƺu(..�4�ҏ�vjwj��zc,�v(�<j��kH�v���&���x�KWmQ~�p�B<��� 򗡇���G��� "�uꄙsfa��w�����O-Z�A���NK��=�����u�.���P�������=�wq���ᑞE���!r�[Bw� k�s(Vn��?���D�8�O!wĞ���U�%IŻ1�ɩ���DU���:�)1��7ʇ9��Y�D�Q�~�>ij5C��,�  ��IDATE�c%���t���m��M�!�k�( ���%����Jۣ��C����DD�o�s�ļv�IrmW���5b{@���ĵ]#:�����.��u>��.�vx�3�?ޟ����	�qe>֥�!]����ݞ�)���daz� ���y�S�lϛ>4�A�gbqm�۸=z�$�1#;�|�̵]�����i��j��1I�t�y	���|�Ï8�z��C�?�];w��/��ك+����z+z��v1{2Z�����ב���V�k'�����i'�L+Q��3��� 9�7�ٍY�Uxv-�EA����q��p��ӧ�^~6N��/�ݴA$���q���'n_�����g����"�`�F��[}"���+����� ���2��%�EL��b�Y������ uCK���b@���^�d��1_�k�̵���n��0�	GNA�� � �l���;~��{��W�ak+��㦛n�D�'NLj�'���xbvtK�1V�=�1_;�k�|��wqgӬ�ad�g�-d�#uD�^��a�uÑ���Q���������H	�@m�s'I��P�T�D����$��\��R`�DO:����J�KP=��� ���z�t��߰��������h-��#ҏ�o�u/�{S��TH�)��2=�k�6��N챴���J(�vm��]�j�H�k��/�����{�csmOf쎰�;f��� �C�I�.�9�gݔ�]+$��3��O�/̔��v��)����;�%'������,S�G�G���q��/�v�D]������v~"yq����o�~��O~�G��0>��#��ڵk��1���Z����U̞H߱����s�{�g{��9	+{>Y�n�������`��d���ɨ��)$�G)Qe%��l@U��knAA�l�~��M��[�2L?�6�<#j�-��s�=��-�AD|�2}4n���(%���~Z��pÃ/��0���f1�����g��v����@D0Nl?���5���4\���7�*�������ꆱ�cE7��MKU=1��R�ߺu�Q��A�Tv�)3��sEgAD��w@w����K�M�Xy�޽{q��W�[n���B�k���1�^bu;�n�W3�녎������a{�������=�=�
O���!�Bw"%̮-@s]�%6qSEE1&�ć����tI*��#r�%���ǻ�T;0����~�G���0i���;F�۳յ]�Ih�*}�u@�>��6&�=L9v����R���O������f=3��.
�����c2ܵݾ���2��ɢ�d���䷕�@�]��]����b���rkn���n�����7ͨm"W���M�umW��T��G�GD�R<�,?�k���L.ve���K��w��ƞVVV��}�,���X�or��7�.]��o�?��O�"`O��=�>�ik��&��s¯���k �C�V^.�,Y��c"{������d��� 	�YA��-X��A���z�����s0�`�L��貳p��Eh�Gn]+_�9��)I��c�'7/��/�D6RԾ�w��T?aXB�0�>��	"8}��@����D�VX�c��n(
��ڡW�PW+t_�)7[�^��$ې*��%Rglhh���۶m�1�M<�:�� "[�ܥǜ8o/{֮�_lܸ���x�(//�j1{�5����uR�>��Y����.����P�V����C]���Yvrg��ףW�A��H�?"$p'�NuyƮ�(��'�
�$�޽]��RD��4p�����3������˗[_�A��D�0b�(�9�0�QX�\��sn���1j��]����b�T��+1�ѵ��	����n@j�^�ve�힀�n��`
�A�������]���]d#���PHn�o��_sG�rw��o~�!�)��y��/����y�@\�1�VL\�@2]ەs�&�hm����g�a���?������~��1t�P|�_L��=}�2�_[_G�KZE^��ܽ\�CQ�U���;KV��mڱcz��[� � x��9W/£W��1���3u�@,��k$r'���	G`��N�����mg�u�X��H���-?�2�L�P?�=�<��δ�=h�m��B�l�%��5D^���������=�\�H�ks��MV-0���u���_o����?�LĠ�C@A��:�����xD~��o�w��.����@&�&Y��CG,�X&���y��puC��F�Kg���j��Ԋ۵uC� kF��x���Cw"����;�@�v�Ђ�I*�{�_�� @�J&UB�t͗H[�l�W\���&�CaQ!&9���h�	.l�V�v�V�_/m�Jb�B1E��d*�r+Ź��@�J�ib7����{�[�>���z+�k���pcu�[:�]��5�۩�kYo��ڕxwve��m�
kyvu�|��z��@����Sb�F;חt�"ޭ+ƙ�k�!F�x2=����$$�nK�k��I4�����I�C9~#��H���y8�<߯���=� ��TU��S��%�h���x#�܆��G2g�s�|�	�۷D~����Ϸ�<�0�F�t;+��G��qd�q�Ǣ������n���.�z������<�$��d������莃ts
A!��iκ�,�曨��=�<L��׋����=h��	���'L���Iж��-��Z�1��f#L�~�_���1:�~n_����9�I����~�8�s s,�Q����'n��V�0�9#�fX:�A�~�����'�����S����� � �����Cѥ��zeZ[�!�x���1r�H�~��I�󤻖�nc,��ϲ1�+n?��!m�PW;�	����>C����.$p'���>E�'�u(.�$�4.�k{t����T����&��xS�p``B�y��aÆ ���8��е[%75",n��3����Z y���\�j"���b��^��ٱ{�'ku�5�ve�FDx�!n׶�b�tm��'2As^���B;S�W���-�� ��Ϲv�]�֟(qn����Y�(U����	���τ���t��qr��#��}�����T߯f�����g��O2�c͞��x�����ԉ���J�y"�h��K�Qo�ќg4Ǯ��nu%�@|��7D�������97��m�sy��U8��YX��;��Ï@���͸��p�M7�gϞ)K@%Ý!��b�Y���ܰ��-p����{$��u����&�tɪ�s/q{$YU(��76����z�Oi�A� Be��F�v���ǵ�B���@��8�O���5��ذu���N��_?.)}����;�!�j܋l�����/��3�$��#K�#q;A�HQ�@?s���B�ݰ@��۽=h��5ȂS/�oO�x=u�D�x�p�w��/��}��(�T� ��0��'Oć+�Î�;@��^XSS�)S��]̞�ZbPc,C��o�E[�S7�����.���1ƒj�^�?����E��Q�����B�$p'�F��$7�x;���Cz%���T���T�k�_�*�O�%��ξ n��v��� �^}�`�Q�PT�������\��`RC������Q��$�?�صB�@m��99��V�]ۡ�k������	��i��p4��r����	��i=M[�-�Q�m���@
\۹�=ۄ?y�Fÿ_g����.�F���}�����u#��?��ǀ�������G��ˊ�՗�[�����#�"�>F�;�#��3�6����N���E8���ťK��g�"?ظq#���j,X��r���w�lrd0�O®u��Wwq�'��d�=Y%	��뢦��,�]{I�NA�lܶ�]�7<q�7ѽK�@��Wn�!^X�6+�ܯ��9l޾�	���_�1�<sfR�{j�G����b_�d#l}�K�9��'�Ͽ��?�y�.%I�s��=��������O�.�]���b����k�D�X�f��k9p ;��Dj8�GL����� � ::�7�I���O�n�Z�3x������?����O�=��X�K��SJ�5/����NB����v[�λ��5C/w������{0���]K5C"	܉�q\�����J�*T��IHRQ�T��y&���Ɠ�>�{�9,\�D�0b�!3~w�D��������3#?���L�k�����ʵ]��K,�YN���t[��mL����k��[�,�6�yU�z,�G�r�:�k��;�>V����.��z�/.��D�y9�K�����	��!��)��=�k�sN	Я���C�ε]�&�6�va>�yB#���qΝ�r�c4��ؿt�H�k�f�	ʹx]����ie�6<��cQUU��=L��<��_�=�܃��??�T2�b�#�mE�3���a�C��*9a庸�n,q�0�bHVqw��jmi�1�Z��j*�v�C��\�\��� Ad�6������^�������0�HyY1κ�D�	��y�bo�;�|���,ڲT��~������&$�ϊ5[�����e�H�����ϳ�`"[�.o��ܵ^[+�3��?D���� 2ژ���U7v:Oo��#��Yɘ/H̍��֨�uuu �v̌w(F�� ��%��τiSн����U� r��۷c�ܹ��{YYYRM��YK�Jc,�uC�Ktq�G��j���{[�������,6�{��o�� �;�$����a#��!}�TZ����$�d'1I$+I�7�d$��90\w�u�#.O`���'`Ȉ�´����\ۃ��|��ѩ��C+��,��*a�BaE�nǭ�+N��[Irm��h�S'׋r����ůlcu��}�79������v뮄�>'ӵ]�A\w�h|h�C��R��4B򤹶s���G��͵=2��i��9�v�db��=�~ma�N //[�ڮ�[6h�����c�?ǻ74yl5T�6�,ʷ����N>��c����j����D���rfΜ�Qz�	� ���VLV�� �uU�+����?a�9-Y���Ѓ{wlĈ��x;ݐ��̙4��kA������>�/?��;�}����ҴQx�@���q�_��G&.\c�+���߸����o��|ab��6�V�s��Ջ~��ϕ�݂�?���[����8@�w"C��݌杦�)�}��m�%��l���!{΋/x�,��Ea��CetD3�x��{��?�˗/���`��3Pݫ'� "W<|(:�����^���V�ϛo��;�?��O��'��*���ۖSRn�Pg�Ů��i�U ���5��\�Cj�PW/���5Ö�ݷ����9`"9�^@$涷�����Ib�un�=I�ﾐ�$��lIhu``��ܹD�S�~|������``q;|���l�c��ipm���Ԭc:]�MgN�?Y쫛�����"�u����Q�61�vW�.+�r"+��k�</�|���wm�9bhe_��=r#���P�Ӻ�b7�IB�n�����|�������;����y�Br�1e��k�t\�; �ṮBnmL�^�Nx�yB#"��qΝJ?�\�u���H�]�����D�^�+�@�6V?���>j>#Sl��{�޷__����o���Dn���ٰ�������I��=�>2�6�#��h��{;����N�#������j�U���Nu�����|EA��\�s�y�_�5K�ۑ��'��k��q"�t�T��.>SGL�������Ó�}�l�s���O��|���3~x?�a��e?�[��u�|���x�h޷�j�S�ƺu(..I�n(��,��Z��������uD/�-t��|��O<�ŋ��JJK0y�tTt�� ��uz��cN8���456��}��~�9'�pBZ����RUK��'��8���n�g�e�Y�Ю��hk�|�P~��6�؄��C�c�=$p'fXUa�IELR�
cb�@��������^I��lpcHgb�~�7bŊ r���v�L�m�n�f�Gpa{Gvm�I�âO5LU(���N=\�#B_^�_G5vu��r;�E���Y�&��z�4���c)��v��]L��:��*���<յܾ�h+m�f	��K�{�إ�#(q����׎ݧ����c^�8�-��\�+�k���^q"i��J�\o^�����˶��:�������
�})�qͶ6ܘ���cW����� �����m���.�ML�*++q����<��>�n�8[�l�n�dnc�a��ΐ�dT��+���$�,�v.i�'r�'�dG���<g���wafM���dA�����Gx���+�����r�����H?x߉���r,��l��;�v5��7�y�>؀l��g১N��a�!��&��a���xqŧ�M6��A�~%��&�lCKH?�s0a{��@�!�G|���YvJ���mRe�K�d�����`�� ��=�0t�p�AyE�ʮ8�s��җ�c�6��G]w�u<x0���:`�}�2_<m�5ƒ�^5C�5o��j�^5� �X��{�ctY>&c����D�VQ�����+A%&�
<W�JR�Ȕ�=]��K�,�D�SճG}���`܃����c�mg
��ԋEe!�!�e�Ipm�W���ڠb{��Ib_i��Wa��ۃ����x�����5�����*�1y�E,�qm��	sN�´d�����MSE�q���}��G��h����cwmO�G+$��3�M����ř�N�v#|�����;u���(ˇv�|um����v~ZiI)���x��g���/��m�z�-�~������c�T$���B�j_;B�J��b�k|�*,x��ŝOVَ]�mFyqo4��ʆ ��f��+-��?��� ����Y�[��/}D�QS��۷}>Pӫ]~��p_���Ys��M;����� ��
0q� ��3����t���;A$����\׀��OS,�;W;�j���=H�PW/t��<�l�K����k�.̛7MMM r�AC�`����]O�|A�Gq��ԣ�?�{�u�_�)��f��ݘ;w.n��6TTT$\��Uc,G[y�����B�Цs��ŝ��"�B�fشg���zD�Bw"!f,D��z�����ޮ^09I*��,&���Lґmn~mW�\i909�ACc��I�1�����"xF�sm��k{X�)k,U��{`�v�O,��ж�d�m�M֌j�4؞�1�z�v��sU�,�vA�m5zP�D�]�kcw&��sq\L�إ�Ҏݯ���L�6�vs��p0²�}�Ǫ{�����x#��<Q$��C�GX#m��<��ˀ��s�o|NL]��`�s���]��/����~0<�H�F_�憄X]ەx4�M��>��P٭;�||�u�L�.<� F��9s�dm2*�|��̑��~}�����b�����l'��]�-[���hii���6,Y�� ���W��K'��#s��'a���:�h87�/�v��VQ�\gdMO<x���SU�p_l=��Eؾ�c��t*�/N==+;�+�G�>��ӽS
wo t�X����X!�~�=��\3,p����X�xj���'c>�9�Fgu�?���Q���-{�� � ���q�������� �T��trl��/�8��_�k����c�]�����ۣ>����vq�j��QҼ	�%}��B�h�Bw"n����ʖ�8XTNJEN81����e��D�Tn�JLR���$U,m�:0̟?��� r�cFa��q�s���AT�\���M�� �����������K�mg>E������{	x�NW�����sm7x�4�^P���	���_�.��\N\ۅU7����J;e�s�`�Q�cMn�Y�Թ��q�?M�q���n��\wAc���wԘ<��A]�M�4�<�]��bqΝ�r�xLu���2���2�ڮóo�h�O�.ە�#�N��O�|�T�����އ��� r����a����R��e�#��*<�;wY�F���)9y�VV�#sa���n9��~#�T�bK92A����k�Z^���6���b���3p�/����	yo���CYIr���⾋�L��{��5��u�qoǸvb�oQaDp&2 ���8㊅ �D9�o+��ڒ�ޮ�٫n}�g�:��mfX��M�|�93	xꩧ@�6�x�|�4���AA�a���Ν��˯�1V��裏bԨQ��W����'��bi�1����n�����cuq���1����8c�-$p'�f�@���PR�{{d[Ĺ=SI�l��:���p�7bݺu r��>y"����!�p=���E�:���*:�y�`5�{���0Uq�:gx���k�(�Uc��ĺ��9�v}[�@V�Ƒ�$ͨ�@���c9�LM�d���q�N��0��Iqmw���&�ؕ��?v^!�Ǥ����ʉݧ���L�6��Ո����r_�]�ݾMi���p+���h['��E�@�GHν���~m��k�]�x�`��"q��(���nM ��k��:-���r;!��wذ��q����{；n��a���q�UW�O�����J*ś�J�X=X[�#�;��ǫ}�A9ae_˙N�J������{6��r�$� �s���-A���4�!}�,��7�}���"
��\p������|r�3{�p���SQZ�x�g���W�=��;N���I2&� �H�!�Ѵc�����¨�vYܮ�ٮ'1�E�{�t�a�fX~m�����{�����`ڱ3QU�AA��T�N���_�ĴD��4sÇǘ1c:DM0������ȝ�Y4�j��"w�nh=صc�vȋ�[�7�o���l��	܉�`C��7��h�qo�ەU|��+I�̾���4���F{��'-q������=��)@;�]��E-f�\ە4m�����3��*����rm��DZ���]����.�uն�A@����ۅv^�튃:\��?�2-ݮ�B�L��+�Y�)e����CP�!6�v7$�����ӵ�_(Ǐ�qmW:P���9�t}A;�r�34���t��!�h�+v������<�6	��kcҋ��i��~��sǝ������a��\p�1%�:��Bl}q�+ұ�;�	�D���n��udЋ�cuqo�ۂ1������AAѸ�/�BE�R�5k:*s&��OO���~	D��ѵ��W0��Z�_;n�����?إ�����ぃmh޷�Jsߩ� ��û�F���+Ƚ]��5�PLuC�A��{�,��a:��|uuu��k�?]{�2�+:c�qǠs�
A��{u̜3/�g)���@�&��l�ܹVݰ��2�z]�u�\3���a,���urg5Ķ6�����l="�X�V�cM�n��{�+!�;G�mž��R	纠�{&�
d7uhA]b�Oܞ�$U2O:2����Op뭷��]���t�г�����҈��֎\��刂u����]�)\۹?�4u9�ؕv��]�]ۍ��U�����d��]�7M�b��f�1Į�7�b��BL������N�4�X�n#n�,pm��,M�.Hm?���~���yا��� ��v;a���>1Y���<b�&��B��34�|�F,�������h�u�]x�j;uuPU���ɏ�{�ņ��A�&l��C=�f��ɨxWA������
7�we�sc'�l7ޑ���῜�]��PIRr	+[�>���� "�{�W�?�n�8q�HtT~s��X��3<���s����NEuebfL,�8��ɘ��9��Y������#/���ʶ]�Ի���i��H�#���~;JJJ���Q놼9�ƹ=S,�fh8�<��\7-�a*L���]w�����~J�X9L�U�s{Ii)� ��KeWs�l��ߥ�U�Dn�j�*K?w�EE��udc��my����� �ˮ�uDo'w��\��b4wf�5��P��F.��	܉���^���Q\\�8�j�vI����E�^I*х!�I*�rcH$���@�7ov��"7��f��.]���;���Nx����.���R[�PU��5�q���tI1�5�A��^^�/%v>6a�V�/�����9�05����>4m��x#�rx
���������z�,C#�v7��s��K}mr>�����)L3���v��?)&k����X5�۸�MwS ۽ɑ,�vML��¾i��ڮ�kjڨ󙦦/�k؇�ԗ��F��Epo���U!9��qo
Pۤµ=�	�$};nZ���������Ea�W�Ax�#,��#0`���AAخCtd��p���=���]k���>"w�I�vd�\��߂��]'n�]t"��]�8r@^��1DeA��O�N���%�y�c��v�� sm��Ÿ��3p�������Eq�g���[/�2���l�k ����4��;+)N�?��	d3l���۳�ݓ''�מ�|{���һ��#��?�q��ǀ�ܿq�C �x	���lG����ۣ�c��v�K?�3/n��{���H�Y9u��a<}i�H=�G�F}&r�^}�`���(*�QM� "(e��p����ŗ���- r�ŋ[�X'�|rR��T?�֒!����.�b�i���Bc,q�g��]qr�pqY�]ú"o �;3*�XC�B�0��ɩ/q����O�ŉ!LbI�lvc�4I��<{�=k�*�}�-X\R\����qڙ��sm���k�4]])��$�ڮk��̵ݔ��b�Ȋ����z�����nM�m���,�k;�Ů�7��r���K�C�3���ʾ�d�vg9�}��� b{�BM~P n_�Y�ޯ_ �\�=�o��R�����(�SW���a쬯���Y��^D�m�6̟?7�t�u��L6�,��69�-�dM��΍3�ލ��^��$��aC���wqw�T�=�yz܂����� ����NDM�J��~�FlmmDG�u�A�u��a�оxಳPեS\��n��Wp�e�D�Dl����?�N�6*��%�%w=�%�|�l���7���2}t�}}^߀��.���~���O,�Y��a`/rq��֝�8����n�sLm��{���$t�Ź��ꌱb�z�cu�a��~�!n���ˠ��1~�$�!� "6
�
q�13��+˰��u rV/5j����<����1���\�ЮF7�r놊1V�=�sHk�常kF~nڳ�kz��ۨ���11�O��m��U^"��M�Jp`��r\ $;I����1<���x�!r_�U�{�Ĵc��~`ǂ�ID��'SigJm�����'nk$�pm��r�vL����r})��ӽ\�S���_�I]OS�N�=bvm�׷�=�ߵn;G n�G~���^�k�kh"��E����+}i��z���k;�:�k��wy�����q��7����웩umc�m#)#�vq�Yv4��i��\Ѻ�	�vZ�yd(�bWVO�����6�4Sm��k{����ݿ4�Li�M�rک(++�KK_ �{���k�����|�C$�R���U�9�~����v9i����&�Z�)��]qq�$���}{�0��'�^C?� �c�|�g8�����o�sY|N�SGįΜ�k>"8��;u*���p_��⻞���|�J������gb��~	����8���sf䀽-����G��:B��{����_�g;�� ⥴(o�����#>s�>茱���b� ��l��������d ��Dnrȡc0zܡ � "~�o�I3�DIi)V}���c�Ν��k�?Ym8��]��e�1�Xӷk�|��K���������q;g�U�j����]?�j�Ņ=�J����D`���
������U�ƿ������r�C
&H#��@�QP��S���g�)>�PCB�"�  �#%��!���{��gvg洙��;{�?���3�9����s��N\��	K��T�4���O�>�k#U>�1lٲ^x�u 
��	㭡���pEO�"5bL�[����նjj����\u��<�N�wm7 ��U!E�����VS͚�#��7v�>vfitm��)�Gl{9Z[����J���]ە�ںK��R��:h��@�|��qb�?��n'�w_�{�;Iǵ�-��R�_I���vn�X�	⡖e���;�dM��o�d��|>Mݵ�;FW�x�|��q˷R%q{�\ۅE=�M�/n��}�|�XT��#�D�z�jx��X�paV���J�q�<�g�ȧ~#�����%r�l������g?G����.��Ka6m�ЊIh��� "��q'�q�_p�/NFiqr�����R<�n#�[�1���z�|��
e�wy�G�c~��A�����W��ǭ�8���r^�7�~y��QH<��&�ꆇ�/��Rٟ���Ӎ��ޅW�ߊ��݊�ތ�#�%�H�L��U����^���]3곟1Vq{��]g��Hg`����'[����/�Q����þ��AA����棢�o��D���k�����g��e�O0�r�C��}��X?`d~?'p��u�w��P5�bn�:q�`�I�ܻ:;q��"<@�X��Y>���!K$1��0�E1���qJn����O��7R�ȶН���Ӄ?��ؽ{7��c��)Xx��@C:7#�5M��dE�š�S�1De��!���O�k{̍ٔ���G˺yj��J�FخYO���Nщre��k�!����
�5�Ǘ��y��+��垟���Υ���޿��^�w�ܪ��q^���p���I���k��e���Η�
��:*/�8�m��d\��� [*K[?a��fjˆ��͖&�v+I*�y!��������ǉq�L5&����ǎ�ˁ��hH?ڑG��AU��]w�(,���q���[V#G�L��(Wb��920��}N���b�un�s?��he=���)���Hr�ˑA�Gһ�{q��^ܳ���&� ���>����}�8��x�:�.����{�X�T���A�(/-AMU��`>a���!����DZ�`��﮼w?��¿�>1k�e��r^�e���f����f�}/ZSX��W�����,��zz����]X��v�۰�Y������� �DUU����US,Nܮ�7���dq�W��W��o�YB����0_�}��Gq�]w�(<�>>�"L�1AA��}��FIi	ֽ�J\�>����kٲe���D+��X�'I����7����ɽ�3Ų�ͦ-V9$r���Dei�5�`�ƹ�n��f�Ht_�i��+nGLX�����ah�ґ.�믿�>�,��c�'f�����"��q��J��T]ۙ�Zjߢ ҍՉzUQ��d�fK�Sa��	_[�-��&�ij9�
�ڮI�|J�k;��)N�}=�=i��Rݳ�ڎ811Et�]�U1���-�w�B�Vl��|�����]�{�趑��̵�Y+}y\������8/���}�G�.��umO:.�^�{	�z�k�o����tt饗ZB�d��<�l�JG��|7]�n �sC��m�*�9��#ߣC��V��{d�س����Mt,�w>ޝע�t��bƄ� �H�;{�ƍ����4��x�7_??��>�y3��3?�r>�e�(+G ��*��xmJ��PUY�|/���Ŗ-Q�3AWw/���w����|��%�q��?�W��?܁u3[;@�}�]xw�nl�Q�rg'��a�]訇�oȞ�>�?��5��v{�g~����3��)S�fX^u`m!��F}.<��h�L�<	AAd�i��DYY���t?U`�������=�O����ڤ����?�,���K�3�r�<��#{�*�&w�g�~C��	ݻ���||���D�Cw"GN�GO]��+D������SQ���f�~��H�x,Be͚5��`����ܸq�`)@��V(c�Ce1���t�vU���k��)��G�:!�*浳L�k�$�t�5b{x�����
��ɔ����Z,K���x	��q�:j?�~w9-Y�v�����=CSW�u������J^����oۿ��{�u7�^���h�m��҇,w��B����u\rmw�SW��fj��c�8M^ʺG�Rum緛Z-7ͫ�Z!x�'�Tc���n�?z4L���$�>r��s��o��5���F�!
�x |0�=�ج6Fe��)����J���ЃZa��9�H�5�`�5Ԡ5G��92�D�asS�����������2���'��� ����[ǾG�S���'9�?�:^|g3��>�[�@���_�Ýxr�F�+�{���C:��/����+�P`���ۺfY����*A�M(+/�>��vI�^�هX��E��8�3�W(��E3,�Q���X6��G�L^Ab�ϬM�.��={@�;d�2�W� � 2�ĩSPRZ��|���
��;w��/����#S�X���1�"a��B�o�1��:�s�>�t�Œ)��Y�oh����L��Y���M��� 
�qVY4n��0J�^������UR㔟����@��F�t��ә�Wlkk+.��tuQ�D��\�g̊�L��ߜċLݵ��_�ӶjjSqmg�+u
�k;':W��b5�t[�-��&�i����Tѷ>��ԕ�Y�v؛Q��z�{\��X\��G��!�����z����b��}��H�rm��;���ә���f7���;�^M�\VԵ]��d̵=�(�J2<c��Ja��]z����k;԰��l���g̰D�ׯZM"��������2eJR�B��ؔ��h�t/c����]��.�C�UE�Zq��Ƚe�N�=o�� ���3�t����0{ʘ��g���9e9���Z�aOcN��-xs�N�#���w�_�Ԃ����ۛ��oEkG7� �e������v��]/rWG}���F{֚bA�Fd��͇~�t�h�-�܂�Da�\d=r9F����	� "[�N��G��=��WQH<��c���q�'��'���X��%�1�)�3<��Ϫ1��/F.r��t��Z�;3�ڊ����!�;��zѹ��奊���E��B�V��%r�5Xɓ����'�	�����A���꫱~�z�żE1�3}c�փ�����kD����WY:��r��sm��q4���J���R��V���]ۅ4�'#&&���|B�!��7ky	ĥ���4ݮ톽w{�]ُ�};]�u�y)�ȶk�������SW��fj��-=���f��F�������>X��]x#n��f�1�um��(w*��7�;�������6��Ι��ի���	�0hhh�^e��S��)G�l6\%3_����� ��&7T�C�V�C_�5�`��Ƞ9Ȇ�7h7Zͩj�ۨAA�	����߁G.>C�+^����`Ѭ���6�^6l݋��>�Հ|���מ{�Z0#-�=��&���ۭ}� "Y�Ֆ��a�5�,n/��s�X¨�na�ϰ8��]~6�3��"�}����������w}�pQ^Q��>y$�
� � �˨1������z�d>ZP\y�8������R؞l��L`c,��19c,n��1�_�!��yc����3f:��E.�	�	_�.FW�f�Qʧ�J7Ġ+t/�:0�6P�'���5���T#T����?��S���;A��}f�wb%"Xg�M�k;4b{��7k�������ea�.�Cܮ���-Ŧ�ڮ]ayC���)�Bq]۽�n8�
���.&�:�r)��[q���u{�uϪk���),gW]�������1Et�\ۥ��s��v���͗o�?��o��:!9����Z��Z���o�dEw��ȼk��y�u�J���#l��튰]:���(����RX�eh��q'M��g~��ttt�(�}�Y�q�8��Ss��Hl���3�}XkD|��� �2XS1/lw��9E��~��ū;�� ��w5��K���?;�j�L��?{0	��̿�݂�~w�ۑ��Q�[~qrR��:}�|�w���:��H�ie{��]�����>�"{�g�ɝ��B������C8����ܹ�:?yy��گ.�����絎H��
��$n'� �2l�p�z��#���D�CKK�e��r�JTT�����?�Krp����XŜ1V��+�_ا1��c�X��ϳ5�-T�(\H�N�r�.t���T��*a��"w�Aѱ��ӵݯ�J��S��r����'���*�V�v���,����Ҝ��Ⱥ���oTdaӆ�R~SCc��T�4�����zl[Kkdj��J�bB��8}��nR��O}�"��G��PY������V���ݝ]hkmX
Ww�j�~$C^>Jc]=�wMAЯ[V-�õ]�َlV��:������TѺ�v�W� 'ώX�}�޽H�7�����{��o��]󒅫]��8`���ڍ�ֽ�U��_�3L_��6\^M�MVC{EE�Z��e�x�H�y���k�N���J�'xd���ղ�q��C��=��9���ȿ���_����D���&�M�����m߲/<�^����,�!l���:��ް�"1�d~	��D8d�x��/[�1O����MUUn���}?���p��c͚5�?>fϞ�5a{>96��U≺(�o��*�F+~�Ag�A���;�Aލ�5^M-݋W1A6yy���s��	�&��g��VaOc��">w>�ι�>���!�5y.8�3?�&-�=F�v� �Ē��hil����>Ø�@��Ήܭ��?��9�~C�Y��/�Q}�:��e��o�������
X��]n�����\�h٬�}��Q=x0�R����a��~��}9�3s��l�9\��o���?��{ֶ���ތ���9��t�����6��|fϷ�kj��#���OjG��=_�\��{,��_~7�|3��o���	c�`��r���3����X�Q�Ց�������7dϗ�џ���b���xe�y*$p'<�:�m{7���<�Hk��5R	UE���/r�7X�7R�+v���F*�h�b�/��R����J[[n;�rU�-~����0�A֝��]���L��1M�R�:3q��ӼJE&]�wnݎa�FX�Ysm�����L�9]y�.�Zw� �v�BN>L���Ԍ1��i�Q�u��tm�Ҹ����6�������L��~�����nHu�%n���'�f�StVVHR��OV~_&0g7��ǎլS�������ob��k�w��vLS�Ѭ�]'�uҭ�[��Ü�x����K1ޮ�R}4y��G:lHdqE=��bt����}�_um��c�AĲ�󄜏��?wj���I�N�����7���s�㜼}�ĥ9�}�����x�"���A���� ?�Z�M}����>g	��$}�����ƆF�ܱ����, mRbq�.�5�_���Va~.��}t��g�v�����o�/�W_}5��N�l�,�3�D��tVJ��*^����M3����1�9��e7���,�8�m!w� "|\p������5ytB˕D�����_|D������͏��>�|�	�%�i��_�l����=�)�'"<G�����BW�?��3���F|v��ɣ��K��=ڳj��?+�Z����^z	w�}7*++֮$.S�|V6ۿX�D����ee�g�t�6�XS��������}�Y�֦f�ز��%�sU~G{������rA��}.�omi����93���[�}.޵)S474�쏶�\�ߤ��=9�?��|�η��o66���b���{,v��{,v�+c�T��ڵk-c�y��eM��Hl����}�����~C3j�U�:�������џYڔ�x��Y	�	OkE{��@%��{5R�SBcU�!}��O���*H^?�0��~�;-[�	�'i�7��2��}dq�)��R9^"Xi��|QZ�r+���uub���Ԋy�,�dK�*��v�zz�(�׏��\S�=b�)�X]OS����-�*G#X�t�B�(*��d@�|nx���3�P��M�ۻ�iĄ˦�&T�KS��q����)���M�:Hߝ���8��4���
W��ԗq�}YF.O�y'G�:I1^ǵ!�7����+��'l�XE ���+����F~�+u��XIܞ���;Ǝ�
�uy�j7��po��`��֝8����G���}C��(���z%o��c��[g���/���"��o��n�g�yfʍQ�uIHn~b�UjC���{.c������n���F+ޑ!�|�r�o����{)ƚ�Pl�@_�:d� "Yz����5���_}%�e�T��H���|���亍�w�%ng��_��/$n'"->��-(//wG{��Y4ǒ��,����Xq���Z��T��G��н��]t��7l[��FC�6�o���)�E]��O�m?��
���rnO]�h����	���~�����,���lD��!Æ�����wo߉��T���Ps��=�=سs�M������n�qֽC.��g/U�5�`T혜��K�۬�oǌ�'~�a���{,���=��ٔұ������^k���������J�h����u��^����ϱ���س��6�*��-c�g7��{!BwB˾�Jвw��HU�i�����8��C�'<�[>�	4�F�x�ݰ�μ�oߎK.�$go����-=�G�ߛ7N/rԔ�����cz�y��{���8�|U���������q�,���1q�R''v�����^r���bE�v��'N���5�)��[w�:��py�N���ݽ\�Mn�h�*І�{b��鬻#l�S+���� .�� v�:u�����A��&��þN+y�/����ߒw�1�'�;�,#u�v]4�=ͱk�I�~��Sm���q�D�^yi�K/����M(i�tm�.�[sm�>N��P���ر�cq�����/�\qr'�ɚ5k�`�|���llJ�|�gc�ΫїO��^�̱�k��>G�ss���!��*{�A�(�ڂe�F㉏��� �����51o���Dr�ߴ���;�yW#
L��_�]�t�DD�C�w������r�a�=�Ї���L�t��'p���+��>�Db�%�_�r%>���A��jv���ȝ � ����<��������BG[�D�D�x�w�j�*�s�9NZ>�zŦk~��X�6Ag�e����X��B�h�c{�r�X�1֘~f�5���
�Z��nBG3�@�5�7�`�ƅ�gx���Sh�JW#V��3%tg'o&n߳g��c��'NQ�^uo��To��5�v�d�_���2O['VS^RS'KY���g(�|>�P7*:��IYK��5+��n/�U�d %�v�X>&�Ӳ����CF�Ʀ-�6��r�tm�rU��vx-�y)@�}�-(�sI��7�2V�Cm�tǪF�ĵ�9Wh��������rXk���<U!�['�:qQ�!��Ju�
G�.��smwʉ�D���v��.Mү{<�v'�K=z�ɜ�W^"�0'	v}�uס��:m�M�#\6_==��bG��|f�~����8�n��F,ٽ���F����QZ4=�I� ��y�J�㮜/�m�i���n~��N��cC��������GGW
$n'"�9�u(��pD�}����E��%n��;��o(bpSz��tdZȞ��֣�>����� 
�ʪAX��$n'� �P5�ˏ>
O<�:�;@���n��2�:��CD���|Ay�|R��bi��B���1Vt�g�K�7dZV�+j�Պ�'��c��-�� �;�0��-��Q^^�
�97uhAۅ!��λ�;�ũ	�E�g���5�/���;{�1���ŋ0i�%=�`�9�͞k�Nڞ]�v��Jz"���>'v$��k�'nc+��k�!�%�|�Õ���\ۡIc�ޯ���eε]ZQ����+ʏe��kҴBr�r�K|��P��-(����ė�r�r��6�|����`<��N(��A^w���O�qm�뮋ќQ���~�E�I؍���]q��e�e��0�]���V[[�3�s6nX�D�ٰaV�^���NZ�\r�0�W?1Fj��~�~�jCUl�Aٍ��_�;Ϟ�#Cql�����)�xhcn�'b���D����<���`F�e�*�@�=^]|Ǔ�(2�iv-(H�ND��*3Pּ��!����Ms�
�~� �vm�!���Lp&�\��e��P7�޽�{;QT�Ï>U�� � "0�����'������.��"̞=Æ+���Ԍ�T݁�o��1z�2�*�:��L��џ9c����(-�EO� j ���P�V^���R��ʫ�J��^$4V��z9/$�ޮ�a#U�n[�nŕW^	�0�w�BL�!K튋�/T�ȝk{t�ZMS�������㺶�����i��XE�K׊�ݥ�*j]��b���zF�ޮ�J��8G-ĩ�kY|*q�:�{�J�a��Y\Z/��=�I�ߚP��먩;�]ݹ�$�[�K�\��U���+˽N�|��a'���.�\۵Ǌ�w����Wٯ5��]���ï�]v<����
)����IQH��ɣ�@�y���������4�������gƵ]9���89�HԵ]�&���ƍÂ���g�AgG'�ps뭷Zn�-�HcP���.���CN#,�]��*�y.d���	�9n�#�0�"iF�VT��GٸA!�/O��������F�$-�]8�ҿᡗ��@���Ad�����n��X�7��;,Ҍ���%�<ڳ�g�?���k`����^q�زe��SQY��>�Ճ� � �p��߇}$^x����?����;�<'-�����w�E�O<c,]ߡ�o���
��Xa�g�!?��-t���Ċ��H�B������hi��1k�
4̠�&M��P���4�ܔX#�.-�������@�&n���L!-�`�9Ƌ��,UѦc�C����f��V=]�!���\Oq�R��>A��'o��]+nW�6�sm���n3��{`�vy=bqZ!�	�0޳�r mw������|1�:De����]KC�����v׋�uu��@��v��܏!�4�i�u҈˕�b���դi��r���\ە��p�7u9��I�lJbwnI��ג�r�r9��S*G�Cp�vC>W��v���k|<AzPѺ��K����v^���4���n�Yumא	�vS7�f0N��Xu�U���^Xc�e�]�U�Va��#1�� ��l�O���{�Fvc���rC�W�#Ck�*
�P�>wu��*�� � B�3olJ(���xw�n|�wb��z$H�ND&Z��4}y.����"w��]5���;��GQZ��ӥ�k�������?����O��Cj@AD8\S�IS�ཷ�AwW�ps�wbɒ%X�tiF�s-l�W?Nu�!p���}�|��)c1��~[�����)�bYi%(i�F�X	�	�q؍{�A{� �E���=��X����v&8O2B�x��ٍ�����#�<"��p� nw�D�*�g�ε=&DU��
��yJ��zK�&���IF5�d>]��<�SsrfY(�m�vE��H��89M��f[���k��fH�خ���%j�����u��i�>�Vwa;p�r���A���>ism�21M�y�A96L��Rum׊����~KS�����c���C����+�,���.�7>�9�xM�8'&���n7ϼM5&��Jݳ��nh��0#}��n���S&��3���W^�����w���7ވ��:K� ��Ʀ�6f	gc'F���=ܠ鸷��EG���{�v�A;�Dh��6V�i��'������ � ��6���vf/-)�s�?���s`݋�������A�d��^t�����\�3�?�+l/*�o���H�_ȋ�S�ӑo}���֋�D�)�(���k�AA�ƺ��O=�(c��G�r�Jx���1V���ҙWN���?�zO��P�7����r�����E���Xv��m�%cu��������
��0���&TT$6Ġ3��5���D]2�H��F�d��*k��ݸ����E�?��= 3f��T���k���#�e�]�����Uŭ\���b{���x� W/KzF؊f�L2���+�Պ���W���o�m�vC�#�eҵ][^��k�sw�<�����vO��'������:�i���C�ε]�&����u򪳝&���Q���~����2�_���/Ɗ��>�c�P�Ѽ��)e�v�r�1푷t�s�RqmOPoh..��	�,4?�u��ƥ۵]7u�}��3Nǟ�����fn��&ˑa޼yy#<ϖ�]l�RNx�=�t�����z�8�����E�؝�t��1w���n�:bp�� � �P��/�:�1���ƿ�݂���ćD���i�)��٘g_�7���h<��C|������ ��3�����3,��P�Ct�	��7ƲӴ}�|?!�=��ܤ�/}���O�~��p˖- �MYY;�H:AAC��ң����z=��e�B�>��իq�9�8i���:?k�XV�~�g���;T�M����+�+�����mS,���Mh�F�X	�	�q�t��C�Z�R�Hh�*�3uapO��T�\��ǫS���a;w�n�k���X�]�P�傊���v^�TH.�n+}ե�� ѻf�.�N��m��(N�N��m�_G~�N�˭��zʢ]N�,e���x�m�nw?a����k�����B������lx1-{��B�|�߶u��A�EN]���Hu���3���$]ۅ�\�XT�|�
��.}�v>��])KSv"������Y�sm��A�;/4yl��b���!��m���k��@0��',mǩ�]��m�;0�/i��3��"��3f�?��_�a��A��q�%�XV����,���wi�V�Fl�5ܠ����1D�)�#ϓ�1W��"}C/r���d4oCu��vӐ�AD������j�߹�^|��>+e�ۍ��v����`B�E�&8����6⫿�]��b-A����}�CB���1���@ߡ�)����?/�}�٘��3���{�n�$��8���AQ�9K�<O=���+��v�mX�l:� ��0��X��D�o��w�>�s/B��X�����w�s�������� �;aq���65&��n-�5R�\	ۡ;щT�6Rś�o�P��?��x��@��I�L��E��A��1^d\�a�;5ǜ-����<E�nih���=Ĳ|^��;�IU���vN�n��B��M��qZ�v)����&�|�����ٹu�_e_T�3zlh�$-���\']�)I�����>�����)c���;���%��b����/�xݺ�ǉz�Y���9E��[�����Qʇv�@��bz��O��UwUH�َ��-��ڮM�^�
˵]'��s��8�?���o�DxY�~=֮]�o~��ƞ\7,%���26q��F-��
���*Sh����|�L�Rc��p�ݥƪ�'��!	� ����G���^������-8���h���_�Z������^�@��7��ݎN���V����%c��"Y�n����N7�����4�J&�\�oii���^j�N���/Y�#F�AA�ɈQ#���C��O[}D8a��]t���zTW����?�=c,Q�K֐��X�)V��H/p�0�b�@���
�㍽����:18�TE\#U�\���xRmJf�\ͯ�����p3�f0.Y�|�aTo�׵�O��!���&�Kл��BaE�n�[�4��J��L�T��@�rrf)}�^ +ocu��	�!��+ǀ��Ų��-�v�U2�P����h+1N�޵]\�%��y	U���F �"J=eq���,\2�ڮ�G�� t�'���S'S�K��������u��Bs������=���8q�N���M���_�v�N	���'4%�OqmWҌl������ �������DxY�f�.]�ٳgn�����D���rc��A�������"O��wc�VT��G[��p� � ���RQV��"�Z;�?��⢤���׏A]s{�;����f|��w��� ���|���h���T�c��j��=kj'p��<�����L���W^y%6n�"��}x��%3�AA6��cᡋ��g���&��lذ���;�����Z��	c,y~\c,��t�c1�����y���w�
Y���7�r��&������X<�-���8.n#U��*��ʷqJn���8��H��<�=��������A���c�`��I�}�(���9Ƌ��n�j='6S��U��q�A��:�3'���5\OjEܞ�k;�tS#Xw�)�]%q}]YA��pc��Nŵ�]uw���^H˵k�U��.ޏ�u�^s��G+l���따k;�oͱar_��BSGSS~����o���I�g�U�kFr���cM�;�E��=�d�e��<�h�9�+ŉ)���#o��ν���]�+yk��� "xum���C�8.ۮ�"�[qԑ�����>"�tvv��/�5�\���2+-^�O&�g�1K�?O��nP�ˍUѡ�}�u.��'��� �PAw�;Mm]��G'��,��v;򧳎���Mx��(D�z��[���� �L���{>v���
}�v?bQ���еܔ���L��|9��^��w�"܌?�LAA�IS�������2��r��7cٲe�;wn���0c���ÐF~��2�*v�
���c,��=f�U,c�l#c����ס3Q�v������C�Bwم���J<A�T�\;+d"� �T�=���^�e��X�|��%���7<�]�%ѩ��*��h����D\�U��	5S/����S�����j���[2��.�O�n��(˺	��,�k��jƅ��Hٵ]~K�g�:vE�}���Y��R�ĵ]WwC��Oݝd9��\+nW�+��>1�F2=b���v��5�����oH�k;���q��
�w���_�#l���C��h�Τk�����\U��W�ȼk�P3vĩ�]�R�Zk��D�Еk���m"�殯��L�m'���c>�)tv��ǟN֭[���'�|r���1K��3��*HW���+w^�n���5V�V9HA����bTU����׷�^z'�����I<�<����J"�~���ذu/
�����6����A�������k���X�;���n��eO�����퉎��3���u_����с�+WZ��Dx����}K�{A� � 
�i��DWg�~��G�+dzzz,c�իW����JK�+���cI��ee#Ic����ݚ�ѕ�����
�pO(AkSC ��"n�x]#�ށ�cx��❴��%�L��Lv��Hu�WP#U��<K�8�q��#������]���Sqm���=���!=�j9�n�b��vmc^#-���++h9�|��2G���z���(���R�'�ڮ�]#����ѻ*u��S�{h~7M=u�U��Ǹ��NH�@�c&]����Y��Ԥ%�ڮ�C�./h�Kε=&$�~�x�������R��si��)�A�������}�hlh��^>�����.]��'�B؞�2�Jb�i���<���L�o�*�L��+b�T��U:��&| � "d��c`��1����ڇ^)8q�́��%��;0����~�����R���C�+q[d�������ЊB�����_�B�v� 2JM����͊s{P������-&����/t�3�E���>B��7�x#�}�]�e���a��fa�R�A�@d���������p�~�z�y�8��R����|.�u��E��+��G~�`1a{��	ڣ�����hَ�����8�	�8��Б�{{�F�D\Dn�|�T2�dc�ڵk��*ĔW�c�'�@EeE�Xӄ�����ѩ��*�o[۪���T����TU����.
x�:z�]��b�?�sm�qL�+kF'\Y�OS�1���.�)u����k�f����[���-Kֵ=u��&�����;�V���1�Ƹ�t�!�/K��Z~|�v8y��v�Ÿ+���>�y�C��mq��[D�������ܥ����#l��+�j�s�\w��HU�_�Fx���]Y�D����.ot�?q�u,l��~q�l��]�ߓŴ�qn�j\T�{�i����|��Fᣱ��V���矯m�	[�S2��k�29�{"�U��]h�*r����|����^5o��*� �����|�q�A3����O�1���=�k���es��`���9�z���S1e찄��8z(n������n�(���{p������Ad�#&�讋���7�>���Xv����v��]���dK��}���n��&�e��i�oށ � b`3�������?N�1�a��)S��0]&W��ɩP,
7�3�|�?�}���Ϧ��9���XEE�M�lc�#&�1V�!�� f��R�46�<%�v��a�I�*?7��$t�����*İc���Q]]�g4�k�c"KU{(ƈ�T)6�k��CJ�햴j�ᬧ�W-'�k�R!hE��t[�.�BJO̵]���5qirm�Y����|����-FYAF�,ʽ>`h���d�j�f�������|�#���\ۍ� �?��j�Ǹ��NH�;���:i��/n�wm����(P�v'��Ƹu��]�#n����Sz��=��Jޚ8;6��rm7�8S�(����f�!V�k�5�V^^�o|�t���Oؽk7�����bŊ�TOk���^BwY�n7^ɍU	��G����:qsq'4� �PP\d��� ����������t����s��ĄM�=h|�������W_���D9`Z-V��E�����/�/�m�ی�Ͽ�� ��$̽��qK��Ŏ1V�3��ϾCO���gܽ]G����W]u�5�3Nj'����� � ��`��ֽ��;A����6\~��袋�}m�"l�d�d<c,Y���=S�c%���&2�
7$p�L*�k���s`���{;�He(U^0�*��r��#��T��r�J����l�?��e>r�o�i��&�dq�.9�Ft*���*Tw�̸���Yqm�V�R_)�]N�,����n7���c8�ʂ|�ZN��J����v�����0�:����'C���o�������'Pwq'��;�꤫���v�D��G�n]ۥ4�~X2�ڮ��-����������-L���@��v���$���/����	๪�/�CxT��	�v�\��k��K��:�v�hs��z�Ĕ��Y)	����TUU���9�^t1��@�v,���bȐ!����g�1˿��m��j����CT����{o/�^B�UD�2a�JK�-���&c��J�o��w<��{��Yh|������;��9h��Ə����]��r�g���,�eZ:�0��Њ/��F�����h�Ą�?r�t�����\q��o�/�}� rCԽ���	��q�X��X�s�"l<���M��ԇx���駟N�����-��}� � ��-z�G���"|<��x��q�1�d]�o~>c9#?'`���yW��)VPw���rq'c��B�ʂ�%hi�Gyy�{p�xQܞ�{���
j���X�T��Y&Wn��w�y��d�!�0v|�oLT�/����+�NI �um�3Ј[�<�Y	V//��Rw>�C�.�Vź��v!��v�صH�k��D]��
*�&��.�"Ĺ�u7��w��K���ڮ�ŭ;��h���Hڷqm�z	@�N��vy��5�cZSǴ���u
(���F���oajb��,�1���+uJµ]WwAH�QwUH��1�KjLJ��X/q{�8�е�[�ƙ)�A���k�s/96�:�L\v����	"\l޼k֬�w��]�F�|l�J�2�J���X���[�^�U�96��P�:#���I���XE�5O���>��
;��d6~z�
L�.�;b�4���[��f���?s���S��o�l���C��-3zX5���C^��m��76�v������ϗ,�z���'{A��;�B��Q׌�2&�����AD����{���X)����Q� v7%�ޞ���t�w�^�^�D8�\m��\RJ�� � DJ�J��#�����D�`��W\q-Zd��曉U�c%��n�)r�Xd�^�	j�2��%��0�:���*�{�,b��C/J��*_�t$�gCCV�Z"��7� L����|�"'#K<���p���Br>Nl�5�vM�Z�n�2�xq�R'U�kIU�FH�k�4/��d��٭WC%.��	q�&.ݮ�8�����O��ƚ��i��I�k����u���쥮ʊA�T�A�(��|��wf��?R�^vC�3"����n���F�����r�ܴ���a]/���"��RkYLyd~wOtxy�sd>�E�|K�����:��Յ����Չ�Ύ��N+N�}ma����7Y�vΑ\�7����k����|9v�&F�p\�5��@���k�V��#X�]�]ۣ��_�L��k~�X}D!�u:�
у
�����Ԏ�ӿ�-\u���y���z+V�X�9s�d�a)O�,��XŻ1��X%���t/�;���k�*nۆ��q���n#�0��+��y�w�����G!QY�c���N<�&���Ԏ�{~{��˛�~�.�AO��('9#�T��e��a�ܓGUEb�팦���bdGW��f~�Y��&���'-���͸��u 2Ϥ1CqǯN%w�	�O�\������"��=�v�з�Px�4�I%�����o�5�\�]��8����C�\���
1�`״ʊ����#�GG�g�[��/Bww7����Y�_�kA�GEe%�F���#��۶m�7܀s�9�IK�p*���d�e��ߓqq�ͱlc��'�$c��A�ȬQ%h��k5R�B ~�AU����ۓso�?a����=�XW_}5v��	"|L�1���㷟�"�Ћ���/:�c��G�v[L�&�bY7O��Z���]+��딄k�����Ă�����tû��]��J�ڵ=v\xם�QL%��++/ð�!�\��j+�4#7��0��g����hmnA��]hkk�&&�ʦM��أ�"U�5���
���<�G��¬�k���(vg"��Hݙ��n��o�p�&I�k;�����	ۥ�D\��"yE%m��q>�����B�8uW ��1N�Fx���n��d˵=V��T�q=���j���3�A���k�{��`�ҦϘ��N=���D�`��]v����:#�vdϖ^D�:ȍU@��*/w������ϭ����n;2tuva��"<�)��� �@iI1�;�8�ww��u���`�	��;�Ì	#����U?:KϾ
Da�?�L�ńQC|�>�p���i��ooC}s;�ʲ�Zn����:t����/��-8��	-�ne�x�g�������g�ԅl�g��5?>��� ����$�ִM�;}��bw/c,�_���h>C���X�\���ه�5��^����7���8�kj@D�(�\�BU� TE�V�~���43f?w�6����L�^QQ��.�0��?��\��B���	��2����c��e$���2tv1s��h��i����s�$3
imo��cvt��=���j���#�ӏ<F�X!���o����Ν�R�\������3��xc,��P��{�������cՂL��	� �մ���k��pq����f�wg�wo��d��6P%�Ho~>�5x���q�=��#ǌƼ�j��+�hĘ�5�1ѐ��\�*"��H�õ]�rBaW��;* ��cˈu��s�Z��<ëRV���p���u��f-�O�n���+��,ȧ��,8+$9����3���nW3���\���q�=���bjנ�(Byi9fΜi��Ʀ��>t��[C�n��c455��"�_KK�5���#F�@EI)fN��\���u�5p�76���YݟyA��ES��.��7{��=�@<Z��#�+Y���N�tm�
�u��g���+���=�v�pm��P�Ο������K�̵�>#��;�#M#n75q��=����>"\���+���{q�����)��v��J����� .�ȝwq�����]l�������B�1
}q��"l����Ɵ~_�Ƚ��?<�0�}��(�ܳ�9y�s��үn½��_qŰ�g����N��-ؼ�ac�Ա���'&��ۼ��n� ���ꆇ���??�Ȅ�-�l�?��%|�gk���p����G�ˑ}>�h� q��3��:��O2�]߃rf���z��}�Ŏ{{q���a�3��M*�b|��2�����^��'�S�`��������KDn`��Æ[��!CPlĞ�b�����1�x;Z�6`g�KH��9�����[H'���̱l���cƣzpuԔ��D`�^L�2v��5ԣ�'���D!2j�h,\�/=��p�^,Z�r%V�Ze����vI�a�&���X�wC2�R��l���X1s,f��tr1�(mlD�0&)Fk��ȉ�<���o��M�Нo������*z��n�bd�q)[�$2�=D0�D܁���=$�|���˘&<.�<�8Tc�1Q�~?��n������n�K������H��׈�=��Z!��E�(W��ӵ]���%.�k�X�O�\�_\��������u���/�_S��p�;�k;k|*��Q#��'�fo_�f�DC}=6���%`���F$���������%�c磡C�bܸq�6aJJ��@q$�Mm-���CgW�}�R���>+o�[�B�ߵ�s���]Zέ��c���iA��k���������v�sH���wu���r�6�+���83`�U�4��L�v7�[.�=���Ϣ�����e�5T-[��F�J�q�{~�]�SYƻn��"`c����m����,w�"K�9h5RIn����V,�P��P�QxT���柟���x7|�]����N���>3'�Jx���R�����8�o����Z]�;m���������>؎�0�v8n��)<�<�对�y"���Y��w������p���2��S����=M�w�
����8���ȝ�<���?�A��b�De�N���(#>{	�3���L�&�YT&_D�:�чx�-����>��;�&N A��]�ƌ�qc�b�0vl-F�n5�3{�޽عy+�m|+�:Vg�_��齵Cf����&��������"�Vl߹���"�L�g
Z"��;o���"�[��2�=���.\�7?��X:w^��cY.��X�n�1����=��E�ZD( �� �Q]託��i���\a{L�^\H�.7P�����T�¼��.r����p�޼[z�(/;(�x�Rum����
R�X�|;w�Z�-4VoNLmy~by.ݳ��v�Ny��.J�=ʉ�P�\�c[͐����T�e��C�>|E��+���*�[���j��N�H�غe�Y�&����������a���GCC�5�_��Ig���c�b�ĉ�0����7[�z�������h�
��O�.�=b�|c%�^B	����Y'.-��h���IU��q�ܒ��ӵ�TӴ���q�X/1�����vII^�C�-+%�z��vq�����I۝5 ���S�w�l��1��'��t�M8�s�������BjJ.�B�{���<��G��C:��In��%g��i(�)-)��sO�D��?�� ������g%$H�).Jn9"�a�'��V������~�V��~�5�{�����ב�Ԏ�;��Ը�^l�݈���NMk��2v7��s��F�
ۇ����4�v"Ӭ۰�=}I����Y��g쥦�,Q�1q�P����X�oj"���}���
� �ǲI��ljGyy�22���4�ﰘspWM�\q����k�����(�0�J��t�u�V�́S��}��A�ePe��P>nl-J"�(�oX��1�{o��?�[7o���L���^/MUF�]mm-�?E�%(++Eqi	v�ك�w���Ad����֖Vl�h�p�z�j~��3fL����3�e1ƲRݨ���(rf�Ż�k��Z��x�h<��D8 �� bTU��[R�  ���������;1�'!���
��*�|i�Je� y2��뮻���!��ߋ�/Cu�`!�4�{3���bL1������0X��U)+Kg˵�� �R����S{
۵Bx��g�@��m���-n�r�ܟѣ/a��g4ή�>�~wM1J��8Cg�7CSW�{P������1���Zמ��>455Zo*3q6�^؍>s|g�p�ԩ�>a2��ˬ����	{,������$�x��h�&/C���'^�r���浜WݵB�81N�FP���.	�}�؅��]�c��C�]�_#��=Z��\ot�ڄ�q�F�n��E�H {Y��o���~�A����G}4�̙S���t7V�.���i��<���,������Bf?����Á�#��j�"
&r���/��7?f��3̵������G��Os�;���چm8�w��_�W�̄�l�5y�_�/������A��}Ҙ�_���-��sw�y��wq�ooÍ?�rܗ#x�k"˰���<�����s�}X���~��y������Ww>ܞ?�&����c1��"�~��Q<��C�=F��Fgq��_�3�E�Zc��"!�˹�S��Y�yI:�~�N���l�&Sv:���k�J�p1r�h�_L#�D�6d(��2U���vv�hjl¶�[��Hw� �Pl�ƍ�dî�#G�Ĥ����}c�Z�[��Mhj�kAd������V���"<���c�ڵ8��s���8�g���3�3�]��>C&rgϙ�VaL�ޗ�1����Hmj@�� ������E��p�1��#���m��D�]i�R���L&����/�믿�r$���E1z��{V]�!��|k��Țk��'���=��)nW�ԉ]ˉΕ��X{%��1��!|��Tˉ�P\�v��ԕkz���q��C��������׵(--��1��)����ض�?��ըB䆶�6���[��`�x���iӬ�{J����Չ�;w����m��!n���1�.)�v���y�vM��(i9G�-	��k���ō���~��m��s���|S����jjj𭳾�?]xzzz@����^\q����+���vTHG#S���l������9��Sq���}V�V��s,���s�Qь�1𜙈�s4��iGb��1��GWw~��Q3��r�������ܖy�e"w<��&|�¿���91����-�A���3.�+6�ʯ�m�v&�N���ڄ��z�?ϼ�N��Z���S0�&�5���&��g\t���I���(-)��g���}Ƅ�x���y��ͱ�?{	��_;_��´�w�O��{�A�c��R�67����w�g/c,�+�|'��U�v�ȝ�?�bpS���&����^x>� �pQ=��,_f��A��oj�hL�0e�l��$����FKK����ߏݻw[����1y�d̛5Ǻ\���Y.�o�lj�����F{[�p��m�1�QG�y����a{`c,+I���Wߡ�gȄ{��X-��8p������� 	��ˋ���qtH�X�0a{��Jpp/vE���:��l����y!�e����۸뮻@��}���}fNw���x�ε]�_�!�+������8Y���S{
۵Bx�7���e�v7NW'���{�֥rM9ΐϴ��a�9��Hi�zj7CSW�# �kl���L7�G�B_o:�;��G���^!W�<�5f�رÚl�{��30a�8k��֎��pi�n|�@<��<m>�qK3�)O:��'N�nJi^������	�|�4��:�v�|I�Htn�I��M���N��EȞ	�v�t��c�&�פy��}�õ]}1�Ą��_����Dxx饗��C�3��LV��3�rRuq���ƪ�.{��#{��s\����ݘ1b:6��� :�z�����d��i�����X��ﭼ�7�B>p؁���~�F��媿=��y�����?��5JA<�;���[��<��L�����TL��s;��+�zDƺ�q�O����=�G?�w�ll�݈���/d�[�������}�r\}������uaoS�;����k�=s��MK~l�o{Ad��Euh�̰����,��H0ƒ'�(�C��-ˉ�4�ϣ�ϩ���2�gfzp��W�H0d���a�G���A�FyY9Ə�q��X�X����K���Kd���
�z�}�f��"�ע�Y#�E�%v����M��L�"%**+#����?AOw7�p�4�~����Bii�����v�vq���=�7S7ƚY�D�X!����'����q��*n�AQ@`;0�N
����J��bv��Jm��O�2����]Ԙ�#=���1�j1g�\�sb��O�l'��.d����ѵ=eq�R�]ۥ��]�iyC�fo61�D�\�c���乢h�Ȣk��um�����q�P=�
��ￏu/�L����w�^k�1bWѵ�4e2�뱧�N:5qCݿqm7�Ӈ�>8���Svm�-'��n9G�-	����n��g'm{�ܥMJ N���S�.��
��X_a;(nc�v�������?��c�{����,]�C�Q��KcU���2^�U�}��X�!r��w��y�b�^ϲΰ���}��6l��Nf"�����m�<�f�OK~��3�\�M��ȫ�XpOcn�}fM����G43�����Ǳ��W@>���>�q�]��/���D��E��y ��6#W0�/;�G�N)&�߲;�\��[��3�]�;��+�Ĥс�;�K�����	���ܻz���ǡ�8ywW����?=r�g��W�ӛ$+����,�+�Ғ��v� "��7�Mu�{��G�na�X^�v�y/]��:�Я�h���_�5�p���Ň/�F=%"q�14q�L�0��?lokǦ�>�3o�"�a�[�l�&���;̜���
�E�m�lh�T�M��!X��<��S��/���5"ӱ��p]���5Ʋ�⻸g�K�3l�ߍ�#��:z�8�!�� �,�+�l�K7R9U����w`��ۡi��5P�d۽=[Bwy�?��<�<9�����j�lIT��%��ϵ]C���r�JYYZ�Rng�>ub�1�%5�q��qm�S{
�5�
�vSZg'.K����)���Ҝ����Ԥi�G��Ѳ���j�?`��i۰����
���A.uuuسg�Ր���oc���<~J�ˬ�hˎ����Cs>���J�	%��D������g3n �<�+�N���qm�+��<h�z�ӥ��{�&TV]o݅@sΆk{B"�hj�8�4q��ݵ/
8�4qb�џ��oێ�^&_Xغu+n��f�y晁�����;'j�n��4X��Ѿ~ΑA�Pe5RI�ڍV-u;0a�4lm��*"�hh��q?�}��8�Ғgq��ӎY�/-? 7?�*n{t�۲���(���[��_��B,�*|NA	��o�'�>��I�Ł�C/�����]���D��>}����E\�����ډl�d����/[��T`�m��ч���-8��kq�/O����/���-{���3/����7��э�?:�e�w�����N�4���!���p���3����/�80my��Χ�[A�gVu3�{K���8}�n�a���^\�������ޮ#��0#�5k֐x)d�p>Fצgd�(0S���Lǐ��V���m���O�� ���A�{ ��a��sQSS���^��4����t���c������A���l�2:4+}��#l����z"]�aƍ��>C��ԥ����$p ,�T���nk(���TE������X��ޮ{�P����L�	���l�իW�%�%8��PZV�-��E�"���p]��r���)nWꔠk�RM�� ���[e)"xC��w��\��;+~�;�[w�K��}���DEy��3�e������o��Gz��(l��w�yǚ#G�Ĭٳ1�f0����������)�!��rm��Q�Ը|sm��\SVPq�sz��54�X?ز �I	�)�u�|�(n����15�X�%lW��ow3�v�D���W�c�v�ܾD8`�O}�S�g�}�.8�T#S���j�\ܹgC��J��VVC�Ƒ!޳�3���ЋEû����B�����߹�oX��6��kG�ƣ���{�51:#尉��Ճ��^'�	-m<sn�XSU���g�r���(�����Ҵ�[���߾�xr�F&6>��wc5sr�v̈́�?8q���!xw��k��G�𷮹�z��-��7�w�%2�E�wv����>��Ӄ"ϸL�<xP����1�>�R��a��J��ĄQCQ;���ʻ�w�'�>"y�y�?�7��D,�;-�2��U?<��l�m؎L�^���ooÚ�|9e7�Ic����)kjl���V4D�6F�����ȹ����{{���Սp����~��+�JQ��F��aՕ�>>"���Ze��n}�����>S����n��+<D����N_�6V�+�g��l_%�̪U���2��g�>S1���� 
v=_;�m�X��Ptuv������������Gcc#���K��Cuu5�O��A3�QVV�{va���8� ����~hjh��M�A���;w��o����='-_D���+�c�ֺ�W3ۛ{A�/ԫ[�������� �V�T\CbPq` <��*�l9&�;�D�a������0��=G��e�v��>�?.��>��Ғ��ݬ3��~Y��0R�z�<9�����}/!I=���ڮ[1�����-�.���cWX+l�f����Ų]]]�uo�"L�.)����::�#S��eu56Li�����푸��N456i�}ut���<�{��(U���*tF���Ǟ@kk�5��y�Ɖ\��;;ߖ���|&�@+����C���lڴ������g���Q��"`��=���҈�5�� ^ �9��ݳW���uo*)a�s��C\���aod}�[N��rP�4U�h؝v��:�w��W��kU��8I��mؽs�&;CyK�v�ruҍݡƱ���n�����P��f��u�׋���m�mعc��=M��Rj�m|����>r~�weu��=�ݩ���|�����.�����D�r_���*���K�.:2���~ˑ�s���o�'����n�VLEc'u���u��7^�`�%�7�&��W��X#"�l��{[q��wa{�zd|�]|뢻��G'�3�0��i���;{,A?{	�H�-O����_�q���;G���/���^�����o|��~��6�^�HC�+�)_�9"�,ށ���`~��;����8�vow>C��gR��t���O:�y�7p���C���C� =�2s�t�5��}���&lۼO<�8���+\�n����#L�<�Z���blߵ������%���Ԍ��F����oǧ?�i̜93�D��,vc,��3�Z<�m��Ld�8�+E{�����q���oq�F � @����l"�b�E�U�9�����ɓ<�嵝�Mlǉ�7��:�dK��%Q�����;)�"	6�$z�������������������������~�6dddH�SsaP��7��i�T���`soקUTT��w�U�m�Ѧ��7��|u�+`@�O�<	#G�BwWW��R��
ٰ���� `�b��=��x���4�V?�/>A��S}J��BX�ݝ�����ZZ)�[,Z�����L�m�p{�����޿9\�
=�g�G<����\�Mk���;��==��W�<��qIȘ�='���cİ������hn;وȮ��M|`e�]�]e�]>xv{��J�ng�,6b���Ŧ��kܩ��۞�F�b��{�{�Ɖ��یx)�bf���]�����{ݷ�C�
�Ƶ]H2VI���++�p�����F(_�@",�fnhi�����D�R����V߀"�HQ���c�
kwI�K�{�����X=.�\�v�l�`Sȭ�|��ʵ�|;�/e���G8t�V�^=�U<��U��*++�i��?���'�^�ąAKcϧ�E��2�ca�������?�<Z:C�}~�1��ŝ��<Al>|	��d�;B�{��?߄+����G��M���#K-mS������K��;�Ǜ�ת��_��7��5L.���������@�=��B뽛HMM�O!���)��1�"�/�:�C�7��#��D�Ň��ۣ���z&�c�>3��D���23��6�U>�K���@���i��1{&j+>�Kks3��o�X�3j�KDj�3�8Ю�;�:���@բ%��^���\�f�ύS�����!���TU��$�lև`�1v�u��Zo��7�`�6��	��:xP�������c�NKG���5wj�>O�`�5��,�N���v`�������v��Y���E��#v�c�FD}��u�~��������(d_�2Ɗ�1�1ݍκ
d�OBsW��">��}�S�ڈ. ��_��" M�.ua���}P�V�op�Hs�Н=��Q���v
.�,_�;0�d$��8K��|8k��� �=}��|����+n��r��,�0�Jd/�c���ra�I}t��i,U��)TT���1y���P6�ӡ����!��'�onh���_��s�ȏG8vE�&�I=��'o��n�l~aa M�/�&�_��%/nnΝ���5�Ǎ+�+%CV�~_����!5Սi�� {D�::p��yܺqӿ.�G������FӨQ�t�y�v��eÆ������?[�6�/¨�\�{�U��bbm� ����{ܭ���S����X"R7
�=a�h����{ow�:cŔ�ӂ����kZ&��pߵ�$Bt�;��\�'O��aÇ��	۵�Iru�i>��>}��qص]Q�G�Y>�[__�LfΞ�_����d��g6�>`~>k��e{"9�!��Z}g��^W������ݮw,vͳc��+V8���M)^RR���Na{<�U���U�"Xe%`�ڧ}.�C_�8 � |g�_}Ъ�
���	�`����~��h)�����b^��]����]A��4�E�/l=����[�c�_�|3�k���|��6����������)�q����������?�����ę��z�𱲰=u)��=Ԭ�����+�s�L���|��-b�S�9�ivo�s�N9r$&"�HaO��*�����Y�U��+V�%�J�7&/��1Ҙ���v�S�\��o�3:��m+����P�����f�x�{v-M_����p��p��ܺuK]�b�c�L�Z����Փ�]���<vv�c���gBܼ�<KF5M~M~~>�-Y���L�ܩ���e�pP���<+���卵���}�����x��H������fw�������~�����ٳ�ڵkcއ����c�}��5�ZSl�¡��}3%׍��{HOO�,P�.\�ʢs{�E�����x�����?u�v��"9����V��KD�$x�߾�,�N.�@'��ۥ��F��¥�yė	���/'���g"��'Bw@�:ydR?S!�XM����ן�r����̵�@\9j},�ݟO1�i�v~/�Ǹ�QܮK����׎�<�|���aʄI��6�Ο;�{�� �E[[~�sj�����%KT�{cK��b!� ]K�?�e�t���	��l_��<|5��>!]��b�(���ZYKE��mR������ }� ��R�:�|���˷�5��'{5���p���9y��p�6mڄ'�|�A�x�xB��߷D�.wrOᖠ��������
���V,��j���nBvÞ�m<�se����z
����I4�?��?��wPy�	!�������o�u�D"w&����D���w���������r�����o<���n$���|�����~�|���1�8r����p��A�G�n�2um9�f�e0ƒ��M�!͇�[|$ʽ=V��v�&��/�& bu���[��U>+W["aQ�2�u��zI��#$���~��.�ʷ����gW�Lp��x��<�S'MƤ�	�xO׮����#�uf.�j�69��so�Lv;�=��*_+;��X�����'�ϓ&M§�[�=�
�ߺ�[��b�y����z{]��[;�L�[�qE�1g�|��gh�;���cg�v�mV>��i�ʕ�0��6�pqW{%}�2c,S�{�����p)c��	/$	�1Kr;�Q�2��F��U����(^\�}�,X��`0�������_���)av]�X���=^�.��+d�v�ې-��D�.#�w��K%(l��[�����w�K2�ORw%�h�C����=$u�	���g��X<N�d����  27v�P�_�Ż�K�򐺶����4����V�o.�d��۝����dg�NMvl�F�."�0���W?��՜y��FyU��t�����=�h�!F�Ǘ'�hݲ >xK0䉗k�T�-y��򅯿���Y ��(�"��v�9QM����#����$Ͳ���|B|��}��O�j�-/E�W��uTWV�����a��^x=��:��l}"�L��Od�I�U�����?�`pq��|n���.�����_�-y$"8z��������Q|~�\V��������v����Dh��?���Ϟ�>���	���o���Q�P�W�����?���4�w�Z�[5xy�)$�^���o~�׫��g3��Z?xq'��	��7����1V3,��3�
�o(�;D�������m�x����a�\�~Dr0y�4L�91Ta��.�3i�Qv{w&f@(1�a3���+L�6�^���N��p� ���̹�hlh@��� ��ŋ�q�F<��S�	��K�/d�;;��jB*��1�!�� eTf
��k�#n��� �G̘�ۍ��@�&���c鼠O۱c�?��T�>��(AΨQ&k���˅����ɒ�z�]�}�v�>��Y*l7��Lx-�����˅�<֮����ȵ]��c�n���o�h�PE�������yy(�/ �B=}�::� ���b���ôIS�k���rQ��	>��	��[��\L��[1���<���ۏU�v-�����i�x���.�g�K��&�NH�,l����k;���w� ?���S�Φ��o�����`���&�K�����U|�*(r7��vj_�ߍ�O�
�����[��1o�h|\K�*"9hn��w~��N^ŏ��2��s������?{{O�<��u�����`"�dvr�����]TЬ	c���hn��s�K����g���'��6��k�jr���tu��/�{3��sA8���;�0�sHc,S�w�s;����Pt��xϭ�%��QWW��^{Dr02'�K�� �"ƍ��������chooA$�<�VvM]2331���\^U�+���>�	b�����u�hnj�l�����ǃ>��}K����l����ylJ���1�n�A�A�����y��v��/H�O/�2P�|�*�ta�qB�)�y����n��W����$aڬ�4m�����v�0�DH.1�5�]ShJdA��
�QP䬭��(_"0����v�A�:*�D]:'l��R���k�"pmαx�=�}��v]�>�6T���O��|*b�ظ�+���q�����=}���ܼv���{�X����`KAA,Z���lܮ�@k[�(v�a>{|y���a�(�H.O<]������D߶�1Z�vA�Ο-Ͳk;�|jJT�L�,����	�%?#�N�Y>+�v����B|�k_�+/�����7��g?�Y�?~H����b���`PJ�˝�mOc�*���

�-�����#��qm:"�xs�9��^�_���1k�v��?��P�L�D�|p������X�����a��2�e牫���_������7��BZ*�JI���q��m<�?�_��Ӹo�$7�����ĥ[w@�3XR�Fks�32C
�������f��r��;L1��}�@P�.�/.�i�!t�v?�楗^B}}=�ÌWV�_����P!;+��C�;W>��}��� �BGG�9�~�0q"�_�=}�8s�<ZZ[ACw��k�`����%C�SSS��_�>�lT}x���hc,���P�7�"�9�A��A�;p�Vy�#��]��)e*>0%����E�8/�$K��~�|�M\�v��ۓ���QX�l�dM���r���AA��7�k���}��� '�����k	um��G�W�O(���µ]���=��A\����K��z������)���҂㇏����L�F`Ͷ�sa鲥�5u:�5֋�6?X�D�)
�%e� ި��%̵]"��$�GV鶰,ngI����xq{��5b�<�|��Ua���*�KKp����!gÞ�/������>�6�]��*5Ű^�T�)X��S�ۺno����}�����Mk��Fa�4T�� Z,��6��)�5Y{/n�H�ؑ�Ă��s��o=�ov9RB\�N�9!��˻��&�C����/����O��>��z`<~��G	-���ǎ2OwOZm��%& ��^�o����礶�u���K���������z|���Iq��t����>H���`�N�uQN#�05��ݩ����b&x7�����'�'����vh1c��dro�~nܸ�6�H��Z���`�ݧgϘ�����؈c�F~�dn���Kzz:.^�ޯ+k�q��U2u#=#G�`��R=p��y��W�裏���hH���TQ���fc,���e�X�d��@H�>Y=х��.�[��s�\���b0E�/�k�!����8-��}3����_~�^�� &�\�~�:�'z�vN�n��X������]�k�v��vH*܁�8\����ܲ�]1�ת�=P'����!�G�O�D��mM>�յ]~q{aA�

��vl݆��~D2�\ݏ>�~�>cF���Ģ	�]Yaȗ�v��[�{ty�u��k;�ñt��pm���F1:�SX��)䋽�]�ϣ������k��n]�n�����O����(���|��x�'0o�<
V!x�V���ԃb�UZ�S���Yrd`"�^%�c{�^�Y��Ld���u�[4�4��C�wb(���oC��w���M�Z��l?	;�����=�o�;����()��d�����:�����@����ϣ������=�4"���:��O�E�c�����?|���ͦ������C��d����_���S
s��l@�W��5[��濼���^����O�pt��م�7��K1�-'0"3]�j��kUu��ߢ�N�R4�����:��D�.��ٞ�����`<Ÿ(��+O2��t?���/U�ٴ�4�f��b���<�.���|��6?��ΜA$]]]W��EEx`�Z4�����b03a�$ܭ���+4K��ь����!�F�X�c�rm����1��d��$H�>��C��< ҉A7͠��H�Sf�*��bD�-�>�c���o~�ܽ{��)�o���K�޵][��+� �tm�nle�vU�l&����	�?.�G�.
�9=#45�Dr'�v1ݪ�=&��|�$_�\۹�R_S0}�4�de���r�ܶ1)�z7o���#ǰd�Rd������T��C��M���=.��ϣ�)��x��C�fq[X�C�̊�k{0yyѹ/M<��	�}k�x4���{��v]u�y��R������_~���N΅M�����?��e�y������PdmH^�\R�a���`�*��B��j�F�{:i�NU<�������KX�`�asm��;�۽g��p������b�K���{�ǌ4�?r����7��i�t�Ld��߼�GJf�ϾxM��D�|t���>U�K����. #͍����w���k����u[�����g����ϞT���0����Vձ|(Q^ۨ�K����0oJA ���_�����8���o��?�����gJg�I\.��>7�_wƹ,�g����{N��G�Y,�UdX��<���l����p6%���'o'�֋���jz�i���M�o�m;}_a�vk"����ɓ'�k�.�'wL�.^���>�������p��1455� �꒕��qc�b��8y�4��i�#bp��d��Յp6�1����#�#c��c�u3?��?�(XQЇ�i��� �� c��T�46 #C��.�XCM3ȋ� �T�.� ,z�*j�e`���
o��&�3�x6
��Ңwm7���K��ǵ]"U���%K�Q��x~d�҂Չwm���XL���r�JrC>�$� ��1�k��p�`u<�܆Ӯ݃}�X�~��b�������xu5b(��mߺM\���"gTʫ*����� ���O�	�=b��\m���u�z���D�����DD��n.l7�v��HωGH�.�I�eq�\@�������/�$�uq����qEޘ<|�_���
��9p� �9��+W�&H�?Xe���`���tc�
)\�t�f"w5�D����������`��/��U|���X<�	�\�U�7v��E�����N^��k�{��xd�����������32b����j�$A���{����U�a� ��o��U�e�{�syy�)ܪm��|6#GY�=|��E�9u�m���E��\��
s���^��}�0f$��:�ܦc�r�Y�%u����}S�/�5N���/n;��^z��l������X�h�.����3Pq�I���(�<��+�j�T�Z5�2�ۃ}�b�a�i[NH�ԉtmV�dro��_�}��/~��>�w:���\w���&��F��ј;c6z��������AFZZZPq�G��E��3z�^��w� �}�t��޴�g�F8�x�����rc��˥cU!�=]�C��)	 �� c����Xwo7��SR$��������|K����N4YM�~^z�%��(PǓ�;
�hѹ����6�]���N�-����u���ks�vQ�������-���H�G�W�Z��0ߨ�ET���C�1�c�iV]ۇefbެb4����ӧ��:��B��v�ڥN�[��ESǣ�n-Ztׄx?���C�֍�v�N���˵]�BrѺUq;$�,�k���|J�]�%�: a�o��ඞOvB��E����a�iy.^�Uk����πp.����_�%%%��@KJ�*�o�d"r7wc3ݠ_�n�B(`ev�x������o��T�GwO^�}F]�Ρ�ԅ �2�_R"4�n���^�"��O/%���֣��1t`��{O_S�������GjF�Խ=lߡˬ�P��l�2/P�C�W�fǾw�ޭ:��g٪Rd�A&F��C��Gc}�ۏ��~�P���8zT}�3w�ŵ[7p��M�`aD����
� ��9x� >�U�V���7T��y9��[3ƚ���7h0�S �� b�pZ�j���jY��r��Tza��yAV�[ě��D��֡����>g�DF+֮Q��d$�k�o��k;?�D�{�]�a.��"�%q�dP�~[E��>M,'�$7��H�I]��O����q�u������?{�[۰w�nܼy'NAu��ȁ��#˖-��)�PU[���V㵪��nE�܊ܵ]E7Ї�[��ĵ]��>�F�4I.�̵���c|\�u}Zt�L�,���z�ָ��|��y�~�ш��|�I\�Z�� ��޻w/z�!�Jv��I\��X����*ƀ�&r�̑������T59�AA1xpy�Ri�����.��=Tߡ�oȷ����<�����;���/�v�~f�-f}&�d��o�͞������7�Į�4ؕ��g���/�˴�����5�t����&`ʌi�WC�8��������$�˴}��G�ͮ�� �	���}�S"
R�������W��漠wn������[|8!��H��鼜ϒ%���������ȥ��rm���B�(c����9ѵ"��SXBx� �Ӌ�����C����E�\^�0^�gb\�e�T���GH��ڞ���y3g�|�w�:�� ��>~�8N�8��K�B���*�wt��:�^)T����1�Qt1�E�0qm�vF!n��%sm%nx>���vs�QU^��[#6�����G!X7�g��r��`>�ݽ���^��^����տ#��x�;t����0�3M\����*N9�k��{۵��SY�Ϯ~�������a-8�AAA��w�������0�?��v��0�k;'n7.|�=H���E��-[���ŋ �ͨѹ��x!b00s�L�8	�=��'O���999 �VV�.��������nC>����D�d>ܾ���ΩS����I��`c,���ڌ�8[C�XN�����n��~����.h�(.� Y�
�EA$8A�m�>��c��A�����)��%!����/�Doѵ]-�#�{���n���ź+�W�*�	�e�p�w]��z��IZl]ە@5![ˉ�e�7�l<}-��RQ<s6��{���>BGG�{V�:y
gϜ����0{��WU���w)�\�RخO�u�zL\۹�,l�p���񣜴��]����g�fY�.�g"���w���[�G/��1|8��������\.]���[����=��}�i�! lS��I���c�����t������g6ژ�Sp���d&� � bp0!�m.�i��l0�6�8`��O���Y"n7������4M����/��2g�Nu��U�o� ����&cƔi�x�cl;�A�S]U�.�&M§�[����q��5D����'���}}} ��/�K�[�iii�w2Ʋn�%ӷFl�%���c�ц�Ha?$p$����܉�����9q�4��P������'	�����_��4Έ�l,)-7�W���3qQ���xѷB���e�vY�|Zl�b{M�m�k@$��ω��t��Z�;׵]�}b\�� w'T���O�wc��Ӯx_�\�3s�S�8|����AD�F��#Gq��	u
�YS��Bw�,�iq��h]�`-�?�"y��ۚ��%�)׻��uH�Y�vm�ϱ��{�v}]%k,�5y��XK\�z>��	Ο9¹0��~Xm�1�┐��oo�5��U27��x�_h���v�Q�J��µ�Y�mE��@AA��d���p��i>��C,�}�f��C���ͱ�&Q�Yy6l��7@8�ťˑ���HV�L���i3p���ؾe+��έ[��eʔ)����e�v���Dr�������� �KYY�j���㏇�_\}��1�2�il �X|���n5F���v2Ʋ�ƻ�aѵ]V�B	��`�4���=�/@�n�<NO�~�;�����p.�w�b�j��o�:Y�N{lUH���%����[��[�R��.VS�򺛊��:���a]Hn&n7�cE�����˄��r�JrC>�$_D��2��(Z��#�9��P��Aa���;�\ձ��#h�i�"&0���C���ѫV����B�WV��G���!^ky�|f��X����B�"�ܵ�w�t�k;�ٶ��'V��r�
�#�+}7auI����eܺq�M� �	����{�җ�dk��,-^��xQ�)>�_� sd���)��z��̉0l��.e,�<!/j� � � �S:��u)����Rhq�Q<R�-��3�Pt��d1��Eymmmx����E�2i�L�:��L�03&Oŭ7�e�f1p؀4�L�6�{ ��]Ey�mD�1m�L�Vՠ�v��y�2Ɗ�1�|�2�"i7�����6�d�C�A��l7Z�� =ݚ{�!H�2�1�"���휸ݸ���I�x��g��N8���`T��w��V�ߘ��Z�+~��k���~�:���V�����u@�/���ta�T/
�4q� WO���;�x��i�X'	sm��! nl8���S�"od:��&{����o�>�U:֭_��a����Њ@�.�!(n�%�H\�%w]i�"ӗF(n7�y��C^+�v���{����ػ���)j������Z"�2|�|�o�����p&�~U���琕�H�;X�� V����Bw�w1h%�nP��q��.��A�r�{WW'J�Rq�6��EAAD��N����:ҙ� m���L�Yt��`"�El3�8��*V�������\�g���� �d�pl��*��7�k�;�_��.�s�����ŏq��]D2�l�
��`3:�;@8���r�����l���<-^���1�g�1VjG���)�		�%��誋̹]&n7��%�Ԃ0�ۍ��z������}����	���Ɍ��Ys��u�:��ت�\�E/J���<f�v~[_�@\�%�A��ZZwSq;_��\���k}�`5ż��Q��,D�lh(�|>�x���|@��O�0����[P�����3q��y�<tAğ��.�ؾ�F�ªի��׃�u�L��V��rm�܈���vA`nL���o���G&l�t��@d�v���E���s����1pm�y0m��}`=>ܳ�3�s��z�-<��3�V�`���]��Tƴ�jS(`��x7��`� � � �����i�c��D����B���?T��!�W�XųOO��Z������p.췺|�
�SI>A$ÆÊ%��\߀��w�G.]��O.}���c���8x�:;A$l���W�Ý{@8���G%c�c����l�_��ڱt��*{@��В�TՅ�ֲ�B -���l��pn������ro�W��`�u�|�
��OO�]�%Jt��\gYl���ĵ��R"�6�K���(:M�nȫ*7��3{A�D��.w�W�k��>�O�������뵥���_\��������to!hhh��M�0s�,,^���5hmkU�yL�Ӳ����KH�k��B>�Ԕ��p�vm���Ks7vc�Y]��!B�ɵ=�5������K�����3aS��_@vv��ݩ������f"w��]�� �vPk��E�j��E���h�AAAD22Vi@��m�Kߎ��w(k�	�7�6|�a<S3�ЯhV/�oXWW¹̞7y�� �d��w�.X�w:�݇�]D"`��sgϩB�e%���=u��� ��_X��g��+ ��ݻw���o�w�w(*��XVL��n7&�5�2A�	ܓ�U��ֹ0D�&�/�J���T����*�o2�%�.Nvo߳gN�>¹L�9Y�Y�f�/4�q���\�e"k-�~[3q��]�C��T�.�I.���Wz> ��µ]Z��v1��'k��>���n���F2�����;s�eN�A�˕˗q�����b���v�8V���(<7�G#n�l+Л	֣qmW˒
�c��$�ĵ]��Do�	������=��<nw*���o�?�	X
��f��drq�E�^į'��4��V2'��������X�xi^*�@AA�tL�q���Խ�l௹1��H ��d��0��3��8�o0Z���ذa�=r$��A$3�M��	�q��a՜� ����ݍCDNN\�5U�t�DÄ�Y�t1��Ԣ��:@��믿�'�|R��0�+�1��g7c��ZfMCuc�	ܓ�|ԣ�saH1	T�#T\:q{�i��(���`Uh�����h�ÄC̅�p.�y�QP4� ����L\T%��������PBtױ:y�-e���g��.y[�K���=$�vUyi�k�c������Q$e��L]�����8���]۵X򔉓0nl�:�zru!G���G���ӧ�z�dd�����>��$6�C��s�`�_ [�=K�"��+FQ} �xێ�k;W� n��.�Lخ�9��c0�#�=A��f{��������#��,�n��)ʟz�!�
&�ި$"wM�n�������w��.���B������
�)��C�B� � �H2���A���{�m$�K�7��"w��1�P�k�����HD�T�oy��E��d���a�칸^V�m[�� �ill���;0i�$<��~��p��o�p0��d�J�ٲ���
sq�w�ˏUc,m�gK�X)�����,ۇZ@�	ܓ�i�n47�I]Rn���ǻ��+����]��!
�<g�b������̙3 �Izz:f�-&h�A3gT^T(|�BA_^��:�/kБщ۹􁺶+!�n*n��k;$�C��k����;/�O�k�$���0��Fdaa�\\�pg�� A΅ͪ�g�n���㾵kQ�Ԁ����z����v.ђh[����bw��&l����Bt�$-�7&�v]f��ٶ����ۍ�ʵ]�j1�髩ٻ���t�o<� .�?��@8�z��w�j��ؤ�׮}[3�+�̍��R���lf�~��u�>�#�q�3q�xWW'V��ay/� � � ��47��X%�q�L��3B�ۃ}����Pm2��ݸc�z��_���{��{��)�4#Ff� �Jff&�/\���&�ٹ+�ށ ��s��-���c��%X<w=�ήN�������sq��y΄���O��Xc�I]�����-���S
�K�Bl��I���Nt��S))a�U)~��@�ʕ�]����S��� ��;�`��?���Ԩt0KV� --��/�Z͊k��R����Pΰ^'l��[J�إ�v��Zs�5�K���=$�QW����!��M�����.�'=0���E�v��.��M~J`|>��9�̜�t�[u]�룩m"Y�s�6��6,X��g�V�mt�#�ik��"�<!���$ك@���|>����O�k{�"x��v��]ۣ�`]���]�r�M���vr���?�Ia�����\����[����??Do/	v�V=������V��`����Py�˰�RGp�^��9��J��>� � � �H�Lp���7`����,�Cti���>�C,I!�@�7��b.�X��D���|��7ɽ�����#���T�[���G��G���� �{�:qX�z���Å˟� ���VU���=΃c���{�ַ�R{��$W�`�4Q���1�oq���f�}!���~Cf�UZ��A2Ʋ�')�.ݍ��\D�vލA�j0d��T�P8I�� so?u�gR4y"�O�����������8�Y�v���,�Nt.�˫$<�<��O�ĵ]�ˏSVnT��]w�ssFaެb=rwjkADrr��9\�z>��:ۍ+-��KEےm�qm��Fat4�u�>�m�yC
�u����#I�ۍ�v~�yyc���㽷��<�`����o~s����Py�#MB�2�����.�v�>M�������i�i�!AAA����:t�ܦ3>��~�3>���Ӻ��j��a�C���q�0=�fXx뭷@8���T�ܷ���������ƪe%�p�<�ܦ�	"�������{0�����!:y�m� '��뗭^�]����Cy���Uw2Ɗ�K0�һ�{ۿ}C,��V�o�FaJ��>4���=IY]�BoS�%�k]���]?� ��`U�nħR��Ty<�4`�.�3IKO�⒒`�U* ���M\�Ec֠��߫�=�ϸ�����E��Z*����a�Bµݰ_]����qzd�$�#6��&�u�\π\�ŀW�+����s��m�n��G"b`ttt`�ƍ�2u*�F�Fzj:�{����8½]M�=Q�n*l�P��/D��<�1"�)n�۵=Z(�{�哽���!B�,X�@oR�uq���V�Y�sg��z�5΃�łUYY�����|N	8E�&��h�Sd�`pJ��td`���Y�J�^hlG��htn5� � � ��L�FksC���%�+��{x3,��v�;��%}����TN�ӋW����F���e���6|8	�	G���-FzJ*vl݆��~��TVT���
�J�ctv��8�pY�٘�p>Ο:�y�1V`MXc,��P6��K����#���f��-�P�5�-�~�hH����)��\t#HB�0�����]t`����k�!�����i��4zک,)]���t�Z���Ep����µݤ���U�D,:L^��\ص������j�H��:�H�ڎ`Q!��Qsc��Zrm���--�/���Sp`�~
p� ���U���by�r������ڿf��*Ҥ�	s�(���=��`ސ�v]Fö�|�\ۅ<�|\���!M��״�S:�N��t����em�/~�+�ɿ���4���`S���;�`U��ݭ��/��LD��E�� ��@�"���y<-5p)c����AAA$�Ey=�g>�W�w(k3�	d���c��oێ<ɘf����6l �L��b��� '1&w4�-\�ǎ�qB� �6H�ؑ�HOOǂ9s�����M8��s�QUQ��;��t"d���	o�e���h�H��3��O�n��?@|�~lj�`H���f�F�\$��.��L(`X�
�E�􁪡����1�vr_v&�E�1a�$�D�m��-lε:��a���Q����e4��Ʋ͎3>���9�����^ʱ���+͐&�� z�v.��v��d�"�VW���A^X�j��m�0aV�^��;5�û�ޮ&��۵�5|��\�u�yq����`����K�2�����p!%��>i^�X�\p?fL>���`��A8�z��1b���@�N���G�~!�o+�wi��_*�0����}yu3��׳�d�KŉJBAA�sq� }M5 ��@^i[�\��"�4��v�g	N��3K���o�[��׃p.�O����=�t�2�vucۖ��9 �AHCC*++�?���g��#���A�{o_��;7mE?�&��\ܿ�o$M_aB�� mT�K�Whj$�kO��ZZk�w��>��0H���,ۏ޺`'��T���2�v+.�`�4P5t\��:�cǎ�p�iiX��DP{��jɵ=�?�vA�.���9��*���@!\�����|V]�5q����$�XssFa鼅�p�>Q�JĠ���ۨz�m���~�����j�\��4�ʟf�G.X7������d�3��vq[�$-(n7B���=Ξ9�۷�A8�z����կ~5�A��m +�����q;�'
1|�b�Jtd���'N�h�	d� � � ©,����.ddd�S���?�c���!���5��,-N�k477��7��L�/Y�~L�����q(�>GFKف�`��+�>u���XW�
e�7Q^qa7Y#�Q�`.�>�y���+��;c!l�ahc,En��}���%���XT����= 	ܓw�x�iLSڈ�8�0���]�o�A#���e6,ӐpI�r~�*e��k�O�΋��ڮ+Ǫ�]�wK���vC�%�z�8]�����D&�W�k;L�)����^[<}�\���۶� ��saؽkƏ�5k�Cyu%����qmW��{9����&���u�d[k�v-_���H��d�3HO(�ľ�Ƶ�b^]��|L����~��Sg �k_|�_P�-e8�Q!�i�����~4���M9h\�-��R(k?Tz1��sk]-FeNAC]+AAA8�"w3��n���C����X��?�T��� ��&����<�DRg��ΜZ	�;&�f� A���.�3�2ұs�1t`���ڍ�`M�J:~��iۙ5�U��PG392�
|���g�e�m̷���i��pi 	ܓ�Ņ�hom�0H:��S��ȅA�Qsw��c�v��y|��G �G��BL�:9�]�K�r~tB�D��C���k�(����I^@�ڮ��k��H�ٍi�pmgI#G�`��blݲ�UU���AC6��;oo��~}#�q��^��dQܮ�	�O�����>�u+��y*l�ok͍�j��`4��������jM��ྠ� ��ضygQQQ�-�w�'�x���Ĥ��h�� �'D[5���2���I�*%��r��������~AAA�cTf
Z�� 5-U:����p����]Z�~@�﫾������+���6l �<�o�d�J�~�����\̘0�.\Tg$bhr��9dee�����3�[wa���ؽi�p l ��6�R��=c,��=�1���0\���;lk����h�r΀���1'lH{�K:B$N�\��`�n��M���qo'��������R�tWn�@2����9 ��ӄ�~Kq�_�pI|9F��_"l*�/W�2Z�v�X_f�8=jrt���O�|�E�R�����wmg�3�NG����y�F5�M������͛1w�<u�YQX��"O�˺G�g&l��k���$Ͳ�]k������Ͽ7�y��}0����{�~�>y�5� ��k����{,���@R����wQ�z1�PfV�vw׋܍�7��2גAAA8����z��Zǻ�)��1�����=�)����x�l����x�}���s��1g�|���A���������<r�H1tiii���[Q��S&NƱ�'@v12'�����s�p�o��V����<�۷g�1�L��c��f��z�;?���=V�K��} 	ܓ��i
�j�v>H%��i�1`&8�waЂUZ$J��ȅ!NRݸq����)������;UF��/W�{5������ⶮ�N���:���!h�f=�bf!U�s����y��+G�)���Z���e����._ՕI����ȮI�n�z�xKs�wi���2nb{}}����㧡�W/^
d�����K6f`B�����~q�:����W}�ioo��z���]S�655��͛����ݭ7���soױ3�<�������.v`米�\kk�z���k�NL�6]��o�D��5hjl�_T|X����D�ht޾U����o��ʵ} u��>盽Ϛ���ЋDD��[����}�;���7�:Uܾ�=�F���9s��Ҋha���h�5?��o�����~<��pjp)�4� ~Ќ�;��.f�
R����Li-��5&����	� � � � ��.�Y�!o�e���o��4��v�_����x��> row&#G�`Ɯ� �����}�+��s����+#bh��GAaa!Y� =����/����媶�p���:}�Q2Ɗ��0��d�g�Qf>����gZ��(H��D�,r��ރ�4y�{��z��=���sa��D��7��8L��a㋩ݎ��*?'w�.���M�\�����ѣ%��&��H\ۅ-}�n^)Ô�Ӎ�T�b�������#pm�'2q��Y3��HC'|}$N�fy�\�YBխ��?��c��L��zB�O�||�Z�¥���'_��9s��]���s�k{Ѹ��_�}{� 77W]L��Į�������rL�8v����'O�����F�ߜ{\W�<v�˿{�.�6��`���c���SũEEEa�vz�V�Z���
p��RM�ֵ���S�9{&��Ͻ��EwwF���L�~��uƆgĮ��Me�~Y��	�++*1�!_"\ۙ�}��حmm��;p���{�y��ڈ�����:~�(���۲����q`��߾�꫸���uלSI�[��K�78����N����b"��E�����Ơ�j�������t���AAA8���n��4###Cp�sE�w��l��uq{����B�	��X�m߾������v'ۇ]��4��Gf��0q"ʯݐ�okiEKSܩ��&��1�5[�fq����4��<�D�?zT.��x���͵��K�m644��4��|�g�4v�i��~����3�rV�]�;���ifx��Xݎ;�>��[[P����P������T�]���R~2��	�'��{S$��;����<�8��6�����
8p �ׯ����d�e����3���&�Ҳ�Қ�1-w4�Փ1V" �{1������;1��L��N����O��6m�,�osɊU�.<��d���L@&s{���ԯ3���	*�%�Ac<�t+��>5�Dh*$�i"n7��s� :���Mq���Vw�7a��?��瓈��`1�1��Iqa��E�}�&v��$��{�9t�*�_}�ܮ�R�\$�,EģO3�{�/���Wo1M,#�1��ݷƚ�=�|V�޺�<o��V�������{���p��y�f!�9sFh���:&�{�4�����KQ�>h%�vP��nɍA��94�4V#5e<z��AAA���Dg�[�p��
S�s��� �1�T������3;�Jc��z�~�8C�8��n��=^�O�5��3]_[Y������D�Dg�gL��l6�5����h�-��y�(��{W.]��ڻ�t�����3���ȑ�8es&�����V�ف������9ոq�l)����.��ܳ���3fL���w��K�b��I�{��*���~�3�d�!6��$�g3?�߸U��>�w���<���~��P��c����+�`ݺ�ɜ��
�j��ۧ����PhCs�� ���ݸVO�X���I¤Qn�6�#==���nű�X�F�D&n�[=��������r�3y�<Nx���)�=q�\�9�z��X�D`�龅]*�D���bLԥs�v��㔉����cހ�\vi��ۅ㑉�}*���2M�|�Q�"x��S�-��m.�8x@��G�K�9�,���{<�Au�����~m]hni�-���
u��N���h]ۥi����NQ}�U�j�/��v �jM�n�������ǟ~o����~+l�(&pק%C�i�if��N���v~@w�@�U7���N����AAA�M�KAwc�|��žC3w�8@�_���~5�L�-���E��δ������� �EFf&�-Y�H4cF�a���8��C�g�$"����eTUV����ȩhhjA$��%KQ[U��8B8�ӧO�ĉX�|�c��`�e6[Y8��@{��kzݾ�Z���y�?10H��$,݋�:]P*Dp�J��̉!.�$D�JcS'���{ �R�_��Dܮ`K~�qrm��A|-�[��Na-���]����]�%�Y^��H�k�pm�y�ߍ�vݱI��Ӯ��� �ǍǖM�b2z� ��s������j�j�E��Z�z���%I���桄�j�GL���2���ֈ�h���Cɵ=��k�(/]��G��ڕ� �Ç~��/bΜ9Ip�E�Q�΋��-fA*��g�C��f�AAA�ݬ.b3M��΀�����͍���ji�~B
d��x���~Cso'����K���
�H$�3faTV6�o��=� B�钶mي+W���W��� Ezz�:H���c ��f������������\�.���ٞ��nf��|\*�T�7K�P��IBJ�]�&��Q�n����T���
��B�mذ ����epkA*7s���#{ ��vA���Z�ih����vIݣum���`]�ײ�}���@�>_p���>\�(�7�$����\80q�@(�v�iάY�i�P�A������<y2V�Y�k�7}�$��u���|r�k����5�_�/_�I>������i�{?�;O�?~�o4h�Ah�����4������~��+�w��]����	�].�Ck}-r2������ � � �%/��n����)�����b}���/�HD�]�ģNgΜ��#G@8���0y"Q��a�e��s��AD����Çav�l�[�9Dg��1e�tܾqwjjA8��{��ҥK(..4"v�iF�����Bd�������R��f�I_H����FG{+�32MU�L5ȏH��Z1Tm���n��� �E^~>�&M�}�\�}zf�]�_�lTm��
�u�"qm7���#K�ב������-��k����r�:Q���������]۽N�%K���Ө��AD<�y�&������|w��3�.(n�!�4E�����O�f���{�m�H�v}M���g��ĵ=q{l�o-���Xǌ�Ǻ�Ǟ��@8�;v�;������ޗ�(�N?�����V)-����]?���G��B��� � � �6Fe����RS�B��[�7�������/�^�$ 2� ����/uz���Il�0�oq�rD��H���Ukp����׃ "�|r�����u`����>C��'�J�aצ�����4c�������#b��1���=E���$��@ߡ?�����&���ڃ��I���.t�����*E�2so���߅�N�����q��m΁����,��ٿpm�8���wm���q���Ţc�ڮ�3J�����9��#�Ӎ	�m���\�M>	'^	Vǣ�m8�
Ffgc��b�ٵ��� ��'l��o���yX�n���	��Y�^]#����,�ڵ=�zE ��k�l��z '�CsS3g��Յw�y���w#N�`L~�`A*�~��D�M?�;����r�6��`����ټ�@AAa%����+!�ۭ�bE��]��=\o^_����fR�\	g1k�1���Â�s�k�N��� "444`��]Xw�z\��	�6�sFb�외z�΁c=��(,,�z_N�So��~
c̱,c�wpWB��9w�Ѕ}�zA��;����m���B�a��~$�o��26��Ȳ�i��{��Y�(���#�ߴ���xKP]C&lק�E��nاt�M�k;/$GB]�E�;`��n̄�\ۃ�����w#C�+�<a�rr�y�&rc!"a��۶nò��1y�ܮ�����z�x�
��|��O�f��鶃׵]��t���f��|rzz}��x�A8����<���|�j'�dt��"bB�4q�<X�;1(�*]��d�\�Y9�n�AAA�d�5�C20W�X5��-���u}���ZbE�8��/Vi6l@o/��İ��1kn1",�7nO
�n�� �xÄ�l0Ͳeː7:�/] Aě9���-t�w�p���x��w�G�G��+LL��Q���3�c��!ۺ��o�+��{^
3�"~����,�Fwk���	"�
A��봗�D1���U��
�$`�C(�-�ĉ8s�琑��}����.�A�@[�݊�vٶ����������Q_m(�/DV)-��k�I^K��(]�ż&�<�|�pm�pi��d���}�i��-�� ��U�}|'� ����㨮����vu%����tc���$-J�vY��|�qm7����<a���&N���!�-X�G�Ƶ�2΀Mm�e�|�_t\*�ei�Q�7-`�}6����~]�"P�:1D�.,��AAA	�0+-�u� u���P�wy�v����B��=`��`\G�o(�?tj�_,Қ���y�f�bQ�R��$� ��G�)Y�[�n�֭[ �H$L�4e�<�v=�<��>2c!�Gjj*�.Z����pl��o~�៵h����iA�?}�>����2w��tHM.7����FeNECG?��@�;�31��.�(�S/H+����a��d	DE[>sM$�fg�`�b�ݩ��o���BP5�/kU����ص]1�D���z�u ]^�ŵ]�7�`�����vC>Swx;\۵<BZ8�vv�,]�gN�DMM� 줲��>؈G{Uwj���T֠SG*s�0+���۵=�ےk{D"z]��������/<����O�Yg���o�駟���������ZV��$�̂mU�J��n^��$.�������_�{꽥� � � "�,ۏ�:]Ǻـݐ}��6��s� r�(��͈W���B��7����s�/,��	E �x2|�0�[����C[[� ��ƍ������PE�]� �x1y�T�,��{w�p��߾};�z�)�	���W)1���C���������ٟ��]���Bۯ��$pw0�n��� �`�5q�1 ֽ="�&Ó,��pTTT`׮] �Cn�hL�2% (7���=��Y'h6�KU<bz(�v�X^�.��È��b��.�ˋ�aP�&l7n�H�D�Ll� �v���ŐU_���4�,Z��{����,:	�p,`�����㏣������
��v+�vc>���\ۍ�����s)��[���[�ApA������;v,V޷� ������GaݺuI+b�4���B� ��o����e��pmg��-l��؀)��p����'� � "��uԡ�dj����B{�Z�ڦB��P3��	
���x�/��������ouq�2D<�;K�������1� �inn��m���C���3�oh AċE%K�{�v2�u6l�O<�����Kop�����Xs,����9��)���K�AM���.����7D| ���)�B_s��P��.sq{�O��nezAх!<��
�ƂT��� ��=.YQ���=2I��k���a�w��b�mF�/QShG�ڮ�7�B�(]�un�>�˫ ����+�ε]_a�����o��������9رu]�A8���wՀ���l457��Z���t� n��]ۣ���A�e�Ć�Y]"��E��ȇ�k�,�C?�S�O����3x�{�3����b�2���*+K�`�b�2L9�sF�?�7��� � � �2-׍֖fddd����/������Z?���e��ϲ��ݫ:��az�,d�$Q	?&M���c�c׎�$�#�1�>Ý�w`՚�(����JD<���Ŕ�p�Jgp��%>|�W�vP�^|�7��ͱB���K��6��̌��Q42Md�H��`ƺZ��rK;�C_\���Aޱ/����H�D�CɅ���]�f�p��OC����tm��D���)��R�9/�W�A����!/X7�S&�WT��KC\�=��uTI1$j��g�1�T0[6m� A��ݟv�܅+W �`,���	n��5sa�>M��]�%"x�h���/76��Q;�'�k��,9�6���g��[@8����˘5kV������1���Bwq�A޽P	��9#���zK� � � �D1?�]u.i�z$�X�@`����~	�dcoE����>�1�8���L/����f��I��?A��`�$|�%˖"k�\�r�.^��7��C&���w�Q�N��ބKb����+ |7�*��B���ںE�}�hH��P��S��xGuo�M�n�� t҇R�tr��t�v��_��i�&ܻw�3`��y狢,�k��z���#����k�V�G�B����J@6nH7��<"���n���W.�W,����%"x�x��E��n؋�OwP��L�2q�S\عc� ��#���x�̙7�5�j�(E�&n'l��(6@��؍��sm�ZD��H��$�v>���R50z����h�K��_�����B�߯�@k}�5L�J�&6�.�ܬj�m���_�wȍ� � � ���(��ܕ�b�3P	��|��8ت��8(Y���<'^��.��ѣ �ü����
��%�����]�]%�Z� �ͩ'1s�L��u��ID�IOOǜ�p��)΀c���a����ǲ|�1���o �X�L�MM�t�r--���[r.��Cw��b�OL]�M7�@�Tq�J�q� =�/��F;��s�=.2�3&F��.�������#qm�jl\%����k�>���ntO룉�c��.�'�{N�bH�;s6���� �H&.]���&ܷn-�S�tm����ѻ�G�w�G&X��W�/ŕ��>�(^��@86 ���1j�(�{����W~�aA*�t�)r�>ՠ,`%k��\n�ٍwR@AAo�MCg{��Tm�K��z p(3�@���=�dxe�o�������IӦ� b�w�_u.�;�ښA$W._���qx`�Z�=x��ND̙6{&�]��֖���۫c������.��vc�V���X6Ɗ��P�����{��8�3��IV� ���pW�"EQe[�eK��ܖ����ǎ��wt�an��|�ϳ����;�s��ZIJ�7p�DQ�DQ�	� �}���UY����D-�
x~VU'��s������y��@?��7��i��B�{�R�>���0�,_2��=� UR��,'��|�g��ӧO�ƍ �Ał
�۴�,��n��$~�r���VXk����v�~��'�>�l��;���?ˈk��,)�t�x�ܶ�?����!�"<��={�֏���A���z��L&X�������N�S=�k�;*{��N֯_����p㫯A�3<<������ T07��L���|����=]�%+�M<��9~L!�B!Yd��Q�N�FX�ܡ�jT�A��/�c	�9��Y��fk��ʺ���o�>��a�s�CM�'$e�exu�wp��qR�G)0>x��a����q��Q�ID_b��m8u�8H~����#jjj����K�M�c��{cY�"w���xl���7��d
��ڊ"�<Ei��TЅA3��I4�A*/��$R[Q(
ͅ��M�pFc����m(.N\��"k�k��Ĺ��w-�v�X�v��=^h�3Z*qI�5{�Ե]��.wmr���<��%΃];v���sx��B)d������g��ס��$�����v[��vؚ�ڇ�4O]�����+6ۮ���'�����?����>~��_'�w*l��OM��:1X_�'��I�w�[&"��ť��9	B!�B��X_fb�I�O�N��.�nu������������e�C�y�l�W�}���Z�-ES�b�I�V�坻pp�LLL�B
���~>p���uܺq�d������Ԅ�O���GL�۳g~��_�+�1��ϸʴdް(�7�\-M"rǰН5�d
��-�/J��l�%�T��|V�T��*�� ��H~d�彳�G����b�Xb0-�v�l��N�X>�퉢�]�����rm�	��2��n����Ů�xa���8~B�B�\`||W._���;046���Iq{�\۝������]۽�0�]۝hiY��/<�s�ς���͛�jS�w�V*b�����qA?%����čA��En�Bcx�%%"�H�k��j�ΒB!�B��֖bL������8�Cw��ļ5Q?�|��4�>���<`��;==�c��@���=��LR]U��݁O�����!��9Cq=k[����?0 B2Ŷ�w����h�'������/�"k䣁Uf�+��*�5�r���4k�9`�����#�ho,�W]S ���<dQ�����9H%��bj�'*���� f7�����[wn���E�u@�v�ص��ێ�%��$��rc��n��m��䳬���bb��w���Z`G�2�ɶ���կ�=Ч`������l�\�ni�k�Ҡ"r��,����D�
�vg��o���/c��Ey�����
'�L��M��C�����P9�!t�D�U��=:�$�����PB!�B�m�c+N�I�}�T�C�1���s)vY�I�:�X��m�l^�����q����`պ5�^TB2E]m�oڂ��|J�!d� r��~�-��?��^Fo?��HfXTW��m��{�6�z���K�={/��6�2���Xz�=(�1���.���ҕ���X���5S��$�P��gT�i��BII�+q�=@��`�A*�c�ʌI�nՃS�n���>��#��`��%hji������ۨ����w�M�vc�A\ۍMA\�ѹ���y<�c��y��%�w��5����Zk��D��a�vC/���w���O?���!d."�e���?�'o���؅|tl̼�ˊk��|�\�>w]���e޵=���=�������k����O@�s��A��?��.]��σP�߯�QC`'�>�L����>:2������$!�B!$�hZ�]Rw8,w�l��_Ja��r>�J0H]�m�1E�yBII	6<��d���&<Ӿ�����2��5q}{�W��W����B2������}LOѭ:ػw�.p7���XF�0�1�S�n7��qsw��c�Ǟ�Z� �9(p�3�o)�4���P�z}ø��h�G��2��L���ѣ�{�.H~�L��-����P�����̵=)7�#ub�	�-�s׮�qzRk��K�f����vS�n�gݵ=/�2  ��IDAT---��gw`Wh ����������?}[�L���H���_Uۏ��>L�%l7��&=�so�u����h��M/�et?���a�LLL�U��[��PA�<]�
��]wX�d����*M��v�2����XW=�/��B!�B2��R������B�']�J�$�5������=_h�/y�l��?x� ǎ��mڀ�
�	Z���m�n�E!sq�s��a�������o��q'I����}-��vD=���׍����=ch��'tw���9El����A��[��=���)(p�3�!�H\�|�}�f?H�ωA�C{�\�{;gg���VbQm��$=�v�Kz�]�e��x�Tl�oʞk�T(���P��rѺ}q���-vm�|q�Z�⎝طg/���A!�q?��{�����? RY�!�(���^��Y�g��=��h�c�/-+�k?�>>z���������~�;�	
*5��Tc�*j�ud0���_���%nw82�Vڈp�i!�B!�d�5U���H�^}�1�f3ƒ���r��	B���y@?��/~�ᇘ���]�@Yy�lh!�`Ų�h]�G!��u�=͡����zN��}�~��ٰenݸ�ɉ	���={�����=����D�n�c�'��$b�'�����X��uS���!(p�#*J�0�߅�H�+a�-lפ_*���U�@�C��08eE8��<yD=�ܸuK�U�_���m{�)nw�G]�n �k�mC q��Mqx]۝��Ko����Ч��n;�D�s�\���w���p��45c�Gs�2��>}�!^}�UT-����`V\�eq�˹��&��]۝�عk�9���~��'N��W^)�A�p���V�_��A�V��g�'�˖tNH����{�B!��QF��+�%� �C�Y�f�%��r�����wOI��g��S���A��lIN�'$U�`I}#�suB�<���I�|~�~_x���%��X�q=�]�D=��~��ߢ�8.	Η�_:�M�3\�/��0��rs���M�D߼t�7ւZ��@�{���с��gwxT�]��.)��v�`$�UKi&��P�� �>��LMq��|`պ5���,��I��-�"l���K���\ۓU�Ɋk�Dt�ˢk�=�������nۃ-N���sm7��[7nƉ�G���B��>|���z\�><�ؚ�k���eB"V�HGܮֵ=��`=�>�܋$��o����
���"�ֲB�
��Ml��<��]�O6����-�XE��Gk��M7!�B!$c�o,���0���m�mgc����4��rq�b�s��B[���}<x>Qς�J=wHH��_��zp��iB�|���s�ȽdU	����k7��ͯ�����Z��oGG����#c,�5��Yc�'�k�m����K���C���1V&��=�h*�H�ؖ,���v�s�ҥ��b�l�w�C���a�����G��G����v��z(�vȄ�]�!�D2O\�M�e�RѺE��Ի���q9\��KK�u��۳'�u�B�"�[o���bhH��WSq��h�8?q{�D�����`�v���׵m�v=tO��@�"��ݻ�+Vx�� T�A6s�f~�����1X����1�	u{=!�B!$S�/���ӈ�D�$ͽ�vc,-i��7��O��웙�.w?�I�s���#L~Q��_�6nۢ�߄�C���(ӊ���#cB�5B���Xݶ7o�!�E���߲	��^ Qχ~���1���c� @9!l׵��9Ck���_�\7�;} ��<�4�/1���5He=�]�T.�T�]9�dKt��:��C8�vQ���%l**�ύ�&���E�����um�}�o�og���]�>�vm���\��m�曻�ř��D�L,���q�2�vY�]����f����`����d�^LOsV!��]���[XPQ��1�L�L���q����44���{���gB�t���G�"�����?�D-b��}����ì��E��=�~Խ]��`sd�LO%rO�1`e]3n�p50B!�BHf(��������B#?(q�2Ɗ�t��š=S.�n�3g@�#V|^��������*���s�A!�x�v����Q|{�6�-�֭�7׿����Z�;�G�����3f.�N��F�c,�O6����&�֮������D�[6�k�"����=O��R��i���H�4�#��Y\,N�A�t$U&q!��l�<8e��O?�C ��6mt���X��r������>����ԉ=L,�Y�vY=��>�"Ϋ��W��h"NK�h���g~��6{��G��%��-).Ƌ�=�=}���@!�ξ����O��/ޣ��zY:��a��abú��#nόk{��l��{�fGp�q�&,^҂G;A�"���o�F����B����hbl�N���ܯ�l,3�pc�<#�n��q��B!��6+�1<4�����vc��e�9��W��&��`���՞�e{�졁N��y�V����Xֲ͵8}�!���9}/��&�&q��2�}��-�q��4�Z&&&t�;�7,dw�p�����x-�/Ku�!W��EKU:g@҃�<aI�F�	���%x��̹�)�U�]�.�n�C�_Ygg'�?���½��L����yn-2��<�mv#^�(� �(ϴk�m��`�q�qm��M���.�w�m�pmכ)qm\e��8��ك��"�b�ھ{?ޣ߸Bq#���}���w03����������26[�����;c�9�7�������Z<x�;��޽� �f�s���;:����67-�CR�n�2���u{-!�B!$]��Mc�ے7tN��zXr����9�@&l��������K+�}��' ꩭ����A�lYҼ+Z����	Bqs��i|��W099�GO���кz%����@�"&���w�����|vgϥ1���]�W�����a��#�� t��	�y@$�����r��E����C��.�Q܁���/*�r�̰o�>:=��%�X�a}�\�MSp�!��#^����G%���}Kc��v��ZM��]�ĵ]K~�
r�ڞ�b��]�vK�%�6Y}��Y� n*^��8��5	!�x#�����?�+���X��q���.ͥk��~YdỶ;i�ݷ	� ��X�J܃�矻B�:mw��*xRe̍�)2�=��RՀ�A��B!�Bңd�ӎɵ�>�<�|�g���*�M���0�r�'N�����AԳq�2[�zy+���!��q����꫘��BwO7	��;lxf3�� Q�͛7q��y<���y)JOEƌ����c��E�r��Wfh�`�/րj����=�����8��+�K��]���\�Y%.��@�I\��R����s�0��6l@Y½=�E؞�v�����#�����k�`]�k�{��$�qn��S�!�k{B�8�t]�ݓ����]/���C!�������������������Wn/�����\���2lW|z��0��vmڀl	����o�����<x��O���ڸ�x!�+������ʍ��/�����F�1B!�B�cqUC��(++��z���'��V}����̱�h�G�y�l��d��� �YTW��eKA�l�]��׮�Ⴧ@!$5G���?�.|~=�� $,��Z��g�cr|D-�?#�A���X�|�o_ؑ+4��F�:���e�gC���ۍE��762{(p�V.���x$� U½]���s`���w��"��M�th�C�_�x7n� QKqqܽ��"nw���\�m�rm���]��h��k����|a�S��vmw�W=�x�-��v�:a{�˙^3���o��-��k��j�x�{��8q���!��azz�������:�cj:�<�k�v��P���ꚳ����� �{��^__���u���������^��
�vc��RirQ�ǀU$��Ë���P�/ !�B!�̖����POQ����?��#j�ի�} �����3�Y�~��B�%Z���ѣGAԳi���쨩���m;���} �q?t���x�7�q�,��B�a��v�"�Z����ӟP]w�1�\�n��W�,y���q٪k[k8z$(p��F{��x������q~�|E�H|�-���6k.	a�9�%�,ȝ�*�PAii���%%%���&<�wI��TP�%u�6�
m)�c�����zLQ�Ġ=4N�xow/����T���񑆛��+~@�O���_&�����>�"�(��2��m������K��S���e�[��������./���q��m�`rrR��/�ѿ���e����X�;��ק�~�Ǯ�~q���K�7G*�]|߆��155�����!���a�O��B��v�j����]>p!o�$���gltT?��]O=#�n��0����8~��_d�}�W%��ݻ8qԲ�n�z�4��`4�����A��2�os�!p7�WQz���0�֍�.�X��VC�OQV܊��|�!�B!s��� FB���XEvc,�������6�!��Bth��Ǿ}�011��o�1�'��U}N����n�8�d�W�T���ÃCY�{|l%#��Ψ�ǋ�Q6�Ϸ��9>1>���,�����,�_�۟=��;>�hEh���:�s���+\[e�����8�t��'ר<�D�Je��n��R5���;/�=U���;���^x�E\������W�[#�.^o�@��|]C��[��F���!�Vy-מC�����y./�ȶ1�������n��}�g���9A]��"B'�&>W��]1-UE�/3½�>;$�R��A*����pHN}�g?R�C�D���\���1!��'U������t�/>�m;w���~��n�� ���t��(�m�W����_c��u�*�@MZ��vm7�o|�%�n\����-ǝ2�2Q �޻u���(���tm��/�V���K���M�b����X���[�n���*�!�ljjRR�ݻw�b�
�B��U}�B�.�����J�Wy������;�⚯��.+?~�e˖)������G����w���\\��:�=t�}��@�ziڮ�w��t>|�M[6��cϳum+�����r=7��ux7˄����}''���؇��Q��{��T ���O��;w_}�����X���:g��`���1h�����ݱܠ�������~�f�!�B!��)/������D��J�;��~�v��A�-V�<��5,�6a��KA�!pW��?@+�Z1����q��+�
���*���~����ֱ�s�}�j:p333�qB�j<Oh�k�
��]|�)���B�y'�s*E�Fݪ�*?{q�&p� [�y��E����l�T8�j41�B����c��PW]c}rB�
T��}4�w�0�w�|sg����ጱ�&��D�F�:����?6Ѕ�e���etޣ��4��ڄ�2��e
">_������.���> �@�ҽ�(4�z�xq1W��KL�nܠ��uٵD`����v�J�����qM��܆���&M+5Z���g)lO��%���q21z��v�g� q��l��D;����L^p��W���T:dB�\B��p(vo$Dڏ��$��A�".Ll�B��;̽�l�~�*D�A�J]^o��y�N�m;��'�Q��^|��'��]�-�P�^fPF7���=a�pn7��81H��,��6n!�B!���ٖ�D��Y��4�r&�5ۄ��#E��#Ih��kN�B.�/���+W|����XS�˪@���Ps�8�d�/����M�^���4��`�"�!:k\ܬ�n���Z��?�.Χ7^����h}}����ʌ��6A����FI�Kձ�C�.��T��؅�Y�Ω����1��ÙB�g/�7�~q�*H��{{z�׿�5>=zh֓��d��%���������v���U�����\��.�+�㩼�����re�[9u����[�Z�������{c�İ�ޚZ�)�1i���=���cc��\�K�j&���qU�A�El�o���e��Vw���$�A���`�Buf���O?Q�����L<&s�tm��{	���b��y�<�k{ a��<}�voa�۝��{q�g�f�u�y�����I�v���764�~�4|~�*!�d�����K���ft��J"��{��ҵ�u�y� ���f��v[Que��˗�@cS��<Q�޽{�����U
�]!l��:��Ӊ�շN
݋��UIa��/?=$V�R�&�B!�6K�F0	�7�c��v3�n��Y��*v�2�rR(����b��\�ۉ��۶���|�;����S2!����s���/����N�����+׮��s@�!�5B�w�w�m��?̶1���՟5ӈ���]��(k���%���
�RQR���2�^��R7� �u�t���]�m_z��P봐�%;;;q��Y��n_���2Gi�\�=��β<um��~Y=q��+.*�ˑk����5�,��;
��.X�`!�5/֗�"��y���+�TWc���l	�d86#����9֜��=�^p�#�(�|�U�����@�����>}/��r^*eӍ������4.�w�va0����`]C1�~:B!�B	��E19�n�g�t�sf5�r����Y�B7�J/�e��hD-�eu��e $/>�<���s��N!�������?�g/Q�L��x�,��+��cϞ=����\A#�g�����c,��"3��9C��>&��@f�
��R��Xf0���I.��� �]�F�p��}�߿SS�D��½�JP��x,���p��ZC&\��(�ڎD�!������k���\��C7����f�����,�i��̵]<+-)��͛���BH�8w�ެ�ח���J�޵ݽ�t�Ac�µ=��ƥ�y�3ؿ���2��
�]9t�.p�m�ww�ٴѹI܃�rN�^9ͳ�.l}��M�� �B!����o(���(�+*��&��Z;S^	��&w?��\�%?~O��3���MAH6�mG��.}uRB!����{���ĺ�k���o@HD?E��.�9���y�]�vt>0��X����ٵ�=�%:ࡁA�.jƝ�i��Pஐť�-�va0g�_"����V�T�`mV��6>� ׁtVM��UX�pa╗k{\�l=Où���]�����;��C�ni�G=2���k�����<]��u��k�f��n-a�Kvn{��������c�����&'019�,O[��]�%�ȵk{Z��4�P�Ov����@�q��A��?�3����ׅ�0�x� �n��rR%WK�V���K�M�I5 �B!�������d����qc9�8V����X��Su�
E�tG�	��Y**`Y�
�K�cay�]�
B!����_⹝;�t�<x�	E$+׬��Ϯ�y�D�F�s��]�m^c!�9��h���֒���+?���ƺ(��nVP������S��s��t`p|Y���2w�A*#�Z���f���_�ڵk jY�q���ߵ]s��;���;c��칶�c5�vm���]�ʹk{"�ϵ�-�w���m~�s8r�0&&&@!$����{�����/���}rQ�"�,��{�!㱅��&v�Ǻ}��� Fu�����!�u�ʫA��1x\/��E��;����Ace����@!�B	F�D��\�<��˾J���;�I~Y�P0�L��e�/}��Q��vq���:�-]�cG��%��\p��9����12:��~*5IjDf��u�v�
�:��?��?���B=o����X��Bg�ڜL���=$��3�Z���wEll,��ؘ{�A�A����t���ͅ�21s����Q�4^RхA-KW,â�Z_�v�.�*���)�����-�gߵ�v<2��,=��(2��E��f��C�[\�5��C���m�l۴ϝ��� !����i|��x���
�:H"�k{�D��(�WZV�_~I�5�����{�x�B��ۼ���s#R��܍�4�
j^KFl�֋��	8t�B!������zQ^^.u}�2�*J���X���·�ub�Y>1Z��A�xя"w��Ҳ2��YB�P�^�|f>��	!�䎃���;�ctl��bM�Z|}�:&id����nttt��^��|`&���]��c�&���]���7������nT�Uax�ZհPஈ��S����`r ��E�����Rŷy�[�(g������C�@�Ҿy�[ܞ����8��947]�e_o�{S��[l��"H��u�A��pme�˗���C<~��Br���0؏��*:�'JC܋e���c��X��gBp,������8~��r��1������N]��
�ۼ�L��Í�ZH䞘\��
����U�@!�B!����o�_5ʚ\�c��� �v/�, ��ݗ|�E��Fc,��Y��Ŕ/�Ԉ��+/}��}��-!��q�=��~|���c�ჼ�����b������uu9rD�!�=��X�P�1��c���c꠫?M�d�����;�Q:9`.3t��s����U��KǺ%N!@�&�ҥK�w��:����d/̩k�=6�k�D�n��<��қE�b��2�hx��)��k��m�]�5��XX^�Kg΃B�:?z������U�����ڞ��wx�y���4ڔ�Xk[+T`���q�����t��������2��׍!�|���KZ����*�{��c��m)�9�O!�BIA-�0�BT0c�p�v�>�$���ܝ*�e����ٳ �����ׁ� q�w���@�BT011��'O���_��3 $k7�Ǎ/����4�>��XUUU���v~/�>f�=q�縴�2�;�*r7&�['�k�O��џ��R����a�'���RC}=�%�	�\�ܽt��=.{����P�'���h��`�̳a�f�E�\��%9��v[,��z�f���p�>$��QH�y�㊛�k����0>W��Ƀ���������lZ��!�����+XҲ�e�7����ӵ]��`��ڕ���v���';033�C�n��B�t�e�T5��A]�+�I=�*mcc�X���.&[	!�B!�Db}�сni<�1��oc�1�2����Jn�/~������Q�ʵkPV�U�Hj6�߀�7�E?!��C� ���lX��o|B�(�����m���M5����y����yot�~�Q�>4��Ț�-[�����[����Oc�/	�
x�9���vG|��3@2�̠U��{?���L������-˗�_�Ե�^&��pmw��5i��k��===�v-�k�~8~���2�k���W��$â�k���۞�����!������/~�K<z����场��>�>s-"�G�}�X���E���a�F\��9�.^��G�����3�0���m��'OZ:��Wߺȱܠu����{����)\�!�B!�x����c(/����c���T^��u�w�0W��lݝc,���� 456�<R��oRG!���7����P_���� ďu�S��?:v�.p���*l�s�3��˱��]���l%hy�ݥ�D02<���b��1V(pW@K�(Ɔ�]\IrKR}��:g��禘� �l�O�>��<*++A�P�ؠ�ӆ��tޔU���k��c�ص]���U�+.�k��=�gQ��|����[����ܵ��n�v�ٖq������BH� ��}�!���?��G�΍.iN]���fKD8��]ۃ��˻)pW�p�?p� ~����B�}Iz�A*�>���]��`W�����ޫ@!�B!^�����D�՟c�e&��}'�ܡC�n�c!۹���=��ܿ�.]�{�B�j���j!�C|G�m،O�}B!�C�ɓx�7q��1LpE�C��4/i�㇝ j����n444����dB�1b��4�C����G��n]�9�)�E��������N/H(pW�h_ a������J��
�}���/���l
��l$��Hq����>�ʵ��!���v���õ]"D����\̵ۡ��䱻]���/�P� >|B!����0:N���v��ӄ5q���{�ҵ=xl����+�t�2<�wDN��_�>�x۽���`��Z��>w_[�ܠ�@�1X5�׃���Nz�xA!�B���M`&�Z?c,�jSAͱle-�3r�~�����W��]�� �q�z���qh?Wi'��|C�O>x�|�U|z��c��v
�bc�򗿜�X�9VPc,_m�Ĩ:̣ñ�+@�C�{�i��`hp@_fй�� ����b�nq��!vW׌���Ln��3�P�� �ѣGAԱz�Z]���Kݿ��黶;��Brdյ������kΥU4���ˆk�����ϊ��c.�DS]=��B!��ݻw��e1�����u\ܞ�k��a>���Up,6�}�5���/��������>�<��e�<c�I��N����^6� �נU�������>���B!�⦢�C��()-�:�K��i�e:��_��+Ih��v^�sn04�Rˢ�Z,��$�w�¹�g111B!����8._���}g/�!^�,[��j��������=����O���g���K��}w��l��OQ\�SL����1v�ȗ�%œ_���{�A+.�v� U|[�6�%g��g���ӧ ���>~�?ϕk{�ܚ:6���{���µ]3�����0˲��.��uo�������A!$�9{�,����(-)��d<���{�{�l���!n/t��0�Yrmw�nܼ�,܃��!��3==�O�����uW�M�u !��l�)t*n7K��j-!�B!�8��T��B8�iǸ�+<sp�jݥZnЯ�Ν;�v��:�lh!~�]�O=Aww7!��/O?Fcc#V�\���n�/V�_�Kg8B�ΝÓ'O��ܬ�V�Ξ�Xn�e_1ͽ�Zʼ�E�.&lnj*ƕGS ���=�,҆0������E�*�[\7� �񭵖ƙ���P�:::B�d�e�+P]S��s��.���n��=���"K���z��K��N�x@�v�_nѺ,\ۍ?a]�m���69�q�3�pp�~]�E!�0������/~�{��k�G�<.����\���⋋#x��p`ߧ j8q�.p7(�z����������?@�\%���d�z�1�k@=!�B!�ɒ��ޑ 9C�r��֜��,K�3�kn0SBw�^(V&j(+/����.�QW[��E��8q�B�k��W_{O�{�?�Bd��^�k��bb|$�LNN���w�y�`��Y1�
l�%�oK܃�#����)\	
�9DӢ��1O� K&� EfR=���R��z�,No�ʏ|qf0��:�nhϝk�ԉ�ܷT��ڵc�Q��Fyn\۽�SV����ڪص�_ ,_��n���� !�"	x��|��W���q�<}��0�9�ӵ]���۟{Gb�X�ϟǣG�����3W��M��3He�c;����=���@��&<�$NB!�B���w"�#ghwp���}����G��DC����|�;�����k�~4!2�ul׶طg/!�G��o��}GҀ�H��m�*|}�:�N�<�܃�_B�pu���ːǵ��7���&�Nw��jAVf+��j@�A�{io(���8��+R8�[Ov#����z�⽐j��B��2��T�/^�ÇA�P]S���by���ڦ	�ø���oE����rm�8�;�i���k�Ȳ?� =�����)��ĕ���aQ-��2D�R��e�:�?@u}��z>���E��*���=h\��JlںW.\�=bb�Hڿ��#T�Lݚ~�'�t�}�[�0�,+�M<O��`�R���A��!B!�BH�����QVVp�gs�&]�ٹU�U��]�]1�|������K�P�8wW�[B���/���GBH�133�S';����p��9"c��u��ŗ��W��ӧ��ۋ��:�u&rx*�~8M��ew���}hw?�����j�&YC���.[��q��A��=�����Lw$� ��%.�R�V��ևI��T93ttt��Q!k6��N�"�B\@�n�C���":w�:�k��#9$qR�vg=鸶'�е��[k+��eµ�-�w�E۷o�BB)p�����ܣC�;�vyd���g�����+6���θ�v��]!'N���A(�A+w�#����C���=�du�r����X�e �B!��-���I_Мab��)Μ|kN�5^��P���C;s!7�W��cǸҜB��.GyE9����]��100 B!�G__�c��K����� �ɂ�J,^�D7P#�gllL7���O~�W9����]F���Ksk�s�&X����tpO�7L����M��7	�
�sH�t?F-.n���.^KZ$���vr��`&�4^<?z�(����u�J���� �+�vHE���.�;�|��]o�!��ˤk�S�n��̵]r�b���M��q��ELN�B
���AUe��$Ǯ�i�3�ڞ��|D��k�]۝��[W���	]����3g�d܍�U�V2'���@U��O�.{]�����{����c�Z��B!�B�QW<���9CS�n:�Y'�5��rp�c��O!�S!&�u�n�{;�SQ^��e+ph�B)\�~v?|��<~������C��	�{
��ܖ�1�s�碤s�!rO��S�bELc얲QP�~J9����Eq�8��e�*Ѐ����r&�-��Q9`�ξ�^��;w�u�*��%�
�k{n���횵6��Y��[ږ����k;q�����`z|
���!���gddCCCh���Ӟ����rmϥ�<h�k�W쮗^�G��H��'����?�K�z&�vbݬE����N���{����B�>:�����; !�B!$���S߾�s2m2i�tp/
էI�$��jnЯ����ϟQCuM5��@��ﾰ�!������#X�d)�!�+�bxp$�����WUU��=�7�}e���p�����eyC�?o����� �
�s�Ʀb̌Π��18�y/Q`�������Dŷks>,3��}	��c$s�.6ѵq����:��}HE��x���6y��]���tc���5�µ�8f� �&n�����n;N�k�f��~F��C\�6�]��� �B�O�>���8JKKuA�A�\ۥ��tmV��}�XU��N�l݂O�����8H��UB��d�Z��`5��TԼ���`��U���A��bU������B!�B�ʺb������ܞ�Ni���ܽ]�:��E�2
-7���۸�-��ׁ[6l��W>���B�����ʲ�_�.���+�d��5�z�2H��uBO��of5痩��i��m�wHc,i[��Z����� W5���4�?����1=.wr�<�mU^.>�p�X���� ���u��15,��E}�1��*�������d��0��y��n��S��)"O�3+�vs_.Q|"*�<.�k;$e���'j����[���|B!s�O?����]��|�s����У�tE����#nψk{��\��[��l}vΝ>�{:::R�1�Q(�V�y�T�8�/7C��+s����]]U��Jm$��2B!�B�� [�#7��7�2�$a�mX�D���`.���E���������@��ښE�,-��@!d���ߏ��ZTWUc`p �Xi[��.�����#�����I�c��.��Ԙ�m�7�c�9B��7�)�9�=���AR@�{����d��r�0��b|1S�.h	;+se����۷q��5�oڐxfum���S0���2d�v�ݽO?�[���C��9��"xM�ڮ7��ڞ����d��ɏ�T�k�H�qI��n�}<,�k���˖,��{���!������4<����u=ql.X.�ϥ�����
�}�
�1::�S�N�?�AN��a�3Y���A��uҨ�=���D/q�&���ղ�B!�R��`4	�3�����Ͻ�.2dY��PyC��3���g�p\B+V�����Xמ�?�}{��B����x�7���A �ki�rܻu$��`�҂XYLP8+8�ۗ��6�[֟���l��L�|]�#ԗ�������-���}�̅A���pg�8ù��E�:�/���{|���=I��r�d�pa��J�J���-����]��h�9�'��b�]����Ԯ��mq]ۭm���g��n���n������ڞ���w�]�%m/))AK}#��� !��e�<y���Ge���$J�����YsmO������_�k�3nqK�._��������w'��
ZO<D3�UK�X�p���)n���	�Ep���B!�2ߙ�N���c9Bc�碐��3yo4w�$�s�~�¥p$9VErͪuk@����z	�;N1�O!s��}���z�9��x�XY�n-��E�p���91�R�t*c,3.x?;��u�߃���1��E�?����%��Fyy�t�JvBk���e������_ZǈT|����R̞�z�ЅA+V�BIi	��v���H{��C&X���!n��_�OO�6�B�`��k9pm7��rm7���gp��AB���8~����1<2,�N���vmO'��];)pW�����/��/(.���@Sf���[���T�����ܽ�����X@$A�"��@!�B�ǈ��b�p��3�c%�&�W{v��*�xy�6Zn�/� j�k�Ǣ:
8��%--���Eoo/!��]����r|M�x��467�zQ��Ar��3wٶ�d���򑜈�9�~�S7<<8�������Z=�h�D��7k�"dO&ӋBX���`b��O�X�����9��S��u�������ȵ�C�̵]V��8�vmw��)���,�����cȺk�}kC]�߹��B���ߎÇ�ŗw�Q�cK�4�c�H�wV���;VO����k���6���155�[?~��W�b۶m3�4�}şG��W��#��WK�#nQ��2������.!�B!d��^��:D�~Y�m�e`�Zͳd9�B��m����܉�֬!Vĵh��t�>B��\8?|�M|z�W� 6ZW��Ջ�Arϱc��?�)�G��z&����XN�v-�O��׋\ۼ������K������!�XE��*���<�U����Uk�)��~�j6��:u
��� �G̮Nq,bl�k���{yP�v#6��=jJ���ܸ��"x�{=�eڵ�������5mi�btp�B��=�`� ������y���.���-��xY�oYy6=�W.^�-��ELwٶ�hJ���V6P%��8��_7��[��2p5=,�Ț@!�B�����c���_��fX����/J�nM
��;9�V����v��e}������� �ʋ�=���N�B��@w�>s;�ن�W�"&��W����03C�o��}�6nܸ�u��e,��9�P�X��C����Z��L�n�6�	]k�7�gM�bt���}A>c#!b��C�-�cWI�u�j6��g��am{{�Ea�ʵ=�I���x�>�wm��%q�rm��އ�]���{���z�ҥ8�!d^r��A������%_E��(�^���;��m�N��"�[������|h�|=�{_�r����T�"��D���[c�V#��h���sp�B!�����H�+��3�:¹����=˰�]I�Թ�B��m;�<�X�b9JJ��1������8���@!d���ݍ�PS]���~"(�(G�t� �[D��̙3��]�mn�M�Mf����n�O�7L�����T����qq���,����(/��]n��k.3h[rPsX��pc�q��Q=���z�2�B�.�Be{n�6¥@<T՟�c�[Uu�>yj�O222���N��s�%n�z�L�n)��NNOIE�1��6!�k/��^624��;��l�v�L.��3<8��%mu�[�ڃ~L��va�B<�|�z������1���(�[8��ttT�(����$*�]\o�o�����cW]�������������=�8�T�?�֊��|�޾����m�J�x�9M��� z�{PV�>'��<�]$cn}�m����*�^������r��鍝�S!������p�z�.*���~/��%��c]KK��{�a�)�z\�[�U����U������c����� �B!��C�F�~�5o�y�ܭ��d�<�Ù3ķ��W��T��
��h[��XY������B�#';�Ə���C�A�AۚU�+B�����-��?�k�2�rN47��~�`K����C�}XTр�QcyA�{�YU3�'bqy3OV�lk�������ݍ�ĺ�d�X�m�}�?~��K��U���'�u7-nƂ��1V\�]\��{;��Qص]v������������!�����.DF���f=�����r�����>���Y%�~� Y��&����U�m_���_�^����*e�Kq�UU���MNN*=���Re"o�B[Q�8n����[u��^���.�s��{�$���_v�b���M1�N��.¸�K�SS�(-+Eł
�}z�7���Op켏{y�wVK�k����Ů���y�]f�����$�������o��u�x�<2��eg�t�DY�DYGG~�����@S��1�J�C��#����S������'�p!�B!����B��_�sr��d;ۜ��o���(�ܠ_�Çq��]=O!C����VF��&�g�Y]�dp��&�|���U6�2<8������q������7��=59��ё�c,�u/nlҍ:��ef���~ܾ}[I��H�����J�Wy���D��7*�]\g��OLL(�0v�u�2dS�ً���
�*��w�?�_����x�+ku�����]���*��W�;/Py�1:<���^�����5���Q&Ӯ_�cT!�s��W��������?׍�jk�N�\\�����ͱfk�e����iIM�|���=���Р��=�Q�2U��8��35\�Q�e�
ݓX��HY�K!X	N�>��$za�D�@t�Ŀ����V6�^վN��01��ş�']��]�8��K�l]��5�ㄫ��F�Q6��Bq��\��.u9�J��g]�aQ]]��Q�8��sm7%�	�{R]g6�ɣN��׹c�a�}[�dmw���m�ܾ׮|��VVV*�����j%u��1h��~q#�5h�����c����PU��cW]��]�`���W��c����^U�b�l�ʖ����q?��_�����2�ۼ�"tKaoy�~�ײdI8��4���?�޼��-�������o��������Bs�~/�!l7b��\͋'�<�m�v��"Μ<�tQyo��{��.�� �N�a�)��r��������;���N�n�JtT,�� B!�B��CLx�&��	r�6I�<p�0Er0��-^�"�s�~�'N��E�^�qLU�3Ch�Jt��c߸u����ݛ��b�J��񃇨ZT��Ʊ��L�����z���x�Ҝ�+ηm�7�??�D[[T!Ė��y;qݭ��QR��cW]��'O����_�@屋q⮮.,�<x� �/VfΤ���B/��ب��|�ο��k8s�FFG�Rw_w�~��'������z���z�0�=��_��ŗi��{{чƧ�{���>q_"V���<�r�nc���n6�X���9C����yC���e"��"�
ܳ��`�Խ�s	s�����BPQ�\�:u*}�	���^��:�I����wmפ��Q�X-h=n7v��^����z��}?�D�.�vg�E�u�%�bN���N��\��|_ض/�\���	��L!��$��_ÊUm��띕�<e��� 6��ݷ� qY�ͦ`=�8y�<VL�\�f5n}���b�"&��H��B�8Д�z�ĸT4�@���Ⱦܠ��]��><4��M��O�B!�BH�����܋�},Μ����;,�ܠ_��s�@� �	1���.�t?!��Ǐ�{���Ǐ�A��U����>��/	��l[>�g�����:������qq���JͰ$⢉�Xj&��g�5�%������C�e}q�J����Q=���z������ ��u�J��m
��o�3x����2C�n)����p��sm�Ǝ�8M��!Z���[��ʵ�^��,�|n�}�ڮ�o�����Ï@!��%�֮[��/D�vqgnE�qmOI�]�5!M�z�XQT�n�{f�3�+@�4q��E���y*F�]=n��M�9K��ܓ+���|���o(�ɻ�B!�2��[P����x�P�<s�.c��
R�՞���,S����2E�� �o1ћ���&,T��,�/6�[�_~�\q�B��F�,p��-�[�_�n���u����-�=Zqq\N��9�L�!�R3����shC�+?'�;����Pʋal
D�Ydբ�I�/wl�T9��!�L>�vb�#�g2�Μ9Î�"V�l�!w��hy�LH���n��B��[�?�]�݂}{���n�h]�ׯ}��
w!��9�?~�֛���P��v��s��&�����u���˒��=���K�.�wٶB���4�%�V�GX���:�K�� !�B!�����nmZ�|��_�|�9C��$�z���_.�Ο?�����C�vbPZR���&��!��o��?xㇸy��DDg��6
���ݭ�mݺu����+���Y�cYs������ ���b\��]�Y��dc�6o����J]�Iz�,��P��\��{�CCS��8���^�v[��k����r���K�s��no�۵�k�(?�Mu�p�!�'������Eii)�'��Y�g޵=�"�|um��՝��7��W�����J�/)t��x,�U��y��k�s��r�ց*�C��Pl�t�#�B!d>�T>��ሴ� �����v+�����&��B��m�3i�E�!��+���K;w�tG!�'�;N��gw���� dy[+�^��{�1����]��Ps�nc������Jهv��f{��;��2�H�KL��
ܳH�Đԩ�ӅAs;1���\N��`���2`%ܢϞ�M�
Z׬��k�'S�n-s�г���ƻ��̵]Ҿl����ݽ��q��ז��8s�!�/�>�����yx߾a.��k�<�����^�鸶;c7?��
N]]]hjj�_���l��S�b�A�q�=&0<Ћ������B!�B�ҩAL}�ܡf�1�ΤyC,g�О�O�;�d�/��iC�	�$s,^��ee dQMF���!�)�+������@�9��T,�@��f<�|�[.\�������b3Ghbl2Ӆ�P9C�������E��h��r7�g���';��봗z�/�fhXN����^N�r��5W�u?�Ն�������=m�e}\�!�K�M.q:��\�]ù.x.\ۭ�5�E��fM�%������j���q���ѩi��p� B!ވe��q-��Ȉ�y:�����gA�J��`�����d՚�(+/����џd���)�;w?�я�&e��!yg%���x�V`���pf���������r��B!���9��@_�?q���cY��󆎜a�r#�|���c����|�� �g��V"xa�N|�w!�/Nu�����*�8B��;�G�ń���j����zߵ��1V���]9D��}r�7Vy�
ܳD{c	�#Q�I�� y��~�ۉ��%;�ˀ�ŋ�L��բfѢ�+�v] n/�J��p�>$�A]ۍz\��ʵ=�xoB nۋ-�.lw��;�O��R��������8�̆Mؿ�B!��t���Ż��pm+8�� q!bϵ}��vQOqq16lބ��/��+W��w'�ࠐo���l�xͶ
��@Ź��ʚ(nt�B!�2XU_���)����'����2ł{2��4P�s������½]L�&����K�-!+W����o�U�	!�/�1�4/_����t���m.�9���366��.�����Dp�6hW:���������`[���߱�Q�TE�98b��,��2v��Ig\H�\�8������Iy��|��ԀեK�@rOۚU0��LK�ε]*��	̽�c�,=�v�@�g��]e鸶Ǐ=*�<0���)i����zt>x���	B!A8u�$v<���v%����е]�����U���k�m~f�
8u�m@'_2�c��r���@�UE.w���dc��b5��B!�2�YU5�����_�����p�~���}$���!���l�|�2H�Y�b"Ŕ"�w�5fM�*����X�BR�����7ߠ���%/]���x.��w'����˷����2ǒ<���]���kk4t�8`�2KTFG0*I`���w�v��yXќ�����$se�J�jϝ;�{ZW�
��.uI7�,����0^'y�%�V���no��Y(��d�A�C /ڑ�v�h�C ��>��F�ڕ+����B	�Ç�\��$�'����H΄�<G��h����cκ���,VVϊ�V,�����0H�x��n޼��k�zƨv`�4�];�۵�����AE��1�zE=!�B!s���8�Nm��;��^1*�Ê�@+{yðd;?)��={$�,ok!�m}�/�ЂBHp�^��-6���/@�7�W�R� g���A�[��⢽�%Ϋ��1	]�
[S,�(��2a&[b��,19�﹤�|v��������(��.^drPʏlX	��������܄+%�s�v�gܵ]&��/��������m��ݝm7۰�u%>�u6ru!�2w8|�~�֛���1HA�v���ѵ�3>����Ѧg6�ܩ3 �C�{\�pk֬	5��O��t��V9�����f�8��P]ր�q�?B!�2��w%�}��\��R��&��K��-&t߿OQL�)+/CSK3������e���!��G�aӖ�().�����e��e�����$H��ꫯ��ى%K�x�D$G��Ѩ��;�<ٯw�}L�l������P��j;�g���FGFP^^�q!�;Nr���\7��\�_0Gi�ǕO�R\f0�X��*����Q�`�.�v��#����)�w����
o�h����*,w9�[��µ=�'x�]����{e�8}�6!������)*�+0:6RD�I<[��;;�]۝�o�@����������<�
���s�sP֗��rls8*9\ܭ�T�ފ��P�s88K!�B�\��T����.�t�<��\}�"W�$P��P�k�|��}���������cff$�,Y�\?g������ �B�r�dv�܁�s��g"������� �C��Ν;����'s&G�M�?5��)������?/��&�;���PRT�IvamP�����N�Ay�k6�yr�N�K�n�,����By�����%Δ�t���3SHn"sI769bø�����%����_�m�;��um�	ĳ��G�� �umO)6�o��S �Bf��c��w���{�\�º�;��vm[���rii�8��`�Z޺��I����)�	C��K
�d�A��h{$6�'��.�^��ec��B!�2�i�� �n�&Ib{cy=��/I;`� ��s�o�����I�Yֺd~S_W�������B	���f&�P]U�����˲+(pW�0w'��#̬1���,s>��ۖ��L��\��=��=> &�k(Ƶ'\��
�Y��l�E�U�GQ�/DJ���,��]'��چ��a\�z$���ա�:�<��k��L��̸�����k����n�k_Q�W\\������B�l�����;����C��:��rm��l9�#Lh�\ۣ��p�*�E�7n���@rG__�_��-[�d\؞��Z�*�se�U��i��KZ�b��i1�c!�B!s�%�Ә�;����˛����K�74���>N��a.ȶ�^�5�+���󍋛A�7�nڂ���!�2[Ν=�W���8
2iY���źI�b%,k.���A1�pu1�NsJc,٣Ȧ�i��V~��U3����Y�dz�K	x;1���6H���ra�Ǩ�R� /\���@rK�6��":w�!� 1��Z��5�2����"/���M׵QwY�\�]mפm����v��'=�c�mj_�3'��N!$}Μ9�w���.p���*�k{�����7�r9�|_pI&sߗʬ����Z�ny�d�J�H�{�Όg������qΝ��z�c[[�e��k�U][֒�U������ 	 � ��׍" &H"���'�tm�~��5�#���l�0���.)-���/���rJ2���4 �
Ύ�	w      ����1���5��V��M�:h��U�1w��Y��1�{�.�����s�[�1H/K��fk+2�<   �	�x��O�ss��{�Ԓ��h��*m>A :677icc��\����냜#���[}m]w���ۨ��ܡ�C�1�sQc����@������U�Q���l	�v�>f�>�A)պ������KmW�ڵ]��*;�ѹ���&��� ]����+*�v[K��;��j;K�>��S�Z��CL  �ش[Ϟn���4�W&յ�G�(�^���l�.]�L����1w�ܑ�G��FpA+G�C�������fpS��˥�Nfi�N      ��||�pm7�*c,�����Gq���+�'(�$�8���m��_�@ �|��w���v   ��՗_ҟ����/��������G�Gݼy�._�I�0�w����Cr�j��q#���ꬹk�ża����X@�0��Y�T�T,[�R;���g8�B�H��I��=(nܸA Z�f�i�����ۅ�B�p�!����vm']R�g8��k�u�<)�y)��y�qm�{um��W�;�$kV���H���   ��y���&p�,�n��X�k����۱}J]��=f�Yz���t�k��G	�n�M�Ȧg$#�,�)/ Q\��@��O/�d��'�2���      ����,��J4:Zt$�U}��M����e��Z�k�E�9�۷o��\>GK�+����2m�x��%   �c�m����"���&�NV��Z��FFAQ���_���<�y@�(��4�9����{۴��:��쏢������tR����si�y��GX�.Z�"f��w�Q�JA����7�|C Z.u�"	Ƶ]":���ڮS��=��i�]��:yI[����yj\�9�]j�ݶo�?�+P��L���   ��{��1�./���������P(������U�wo�����>��=b޽{G�=�k׮%F�V�L��*��W^|"�ZP�����2?R#      �p��\��(��ɸ�5r�FR�0���24�A��$c��^�ӗ_~I ZV��Q6�%�^>��1����/   ��믿�?��O�ۿ$�N�1���
m��$�?���t}�s��:1_��yV�vŜ�)v��3y��7���W�tc�C�f~�JՌ<P�tbp�0xsb0�ZeE�>+6-D�ѳva݇k�f^�6�v���*yK/�!���]��W���A�]�ڮwD�_�N����&    hX�����v�U���	�}?J���z���{<�k�ȅK)�˵�A4��ͭ[�Z���*��~�ٮ���pI�J�+�7� �����B���W�       ��b�F��1�,�����U��|��ܡ>@�A7>|Ho߾%-k�H/���i��S��  �����--/-ӛ�o�����!p������ܤ��{�Ǐ[��uC���=����}za�L;�g[Z���56p��H�jB�Ze�}qI���*I�J��GPJ�ݻw�Y�����.�;�����E��e�Q2\�e��"u��c?y���:ϐ\���s�����@Ф0Z���	�J%   ���~{�-�����~�LRO%BA���p�U~(�FFF�ҕ���ۇ��M����׎�8�I�c��Z*!X%�J!&(�A�����j� p     `8m���HfK��Rc,�C�z��Y�ۇ	��d�[���]������������-   As��M��_�������3Y_������7n���z�s}��ݍ~ukQ*'���w� v��]�f~.j����@�0�#����R�2�/r�p�NE��̆��B��F�i���ٵ�YF���\�me�g=;�S��pm���2�M�m�=���F��?�F���N   @X�������;ؗ�O�k;��cG>q�ޗ�ݷk��Vytm���!p��/��"�v��U��_��{�s�i�fF3��       �p���f}V.ҙ��ܡڵ���\�3L��U���D�����a���.ғ��   vϷ����VVi����Q���y��~G :�ܹC?����>�9B�u6%��KiPM.}|!_��)
����qs��@� sc:+��h��ف!�u��]�.e?��>�A)q]�Z�o���@�8���]\�5aC�p�������*�����$�#���|�rm7�U�ݵ���k� ʷ�ۤvm7ʊ�︣�C*��   ������\�cgo�,É�O��wmo��X7Z�v��W�#-�_���O��{�E��G��`�)���U2�H�@����$���{��rw      ����zB�¨ÙM9Vҷ�'o��k�Н=���	D��:�����KW����   �oݦ����{�a.��G�W_}e{�=�u�:�*a}k]w���-������?g�e�h�R>;G�:f,`@� Wg��9�8�nIm� �07��'�qu�Ş�$`Ÿ{�.��l6KK++�
a�Ñ�t����\��V��n�������by]&�'��ڮ�+]۹6���ѹ����k�y>
Q����ý  @$0���_3�tm�P��ޠ���u���iii�޾}K ����͛t�ʕH�I����x��,Xe����Un�*����^/!n     `�x>Kک&up�������=��:.yC~�0���A/_�$-��k���WޣG�%    l^>{N�����&������5���M�������n�k�>W���i�
v�/	�y>7���b��N������*�e�X�Fə�vso�.NE��!z�P�0xN��$v����s$�ϭ��T���2޵ݢ}�J���µ](s��5ތ���9���e}��;�Ѝ6��ٗk��}��]!�'�����n�`���U*   ��i��<5?G�GF�v����x��k�X��G� p��H��wPo+�]��N��_�q�nY �E��pp/��
      ��u�7�Upp���(� ��"�ża��C�0IW��c��7����)���$�N.�������   6L����'�����Y�ӓ�P���o��������煵�!
��~6׷�b���g�����l}�A�1aA�dT?��$Q-
�m�3� T�d�QO�r����u���'-�/�/��\�;bj��;�vN�m�͵]s��ޮ \��gb�Z}~�^]ۭ���O����   D�7_C�����]���%X�k�����{٣���W�_��	Dǭ[�(�z$�>v���Ry]d+1f�(�      �tF%n�qޙ���[����Y�Bخ@���u�~'�Y=�N ��.����  D���-��ӻ��ce�=y�@4�>3�bwٺ�ԃ�a�!t7���n�<��<�`�=�eƳY�J�t$�f�pJ�R�Y�r�n���V���۷	D��yn�A_���69�����K��5-b�v�y���.�]��&n玧rm7^��ۚu]    D�m�~C���+�P�pm��\��W�x�v��s�T���)�h`B���=���k����P���s�5��K��:	�UN��`389:�b~�J�      ��r$��w5����pM��T���FEzn'���s���^�{;  �H�q���c��_�+�����{԰��gnQP?}k�i���.�k���xs�
��`� �11��ӓc*FM�����S��r���wb�+j���y��-={��@tL�����D[�ΐ���l[�]�ퟑN�(]��N�s��vᵣ��;�g�n��F���W蛯�&    j~����O���>n+��*vI\�{�M�������X����W�֍���M7x�����X���un�8.K!X%۷l`����F��,k>gw���e���     FrDǇGT(ly@/b�L��rڵ��'�u=�upp�����/.H�SS����V   @�`�X��3��#�����f��\���7oR�T���g���i~嶎=o���2M�}lo�ϼ�d����!e�i��^��xo.KT��=N-(���e|��QGZ�	}�V̽?ZѲva�ŵ].��<#�3Q�-sm�
�%��g��zv%�Y�k��L�^(�.o=������vvsm��>96Ao޼!    j*�
��:y��E���6�*��v�{����@�!�o���Ö�}���y��b�ʪ�ra0�WR���%n���x�0?      ���y�3�&�e}ǒQ�=�tI��7�8�l�6�#��X^]i]� }��w?���&    j������1�귿!�.X�xay�޼�"����Ağ~�ib�a�i.�w������7�H���x��7�ժ�>��g{5J;���X�2�tDE7�v?Ir��~�,1�������V��ѣG�eem͗��.��	މ����J�tm��9�w����@�z+]ۅ���ڮ��a�����.�ӟk�f+�����[�tne��}��   ���կ~E�ӟ��W/�|ֽօk��vY�J��W��%�r��}iy�
a�k�3�|�{\���qc(f��=g	      0���5(Sq�ޔ�����_��;��<�@�0z��&H###T=�P�Z%    j؀ƑL��Uk�v�	�{t�>߃Z���h�Xe�v��\��]�k<�a�ͱZK�.N=ۣ��{@Ld*t&qa�%��1�~8$+Is]�e���w��&�XZ^�ܿ�?
�t�Y�k���BpI� \��7W`�uum'�c�ǵ���� ^�v�h��v���)v7��|X[^����s   �����z�)BUjأqm�R�&�v�drj�5����;�p�֭�4��	��z8p���-�l��A+bv٣����t��      |&�:�2Μ!g�e�7��)�~��.�c�^��"���U�T�Ax@��N~��ߡ����   �����/���|����5�t���J����=J(Q��?2�����_��g|�b���23�<�"[?��
����H%���
�8V�Z���0>>N��F���bb�������'&'���'����J��tG%�{�C��s:����U\��muy[�˩T*�
w����r@��c��
��޿}۶�׶��)_q鈴�fѻ�o���[.�9-�كG����ȓ���b�����666b96��b.l�8`�ξ?�r�988��/��f� �s����z���%�<w�Y;>>n}�����,Bq��0������WZ];GG'���k�}描�iow������n�����׿QU��Wi�����?��g�������I�c��7[��ޱl���y:;-)����>	�W�k�؀��ϟ��˗)i�j�i���d�'���O_���)�n��     �a [/9��]��r�^ך9C����X$�u�Dސ=�m˿����������*d�   ,9;5Cc,0�L��Pq�H%��!f�œ��q�W������wM�y�.�XBܠ�3�S����Ѳ�MuQ��xa�]��p\�$O��q
�ezA&nBp�\�%�k��㡗s��;��kJt�V/w���V��ާ>�f�S��˅��3݋�{�N�޶��KK�!� ��`~�\\��2����ߺM׿�qOm'�L�vѵ�lS�՝�7��O?q�ǥ��ɧ���?�ҥK��_����Y*���}��i���+L���K캋&P�p���������~�صq�{����ަ������K�����y����c9>�?ZXX�mpA����~�3z��R�noo�^o��k]�
CpmW����~M���O?��������G]��i�W�v&l�V*�~�|׺�{��i���}{��wR�$�I�^�u�Ν�g9)
a˸X�|�K�"v�"���׬83����      ���5�����`�s�B�6!��H�~��I���/_����݁4�byC�������Y�}��㾎ͮՃݽ�qB��������&���~{�^��%�Jg��[YZ�������cai6bF-����ۋ��)7gb�`�{7�<w�=�οR��r|f�=��L�0����!�g���o��Fǋ���#]_f�`���	g���;ψ�>�trJ#{�{�p�og��}�}��8������O�Ȼ����X_������ܢ���JX�[��i�`s�7$י�������ww�`���~�����$�[��Ī�lSߑI
t�u���#-���)��v��&�G-q��K���n����le�<�.�_gs�vv�8'ׅ�:�t��T}������u+����O�5�+��A�N����v�$/�s�0BǇG�   ������u�۷�*��Wq{�"�~�*E�rex_u�ܫ+{��Q0/����Y`X�D÷�~�P"2h���d�2����.V���7�%x��_�����     d&F2tvvJ�¨ҽ��b�7��V%һ%=T	�8�l�v����%<3�&q����'�&1;����O��{�)�l��əi�˨��c���{��\:���ZY_�ݿ�����������l�̙�w���t,�O�{���[���h4�A��L̜��|����&����6�{��=��e�(�~o�ʰ����~�/�$]���ۺg&Jq��|���~������D8�X�����k����Y�gtt��IX�����7oҏ���ԃF���tx.��_�_��N�(���Z�ӆ����,ig�R�pbp��_�H7q|p������K�?�o�[aB���y���S�����z|G���ќ\�����\ŵ��;��~��׵����l�̶K���������+   ���{�飏�c
�u��]R�k{�����O��݇`ݯk;O~$Ok����]F������_�����+c`hkQ��O����sA�\Ly�
     �!��l���j�;���`$���E�~���$�(o���>|H :ص���L ]\X[��O7   H
L伲�L�߾!��ϭ���{��QK����:��|?�S(7�r���>�[�0c�
�FC��39z�[�4�{ ,�5/����&f'م�t��	����v'ɑ�<x@ :V��Z�uQ4�ݵ�+ٵ�*K�k;;�����ǵ��.��C|O���v�l����	   H
�w��`���lkZGgYQ�\�Uu�ڮ��ӕ�߃�=B���9�
�� B
�q�;��K+X�}��՟��� ��]��ևP      ���8Q�"IP�^�}M����n%)��Z�@m����<�;�� =\����?��   ��p��]�џ��)c�Xl9�����N3IWA�=���m����1@��K<7I�x�R��0��RY��V&�� �p!���F�I}A���?B����g]�\��=b�W��7K�lI�V�ڶ�%�Bpm�I�F.1D���;��Ѻ]D�>��@�o��smw�ݕ�S�ŅEz��	   I㷟��~��?��/�BkĚ����zw�v���k����k�6��ɓ't���X�M`�.�.x������28��\�����Ϛ��       ��2��PYq��g��D�����[�H� ��	·�~K :�ޞ:
#*��7{  �t�~��F��Uk�v9N�~��`���Z6�m�N���������};�ny���"���s�|�l�Ni� ��N�#)$�v��])d�vl�[�j����8������trrB :�W�h�Kx̮���	bpI��W��ծ�z]ۮq��}����v�\Ϗ�~���/��   ��qxxh��k{�mRW���G����γ���
�����G��0���k�"�{[4�0n�>ޏ��[_����      6�z��.�X�����FWlyC�[�3�<�<{��vvvD����t��w>��7n   �4n~s�>����~���}t�Q���+z��5������仺�v�A�.�Zy?�_�_�=.3�*P���= �g�����<\�F��{8J�`�8�c�A&�����)���ܜ]��~D�my�].��zе]V�һ;����.�D)��e�trt��  ���f�_^���ǺH]���'\ۻ�����rt��:��xF X�KF\�a��bǥ�!`%�M���1 	T�J%�-fh��       �`R-[����ۭ���!u��G�7t#���G�D��-.H�ctttD   @���ۣߙ�&�.0�2RX���Çt�ܹ�ЃA<.{.�{�}n���=oH�~~/9�F�� p}1Y�P�D�¨�sV��y��6�뼻�>ѮX�"��
~����A :Vέ��iF��R��,P��N;,wQ��vm�� �k��
ܵ��&��^x����+��W�}N   @R�}�����M�K������z���um燐W�vq�/]��=Bz$�]�?�н�W���u��ޏ7�I�������Y�     P&FX��7s�lI�]s�N����`�����SD�0Zf��(��H�VWi��   �ʻ�oiq~��w�H�B��f��p��@4����&�ܢ����j��7���F<���r�y��8m�{�\���r�(!9-wR�3�C�ca�1_G0�%)�~���cyu���S୓�ƞl�vN
�ѵ��_O��ƶѹ��$>�4� ���x�
����'    ��{ȓ�c�f�T��S�ڮ��k;+����.k�������ݻ�h4Z�3F�"t���e����b]Y�ݳ�]�b��X��T      8g2De�֌���<�=oh�5��$�y���pp��e��kWާ��/   H*�oݦ��G�����})�����ci���_u۷���~�V|Q=@]�74���z��w�昵��L����(�@��'�E�2g��v���.X�*X%�u��v'9����9+t;.��	��ݻG :�W�5�F�\�ۓP�k��пk�D��E��j�Y�h�M��l�_�v���ֱ����E��    ������O~����զ�<M��A�߫�=.�v�peu���g�k>;;;���I.\�k?�����[�N�ʵo�$-��/V	q�n4Si�3K      ��ce�(S�8���.$�ct�
K�,¼ar��9��cai�@z`n��r9��;   ��7�4c,������A�k���
^�.�{;�{�*�L&#5��d4Z� z�K��>��T�"��������*��#2%����W^�xA��)��FL.��مYA�ݫk�U.�׵�o[��X i{�v*]ۉ���v��wm7�.�[�����A   @���ۣ������ۄk���ǣ��������iu�m�xI |�ߍ͞u�����н�M�ݶU��ߺ؏Q#���מ�,��=�(7�5F      ��c*[��b@�J�Nʁ�Z��!��G��k{_�~�Z@4�����ӏ>��7n   �tn5�>��ݺw�@:�}i�lll���>���v�;�W���uD��(u���r}xO�wS�������3 p�|�LUc$���5�\�|��;N��8�$�.�Ӧ`�x�,�,S6c�j�rmw:����g쇀<:���.i�]��k�M��9�n�;��rm'��]�vM5�|�u���c�Ѭ��\Q  /�=�əI:<:�L��R[���z~�&յ�������\�t�y��i(�MJ��ؕ�R5{�]��|^pue�/��)A�     �`�m�)���Ͱ��9��P���t�vٺ���#o!ӳ3-Go��'�����   ���f�����.��P+�����Z��2���?��XD�n�[��c��˻�;�󆤈���eTg3?�PZ���OՒ}zq�E�-P�p�a߾{8*�	�?N :VVW�c�M�]ۉT"x�_�f:�;���.m�\��ݵ�lm��K�v�#��dmĵ]����6���:��_�[7n   0(ܼy����˖��Q��֕{�]a��˵�����[�[[#�=��'E��q�q)#`��������������ͥtrBYm��z�@      @4*%3O�O+޵O��d}�ֳ.yCUB�%��W�� ��d����Ez��   {;;4=5M�������G3�b�^��"{.�j�E�ۋ}z����z�+��~F���9+��ܭ�M3h\��Hp;.lV%?�Z�낌�����E��ڮ~�t-b�vG[a{H��r��؆(\�ݏe������m   6R�Z�t��k�TD�"�v��vym��v~�������ȎW�ʀױ���µ(���7���q�%.� yv��S9zyP'      �`qvzB�\�S�Ж7�&�53?��uI��7L�@y�hYX\$��]��~��&   `P�}�6��������������x�@4<y"��"P�|�P�R�W���k�@6`�R:i�a��
�}�8��Z�J�Q��*Ub[��e!��[$!������-�bj��D���QF�z�M��Y*Z���{pm��%�]�]�n����9�˵]R��&����G������  O����"���I�õ]Z�����˵��M585=E����ٳgtxxH��ӭ׃���q���f�4e}�â]��݉�-���     0Zy�Z����G�vU�[���@uސl���&!o�P�<�ava�@z�6�H�u�'   �J�
�<��0��@ :�`���"C���l�?+���\�^��۫��,�X*�hb$CǕ�����d�����R�0��2:"�.�p���u���Ar]�� �gfh�P��ӵ�#��T��=��i�߮�܏k�ޏk������pm���{-m�b�3��-sls��y�s�6   �ƽ���?~�!m<۰�G���,�O�]���jT��Ы��v����t�&�[���3�������	��lɷ7��;/5s����jv
���zݝ2�e���       ���T�޾d�����������$�����ڦ��c��� ��Q�'������-   ���=������]����4�G�T�T	��Ç�I:z�$
ԃ6�jI���˩���5s��$[a���hm:C�ә;�������T2��u���]b�cX�)�gA�j?HQ���Lm15	�i"C���:��pkm�Yd���(k�`�����W�����g�͵����\�e?{��G�i{{�   �A��՚i�0��pm�ϵ]��z�����˖�]�p��ۅ�f��gQ6���B*T�eX�7C      ��a���k�9��'�ż�8x�y�a��&�7,���a~�i����_��   w�ܡ?����	f�I�4;?Oo�^6��W�����}�g�r�����������zM��*N�q�2�4F��	�}0��SU�𸋋�T�t������#`�6>D͠9�3��".��4����ݵ]�Փ��w�	e��U�����f\!���m�S .�Ώk�c_Q��P{Y��]�$�A�|�N��   T?~BS�S�z�u߂u�u�9���ۧ��c�umW�Ӈ��Gq���*����܌��Q��)�\X��b���su:Z�K��E      �\��}�gQ�������C�P�7�Ǡ�ٺ/^ o!s��҃��l1c   `�`���,$�ibn��0�/]�40�ޏk7�2��BT�o����>�y��\z���m�#T����5P%�P�\�m���"�@,Kb����D��Ғ��[��nWP��|n�K�ڮs۵7�����,>���\��O�ц~]�e�v�����t�"���   ��������O<�ǵ�O��]��{�7"<�v���>���K��f�d���O�J��]��x����_��/��Te2��^)�      #�2�$��]�>�<�yC��}��q�N3s������s��%>_   ��w�hzj�a��
0�P���KNnQ�S''���I5��ݖ;���k��_
��9�R�t�uPT����`�i���%�ݮ�pe���3<H�l��l.G3�ӝWy����������ؕ�f=��Ei��Vc���)����k��NB�*v��� �:�NSܮ�������drtu�e��f�+����   �J�ѠZ�ҵ^8��5�µ=�=�W]ZY�-$�#�ɓ'�׃��}{��]Ӭ��B=Мwb 3P%� �.g����Y��       H<z��I��o�ж�|��yP��ٳg��]s������G���?   0�ܻ{�Ο;Gw�}@`�a� :�LZ2�#P�︖�O��X���m�~��]>P��.[;k�e���}P*7/$�*2.T�]��}v�@)�Q�6KZ��WDa�ťE�d�d(�"o�;��������!��J�v�#ng�I����v�\�.��mm��i����k�}��Nz��3v*w���I���#tt�Q�   ��_����r}8������ܫ+{��k�������k�G��ũ���u����2T�:�A��]�H� d{6;��D�^a�      6P��U"�9C�AL�LS~$O %4���   0�T�U�e!�L��Q�����cᣚ��W��[�4Iʚ�+���)� x7����R9;!܁/f�Y��+T,���[�@V��^7�sJ�#���	�#d~a��$0�v��,�ε�cۉ�#k;�//��f�mD�fەu�cyqm�vJ���x�\�H_}�9   �Kj����r��+w�nR\�E��	D�`�'�|K)L�v�:1.Վ5��!�Px!�!T1�+|}���d��dw      ��b�*�*�9�#:���i��
�ffn�@:8���2   ���=����:�w�
��m�hx��!�j5���`�(P���jQ�7S,��-. ۟�C,�JT�iT�����Y�ʐv�=0e<��0
C6bC�����0	�^a�v&� �0�0'\_N9Q���Q �	�Cqm��k;/.w�������~;E�����   0�{�Z��(󺭼\Z걞�nH���� ����b3��x��yK�"����1�gF�����oT��,b@,����     ���>�E��Ǿ�8.�m�\.���y����K�闿�G   ��Ϟ�'��)mla6�4037K/6����C��ڢ.���A�-�D�$�[u�}{��\�E�.�X���n���=2W�)S񗜶9�u�#��1/R늷���oP(��,P�񁝹���3��g�v�5qs�L�-���xsm'y�I��h�F1��s;��ڮُ���d2tV:%   `X��ݥ+^��f��+pm�����%n�Qp???O�l��u8\G��f8�d97؅�f_��������pE�C��H�       ���(�f���#o��q�@l���	�@:�kj40�  ���~ϲZ�@:��jt���Y����!Pb߬���4��A隽o���d2�L=ޥ��{�L�4;u�G�g���Q�ū�h8V�� ��#��ׯ	D=O�L�J�ݛk���[7kr"m�����zDζk��л�m����7A�v���u��A�_�?���
=z��   �a�իW��s��C�����[�
���˫�>������}��@���a�+D���L��bԕ��{�X�ZG�"��:��l�       �g"_��Ϝ!����˗�czf���3?7G��m   0,���hrb����7�GK?�X��[��c�}p�/���u��@w2��~̱24�O� T�{�@U�h������ �vq�#5��L�;6p��
F��o6��6�`&��z�2�s�3��,�L� ����ڮn�L��ŵ�!n��.���bqm����߾�7   ��Z�Fz���jx����um�S7�v�zn���������{D-H�s�$����|��׉{.]2����+�;      ������n}�v!�}웙�h�����H���������g�   0,<�ؠ��O�_n
��4Z,�Y�D |T:�$��z۷ l�N�]��K��{��O��N�7��V'�p�?�@��#9�JU��$�@[�����~����i��aN+�����K��Ե]!�����Z��&'�õ��v��v�ޝoCԮ���=Q����Q�Z��   ���c�f�T���ٵ]�PO��@\�����[,���-�A |666�ڼwi��]���R����vW��U������~�/0��V=k�N       �d����GbyC op�L����e   ��R�D�㈳����Y�z	�{�2�8.�{/������~"��u��]�.�sČ�
�6 p��vfKB��u��dImQȫ�0�D��}��������?N ��;�:Rn�k�W�s�ۮ�s/�k�ŵ�&��ӵ�s��bq�2�v"i�bwj��]������ŵ]<�񾍏��λ   ��{w��ǿ�)m�~m+ϵ]R
�vO�Tu��KK��������imm����s��$,�H�Vq��`�����rvz�|��f�      $�z��U��=oh�)�7�o6�ߋ/D������T+   ��ѠL&C��#nff��3=E�q�y�$�_�z\�X��5�����(h7�|���Yy�D��x�rVrMD3D76���l�N<�2!`�g�F]���-1��v�*`�vC�M�2޵�] ޏk�&�N�v��P~��]۹#+�Wtm�&n�ʺ����[�_�˿   0l�)��h����~]��ԍڵ�K=U]u[=��#���-�3A0w�s��%^�ľm"waq��U��X�ʥ���h_X�}����S�     H:,o�D3*�5����߼yC ����^�B�>"   `�x�t�ί�ӳ0Vvf0032؀㓓����Z7I��^���%�vu��9K�)tw���K��f~����{����T�tq���m\r^�<bB��gs���g_�̍D���\(��ium7��RGP�+�k�̧k�Cl���L�f   F*g�t�um�ֶ�\�=�S���v�C=U�z0R(����ku����n�0���7+s\���<���o܌��z� >C+�     �t�G4�T*T,�[�7v�,o��ؙ���=�..Ӄ�w   6�={F?�� pO�s3��Z�ҫW��>��_/�64�|ܾ����f=���%�����N)��TO�������d���P]`D$<�A*�%�y��2IN����ׄ0�̈́A����&�㻝���8e�j�"!���7�v���7�"uQ��pm�0���ŵ�^o��j��m_���|t��S��"u[�I��aS��5�p���"��õ��@V���4O����~D'k�ݛǋ���{��繳ABq}���޳c�}�����ٱ�����7��\�� ���8���Ϩ01FG��B�d[*�E}����תUr#�v�_s�۷k����F�}��Jɵ]dna�޽y�}�2�nWX�x�sn�"͊^�ZdbT�D)�h�[��x>;
�      I�L���{��yC!�����}�~��@4
-�H4  `Ha��ls8 x�'&(��6
X�mss�%pw����_��҄��κ�Z���-oHB<������4����t���Kc�N��g��"�E<��'��������靤����[�A���ߧW��,���&�q;���)�x��V&
��m�ʚ�b޵�x���KOُ!ݝD�-)pEl��Q[�vx�O�9��q<�Q�|!�M�T��٥G�;���qzF�ǖH�0M�λzx�MNNѷ7����E�������v3y||�=L�W.�[#��������M��={�Y�5��
�<�����󑑑�oN�y��c�yq�γc��I��e�io߾�>��v�w�+}|�~J����1o߼�k�~���������޾�K0���.��P�^�}vo�g����U�0R��ޞ��U�.��}xTΎ��'����bF?߶�>�.��[&�po      �����'ޝ��{�yCqP,�ۭ�c���E���J\1T�s�������Ўͮ���i��p����;0f�����Yl�^�T�����O�OЍ������Ȏ��QO��,�:�qǔ%��]��}��g�+���B�y�,R*�b;�ql����8�{v���q�ާ�3��޹}�ʧ���#*���g���]L�g�,�7����ǚ���z�;/�{{C�������e�2x�E�9��p�����{i+�Ms,� yQ�̖���;Ӆi�.��´��N��ET�*��
�`#~NOO)H�{�>��~0��k�7N<n�~僫�އ��]������j�k�y����������ݵ�VOӅO��l������7��+�폓ҵ�ٮ^]��:�&����9��e?���w����d��O>��^�����������`�*���-��8`�����c96�������R,�g����u���{�:���gc�B5�s����3366F���?�sg�Y�4�����-,,�(��g�VL�o|�����������D쾕����~�S��]۝��r���;��t|՞�U��o��X��_[_�p�n��W/��������3��[�t��4�~�kj�^P��5aiו��+�kj�I�3u��      �b���c��x]��&R���8o��_AC��@�"��{lb��Lx�R�2-P��p=����1;�i����_:�=�6R���!?~�����q��yO�{o�"�y�����q�Ń����W��t��z��atǏ�w>����x��&��p� �{k�1I��Pͬf�/�ܢ�ҳ�4iRѩ�������|�;_G�O�I�u6���D�Au��nIj#H�����N*����X���^����K�0;;�zE�2���f�Qfsm7�qmS�-�1���gB"�fu5�Q&k��Z���m��u"idBr��$�Y?r�:��M���&n����6�T�Vy3   I�%��N,<
��"x?������'"�z����ա���Odn~�@40�;�b�ȓdw�^�W���uDq�:X�P�{�ә�T<D      ��ԩ&����H�'����F$�y��ϟ>c*s2�kV�o����}va��C6�9���*�NK4>5Ic1��ۍ��˥��߽�:���ޣ�Ϟ���hd�g�LOOOS\�y|#n�����3'if ��� �sg��l悸���দ�bsp��g�t&r�g>z����׮���w�?������L�����D��X3�s�s����pp���n���E�9X�E�Π�_�؇mˆ�~��O1���_�s�rog@��y�R���X�$`e<e�"w�rIoQ���[T���LZ0�m_/^� 3�3�6��mN���B�Q�M �ߵݱ/�k���l(߆ \�u������k;9��Vh�����)��@�N�=    ��g�ra�vv����wmW�k���Q�����������{�U vvvZ����Ůu��+E�
GgN��)��Ur���(����A�     @�ayC�K��Wn�ٶ��^��8 ֶV� (&cāh`�-�L�   ?�z���3=3C �6,NZn�-%���mP;_�ꟛ��5C�u����R�� �tI��u��mT�#%��f	Te�vˉ���`]�n��Nr0�딅'''�)-@�L�~�;�o-@�v~?*�� Ж���rm7��6D�ڮ�ֱ�o��������'   ;t���t�>\ˣ��k{߂����Gh�Ph�@�4z��-,,�*0�mZI��c��y��S���.�Z�	�!&       �d�e���q��.T�۝yC�����2��г��B[�^   0����������^p�lf-6;�1�[�.�����w�+G����r�bސ�+����y�d�4�\�����2Ή�(�/ޮ(V!}nM�0e�۷o9m�02>1N��QS	޹Z�x�[_��ߵ��Cǵ]"ZW�Br�%&��m7?NѸ�������sg�ѵ�:?vv����,}��o   ;�����U�ݟ�]V?R�v����}
��
A�.��=ө�������AP�0�V�l]s����ɬmV�b���x����D��c=D
      �?j���^�\��'�|����v黤8o�^�j5��F��������W���   �a���'t��З��^�&�)���R����o�O�C�s���]b��=�\K�to��g��3?)M@����Y�Q�R%��N�=�2����R%!��7oބz`137�k;9�um�H�.�!:�v~ �p�����	�H�o_���{�	��k���&   ��Պ�u�]ەM0�v���1Ѱ��@} ��blJ&t��Z�{�ʸ�w��f��K�0�]�E�vO�'      �T�ʔ�f��Xƣ����;�ud3@�����O���D���/�@!7�r�   �6�Dq��p��Hl�&�?��ڢ���ĘW���/�$�vY���
�X��!�4~`>
��r����'���:x##���,H�)pqb\�T*n���IF����G ���;�'w���~]��u����~��{um'�ߢ�]-R�	�[?|����nP�P��]�   3o߼���q:>9	ŵ]I�޿�<�v���꺝�1��w�ޅ�_=���΍��ҊHkk�6|__��2��]Öٱ,�b�*      I���Z3�es9ǀU�Y��A�D|��ڷל��_� o�095E �h  @���^*)���n�XI�����m"w5�Fg�n�%�%�W�~�r�[f�Ŗ�1%@�Ѭyqے������X�2هA���`�;;;�����	�Crm��J���۵��J��N!��q^-�]�Y����+�H�]?��d��G����   i��Ç��?�1�H�µ�뱒��η`��`S�� U��S+�]�Rv����A�|�S��;1�g
�     �T�3ds]ScY�B�@�7�	�S�7k�5p295I`�-����   i�tF��Q*���9M��A$�9�s��r�gc;�L�k��8Ck��B����c���O�Ƴ�ո�3ɓ�ݝ:��qg��F|�(C�*:����t��Џk{�����n����$
�em̵�l�µ]*��m��������O	   HGGG��e�R��{��_]?݁ \�yFG���7o���f�T���:}s׬];���*��C���w"�;      Ief�y�^�;�1�I�N��3���ʺ8����Z�5o�T����F�����fq~��>yB   @Z`�{�_���%0�����=*T������Ͼ�9D��z���ܡ3o���"�͏e pj���j���]l*�6��V�2+JV��ۭ���{P�ޘ���
ăpm�]��P�յ��/��֕�v��i��������.��rm��'������4�R�D   @���+�+��{=�/�}߂u�u�ۏ�(��P����|\lmm�?IP��Jˮ�x��0Es��֮',/)�B�     @R�.4��+vc,�l�g���]���l�לagI0Ȋ#o���[�0��������O   @Z`��^��;�9#ܣ����`�-e��&M*�f~��yC�v6S,��,���j@��ɑ��̛��rY���27epJ���3X��=h p���q�Eꌨ\�u����T�n4�^f\ޢ�]���\����|��J�е��#�Q��  @�`.��|��ժc]�N�pm����{=���~���4����ׯ_������u�w����U"ws��H�&FL�z��`U;� �!��n�#Z��CU      I����IgA�.KP��^������ڍ1s��5q���;�~)���q8�?��    a��v��I�u&u���kn����|��*����iw����ĳč����mIl�A*պ������-�@>c��Ϗ�ir��rm�������2lr���vq_����gLW��]�p���n�K����N�յݠX��Y�F�  �.=|H}ﻴ�%@Csm��=���	˵]�:;7�{�����ŋcmG��y�S"?�]��q����(s}�iu��     �dR�4�ݱ�bsI�� ��;�<�ob�l��fz��$����o[�RA�0"F�E��!%f�߷V�   �6�:fr����y���?c��l6�z��U��Vi�5��7�����yC��\�n7��Z��4�^�O
Z���+tuq�'�5�zc���8��b���u���c���!>3�3���k��˵ݱ/_��6xi�b_��b{Tۅ��n�Y^\���}ZZZ"    M���4�}2ҟC�ڮ�
�l�nR\��z3�D�	D �L]�pa�T"Ҁ�!l������j����}68n]�%��      Hy�F�1���>��K�����.��+�����Ak�319I`�Y?�FO�?���Q   ���˗���J/67	/�0Ɗ �3<99�����u�,~w�[j���f~V�myCu��܂���V��� p�I��wS�ncOb��m�|e�m�R��~�{{�f����𙞙�<��~\�u�k;_��=7����Ե�YG(s��7��A4�}�]���Um�~�&�ƨT*   �6�=J�Vϵ]V�g]��{?W��lzz�@������n�:����$�+Y�S:�T�-��J��H      ��mԬ{x�'��O��i��yC��;�K_�[7J��!����	����<}s��   Rǋ/�~���9�S�G�u2����q��m�*rW���{���e��|�8���[�ȥG���3�L���w�ywpo?'�l2+I�4԰/��G��sb��q����� �m�k;2��3O��d���N⾽����	ǳ�K�-��V�'z�Q    LjoS��k{?�p�v]�g�aӏ[^�T"FL��C��enD���w+>``�͛�h��2      ��Vo���!���6��u�o���sW�O�,7��C0�:�����a&�e�y  �J��*�s�L;��(���w���ի�0������7�q�g+o(����F9�`q��|���L�9�yubhc�L5�B�j�7G��i_���m���#���a7��2�v���pm���\�M�w���2�z˵]�_IYK�b���"rm7D�e�j�   ��rvV�\6G����P�S��^(��Q���'n����31g������TB��:i�]��k�d�pbw.PU)�       �Ԫe�}�Ù]��n�l��=j�~�chk��i���7��h��'0�@�   ��gp���lTt��m~6-�µݹ�\+l���3?ט�==3?C��Z��z4�N.�v�4��Yg�����~?�I���@Ut�@�Z�.X�tm'��Q�v[|��K��:���n	Qt�v$�G�MR�z�v/m�(��R��   ��勗t��y�~�α��A�۽���\u�;>�{d�)�t�;@V�Kf��:�*Peݫk�x���ئSΦw/htRF�     ��Q��)#1�j?�r�\��&n�d��F��a�0Ɗ�����%�ɴ�   @Z��|f3^p?���_�����>le�6U�L�7Eiw��@s~�"n�<��Vr�O�*����񉎮H�S"�ٵ]D�"tm'��D$�۵]�˶�ͭ�"/��q{�6q��F���9���$    ��|������]A��k{�'��f��RE]YMi�Iq�H�\��5�Z6������V�n��[E�蕲/	TA*2��f]{�J6c{�0���2�m      �D.CT���PuTU��I�X�^��=g����-b�^���7�cp�f�����6   ie�y_9;3C�
C0����=2���"������� ��Frl���s��kYB�x4���"$R����ו�-�@UX�#P�v�@|8\۹�+�X�
޵��Nׄ2_��n�v��r�=�n�o~�   i�\.S&c����ڮn� ���+��ӵ]R455�
J�p�KM��6ʴ�RפS:gg��a�1�%,�p�1@��S`��#      H��l�Q�p6����mV*\ڇ���=Y&a����	��^�� ^έ��7���   ���js��]\��}����=*T���ͯ�B�*T�5g��ߙ�k�:��htRI�������Ӆ�=���`�9�ɦp��T%�m����86F�\�+q
����D�2�k;WOx���zw[���+�N�筝���nַ]���n�x�~\��c����k    R��ݏ�յ�_q� ���u�g�!p� 6�*��
~{~�h�D��b2��!l�����=p�\�x      ���"�p��y�}�tJq3�o����	Ⱥ6��v��ä�_�c�h-�R&�!0�������   ����+���'��|>O��<U+U႙���g~��ڟ�f~feS��T� p��T�y�4�y�t�:�)��T���QQ<r4�����!>����gN�z(��2q{d��rq�%V���+qmo�R&@?�����;�C}���u��   i���=���õ=q{���:Wsbj�@�looS�R���QFTZv�=q�8���8����o��o�:      ��D�y�^�f^����,��|���O�$��V*r����������#�    ݴĭ�v_[�����A��R�&{��Y��r����#�����c��Q�'��`�#A�]��
D��TVY��d���'�h�� �������=��KD�Ra;_dkC8���l������zsm'�����)\�%mj��1j   p�9{��tZ*�^�k��v�k;�����9::���cO��u`P�]�ޮ�8�,�z�`�,�0�m       Y������Q�ԃZ;6m�}�#�y��8��35}����̸`�H(�C�>�@�   �$
��0ּ�=܇�=l���R7��-��ʌ����KA���^�5�@�x��J@��u�A[�N��O��:ʰ���#�۷o	����d��h�qg������/�v�p}�]���"���   �v^�xA}�ݖ��_��JDޏ��o�vV��0���`�� |�����#� W������*:U�p���`�Hw      ��h��4�o����f�0�U��6� ��Y�)c��W������16>N`xay�ӓS   �N�Z�|.G�Z��pR�}m0}g�f~v�˶w��1 �-�`�5h��iw�欋̼H�ܕm��t�J������+ ��	É!��ο�z���+µ���ί'nwݦ�v���PG��nqqv���{�   ���:�86ޟ�9\��u��tmW�B)�o.�p�
э��pW�N�n��+��m�K�U�s.֐3�J      ��P�ڍ�x��^����/h�P'���+��!�� >�&��˹�U�z��   ���zk������M��f&�6����i*g~�*t��r]�|68Q�\�@�$ZS�{wpo��4��*[R��s��~��wmפ�r��y!���Nr'ٵݾ�ו����Nܱ'���ݻw   ��F��ZlD*"���o���������"������!P)]ܻٻ�����\p�Mܮpp�Q��      Y�5���;?PULL�5;�~K�P� ZM�7�q�����7b?�;�1�W���E��G   ����-��{߅�}�-��xa�m���Ѱ�w�g�Z�Ϯ�tup��XȦ�o��F2�K���GY��ic3�kk�H^�0������TED�8&��ڮqE6�v�흝��u܅��xum��-��k;�_�T�U    Q�w��k{���u#vm(���!*،[i��� n競�VĪ�`=��� f��@�     @��i������J�sי���FS$�%�H�	�888 5�l�!    M����(�{���(�Q��kI��9��I�X��ֿ���0�$17���=�?� ;�߁*S|��bN�U����T*�6b�6tC"v�����yumׅ��(�䡻��N'���tmw�����n߮3�E�7G��
b{r�Q*��|�4�u   @�z���\!y��KǊԉ�O�x\��6a
��`��^�=��+q���BA�.	�����      $��^wܿ��V���0�}�[ZPQ)�.R̯��
�Q(��	   ����h*��=:�`��:�b�(rW�����G��{�X�0Ki wd�nsTk?���@����TE�hK�����.��kB-R�	�ܵ����ڮ�_���   ��ĝ(�vy��tm��"*�v~E6����U��2ȁ*�y#&e���U��*���+b	�:n����      H�������A�>�~)5�B�0:�1b0�:    R�����8n��̳|�����f��-o��4��l}&E�s p�T1����c�M�#
�)`�v��]������]�S/��O�MH�y�;���(t�H���7I��]�5�u�9�   ��κؼ�)��;��ȣsm�'��n���"��T)����ciybL�j�s��vmK���&�Y�������      HZ�2���߭�b�Ј�;M�4IA܏t���ӏy�I
� ��F��>�@�   X�wq�����HKͦg�,nw��+o(�se|��=6X�0��t�ePp�ii	T����{40��\>'�����*n�^�Jq���.n���������}��!�wm7���l�Qr   @�x��]�z�N�$��pm�Y7^�vU���c���{�Q	K`/ƨ�AT���
w��=�`�����
�      $�F�b&�����;$�:�DY�Q�c��ݹ�7���h!��A�
*��	    m�ad&��FƑ�H.�k-�f��~�kq�g���l٬���5����{,�����sMC���^��"e���&�m��|>�������l6� ��b��>|Dַ� �v<S`)Ĺ}��v�wg�=xh+SȦ��o��f/h�tpЪw����M%��\��vک���C��3�m�tyc\\�e������Sz��M��9m�z������*�J��1�<�j�J�r9��f&@���q��� ��z�y�q���e��q�;���8�o��z+I����١��#�q����U��w��t��ݞ�W�%O0a���;�>õ�g��tg���q�k���ޛ�I��g�/�̳���>���[rK�|���w����iw�[�ǲ{,�#�j��ե�+���Ȍ�8�	F�@�#H�A>_);3 @F1"��}����,�fξ̺�C6���?��;��q�˹Ee��p8����7���_���!d<�"      @��N;?��Hu��zᬼ�3���W%Ņ��6�.�9����}�\֙۷>�Ã   ���#���G�׿A=a.�,�	�E��s�M��r��`]U;4���y�:oȷ�O�� p��lqc��tO������lR��	2�M0��+Q뛉M\��oa�7n�ѣ?�@)$+�=I���I)��W,l��Z<���ӧ	Gt��\�SOc���x�v?(�{�����,�'T�	�}���z����Ŷu���O?�E_�{������Y td0���۷�L�y��M��zN�g�~��'}����z���յ��	}ٽ�w=)ux��wg�|ϳq[D�~\��ڙ�����}��[6�p�������w~�w���p%�����OON��gOu���]W��>�}r|LO�>�4VwxW�����^��w���������>|�������M\�-�(�Y���s�A>eL�=E�p��x���q����!�j�!      �g:+���aX/��In9g��t6�ڥ�,�-6���ަ�p��`0c ��������ܟ������~rx��5����N΂ݮ]prtl���8:��� ����췫��-=��\��7c���#1e�_�И����kg�yv�̐�,���}W�L._{��3�&W��������>o߿O������q������a�����X�~������k���%ɇˇ�﫸+R�s���z�͎���%�������������9�2A����$vpWݘ��hɁ*�q2i7?�_�@[�Sf0���*X���us�?�����7�)Ru�//)���_L�B<�/�:m���H�õ����:e{f/��P�u/��긄�]!$_���r��m�;�Qt�{A�׈kG�K�/=�����ݻ���AD8Ha"'���� �\����U�L��^{W������\�&\����fT�=����>o\�ۇ}�
к|����H���q������g[�� ������L������h{G���3f7��y��������8H4����:�n�z��Hro]����.�i�y^�v�p�Fܾj�e���i����;�]���6]M���      @�_σ�\<L2�b~���9!d7�&ʪ��(&L*[�Jx��]��p�.=���V�~��7��ӏ�o_��ݛ{Q\�6Lxe����?�3����qGe�����ٳg�
�����̙��������Ύ��8]^;X�{��=z���/_�7,����}���ݻw��������l�����~�?����|���W��{�����1��o����}k}3����F�"e�y��d��]ܣ2}���q�_�/�^�+����)@���ٌ%��7�|S����nX��+8A�l�%q�Gf��B=^����~�X/\��~j�X�n���ɣ����~��Jr�K�Ƶ��P�N*�����}e������"   �'ؙiIyZm���
���3�V�r�pm��s���I�@g�E5�
���E�"w�=�y^��k.D/��      P������O�$s��NɹAZ:\�$t7�ra����\����Ϯ�a   �,��>�?�yC;,3_�onQDm�ū�9=�p��7 �'cw��m��h&,yߞ�db�Y�̎��*��-*U�����ȹ@*/ZH��tmO
Г�<��~FQ���Ke)���9������]��O�S^����F�ΘM�   d����x����YaѮ�i��ڞU�l�v�n�7Uv`w��
�]SN�L�?�i�A�n0���ۅ����vgM      4��`�<?1v�I��_��>g('���椬ݙ�yC;�;!�����}   �t��Xk:=7��7�u����[��u�U��0�=e�7d����kN52�k �!��)u;�L7~�E,�M:1��?
vbX�@���9��	@���.�M�;b�Q�k� $�����.���J��Q����e��     �o���U]۵*v��+������ʇ�ט����&Փd`�K�'��xu�8fO�x^<A��;pp     �:lt��x^��3�5�k/>�����DE��?ߟL&��:]�    �0�PS��Ev`�X�`|]�՗Co��7Ê��۹8���6o�S��Ѱ�@�G�[$�c��7eRԮz.�L	N� �b[�_\\(�n�oϵ�Br&�D
A�\پ�k��<Ȟk{$�����?�6�   @����;� 9*�v�k�%X/ŵ]����H�ڀ�3����e֭���g����v��EU�굪�       �K�෗H2�P�?V/xU�N������bwg,�srrB�|  �9�   I<���L�V`�ټ���Dus�zq�X��;�tbɰ'��{�+z��m�pR] �lrND��v"��H\�V��H�^d��	�///	�O�� ��I��um���]���Ūk���^)R/��]#�O�rm��-|�gT   2�g��ߠ�I�cP1���������um��E�[P&��`8�:�L+ͬ=�<17��uΎ^\!��P���=      Ua�s=J�qIgE�O���H=P��0w��H��vC�� �w    	�kM���6`F���6fչE3q{��n�z��>�ƹ�TS,.o����,W p7d�+�����I�%��X
TUiBw{���e���D�Zq�,l�D�NH.���ޑ���vŻE8G���z=�um��^��t�   ����)���s�;\��ߵ����5F�Q���mbr���R�*���)�G���     @e�D�U�<�y݋�s������3�VӘ ���!(��k���/�ì    ���z��n�1ެ)�>Ʒ6`:O��s}�'n�ŪDQ/�����yCw �n��n��	Qn-�V)+,<$�e��n�^#sGB��/O+�V��5BvI�>���ubm{�풐��wm[ԞS���b�D	q���f�O���     28?�~�W�k�����!nw�ڮ�[����E"�E8�7C ���"����>/�;��,J     �����bWpE̞C��x����ԨJ3([�Y벃X@\��lmmqQ    �紵�Ig���%�ځi=�1���nf�Us�U�-�z��Q��;G�!��\��7�8Yn���W���� �i;t��V�� ;͵�����'���'�*A|)��A=Q��[v$�]ң�u���5��	�u��^'�7tm�w/
�766���   @�- S�Q��ڮm���i3�C>�����m�)3�e��ֽ칽b�<��'��ږv��x��      @�t[�|	{ ��Lɼ�j��dy6i՗�Uiw�4 p��*�eg{�X   �������{M���ln����2�E]�д��a��X<F�7\����^��i.p/̉�<�T�[�V�+����\����RYȭwmOuW'o!���u��1���K��<��|��E�9Iu���K*���    l��^��/���Zy\�]����"Z�����x<��#��x I���"��%��bt!p     �2������S������ �����t!�+ۛ��pL    �h{o�@=�$r ,��䪸��$�T���H��z�"q����3���k/V?�&N)��e���U�`_� ��E�E���Y$��k;�k.�v�pޞk�X�ͯ��������+L  ��ٌ�er2���4'q��pm״��k͒���O��{�X!Y��E�	���q��      *���RZΐ�G���&S�u�]��d��%ǹ�;���Lc,    	�~���>�z��4D\��yk]s�&g�(D���ý�v3�Ș�����
O�
Ik� ��{���:mYQ�L%�����.<��vw��i��������ڞ&��w�T   �@�n�ڮy��9�!n׾�>u:]�e�%p_�����\��
��EnR��b�ߦ      �A��Gۂ�����k�������zTU��=�1lW<PO666
   u��j���ԓv�X[TA��2�-c��?�_����o?tz�T8�Z$x�խ��ڎ\s���!L���	�x�v����r������4��I�{��|)�v�r��/?�������e�vA_   @���]du�v��]ە��uqm����VSq;N]l�m���5�b)4��H3 �a4c�����g[��6�      T��������T�+}�b*nϢ
�U�B��
,�T��`%��e>   ��a�u;]��wk�aޖ�[̓3̚Wy�~�/���e܁��݆�����|ERz�w�V��/O,�0>�E�����]�)w�um���ʶ]۽�v�sZ��]�P�k{t��%�)   >'po�k���������"�^�@�4z�f�J���C$�)�W?�      @shyB�c����K����z�1�
�%+�p���:po�7�%    @u��dmas�V��4?ły[Z.��M�5=e� y���t�f�������)�X��� [ʧ91Į��{i�v�q�F�v�@�N����v�S7wm׋�m�e
���/����u���ή0�v�3   @�l6�^ݵݼ��uӺ�]ۍ�I�f���<�]�@� P���y~R���!�     @eh]�ϧ�'t;?{&s�7�C�    4��:�ƹ3�J'k�V��˕G09Ts��ɝ�cu�TCZ|rY�h���Q�د��.Uv�;[.��j��\���R#���+�����q��k��J��TG8�?!\OI�b/��׵=!�   ��l%q;\�+�ڮ?�N[I�`�y�Z���A8?@�0�+��Қ      �CN<��{��9A��Oe�#�����    @��\�sǘR�N��u�-Ff׺���_�V�924�?�Ғo�7KB�jt�z���\;���c��ڵ]U��k{F�+��/Z�����t�,���ڮoW>&�k{���3    �!}O�ھ����v3q{���Δ��qm���nl�hNr�Aq���K�{�'     P!�8��:�񥌄�v�d}�����`�e�N�Z�#�    h��d�ic�k��tJu'�+� ��(M�/ĩF�D���]x�d��E�J�g,� )`�f+M�!+P��z�^t����5b�Rn��*��+�W���/�s"�\�iQ0_�k;�<a�   ���k�ڮ��޵}!!��Rq�cVp���� ģr��k��{y�      �J8���a����~�7���>w    -�'�ƹv���ݕ�ܧ���7��e ��	X���w����j�Jsm�R\�%��R��j���T�k;Ie�Ӣ�w����    J��ܕ��S�6=CL��󺪚帶�z�E���u=�E�|0o�F��NiE�Ųi�      nH찔7�'��6�n��ua��3    @�x��`�g;4:ohl�%�I�F�����.6�s�^C��D[GJ<����5H�H�A(a���=�H]S��?���I�r������uumW֡�\���|�#   @�j���k{ �^cq{^�vS������|����y�V�K��-6ҭ��U�     P�Ni��ZVN�@f���ÝYoW      �y[:iW�Д���⑿|��3.�nv xv`�Y���]��e��(��M]ۓ���,�v/���sm׉�^x�b_�k{R�ηS�k{�>bT   @*�Ʉ:�6M[�5Ƶ]�ĺ���k�O�>��Eշ�>��f'�dm�     �
��3P3V1�B����f     P?`�e�ۊE4�V����Z��!ѭ�%�j���s��}��m��l^�k;�(-�۹���%%w(l�_µ�����>�ye;庶׎�   �e6��_%��!�^]����B��d�qx�\�yZm�l�T��^-�[�r��     P��s���OJ'���m��Z<X`m�C<     �c�a�{�r��"h�!p<e"�zcV]@�@���\�M��Q�%�v�NX�.��-3���   �c:����pm�q^���pmO�� �0o��JK�1�     �2���sO)c���1p      ,&_Vh�-���I�����E�B+͸�!p7f�L2�U��C�k�v�-:��ھ����	�b�L�v�ڎoE�B����*��2���c?�b���+�����Q[r!    x�[p���k�Yai���4oXQw5�v�Nvhb���;˰!���      T�<��RWc6�����    @�h�0#��m��l/�O�F��8�t>�X�t�h��]�c��\�.�U�k{|J
���?}��k]�=�A!��T�k{,n'",   ��0���祮盾�e���`Km+ PU,�;`|     @u�R�˴c���6S�.ͩ0��vī9�+    z�=Yk<���y�Er�Ư/���]��g�V�]�k�T��ڞ��k{xNĻ�S�Kqm�����pm�1�   ��f>��#Sq{u]��륹��XP�k;_	Y;`a2      ��x� �M0���)��2    |O�*���F�O����!p7��Ce���̵Ԛk�,Ҷ���I='*��]�vV�+޵=)�O;'    Ȱ	���1Wwm/���L�^�v����R����VN6@�*/�     P��(�>Vh�ٲ��Z-�M�   �`�Yg�X����H���Mi��P��b���^�k{R�mѵ]�/�'i���Zյ]QV�k;��   ����攛d�µ}q{����r\�źH�١�n�      ��G$�&JX�uma�3    ��xX�l���Ҕ�� p7��Cu����ϾX��V�n��NI�5'$W���"ɑ<�k{xNJ�}R .��+�'յ],Ksm_�it�j���<n	�v��    5��۟LVvm�S��庶���w      @S�@?(�?� �����F��G   ��k��v���.M��A�n��1��}�@�n���ݡE��=N���k{�%=͵=)�����	ι:B_�t�'�NQ��r����.~�,��>_}�8   ��m�<�%��k�ھB�"\�5��>�"��g>U6���X2ߓ�     P0>�
柖@
��9a��    =��,��m���M wc��!$�*>/��v����[z�>X������y��>�L�g?���I-����5(R�ˇzRm���{�O��O?=�w��,J�K.8?;~�y�J(O��g��� ]כWo���cv[�z�L��.���c�bg��?.<}rr�(��`0���sg���驳k�����Ņ��ٵO�Sg�.����ap��\���]���w�}�~\�����}�M&'����{�._{�Y7��>oٿ�p|Eak�<��d���7�����r͕��s���o���n��n����k�����zZ�Z����ѿ��E��NNi{{�l������}^U��2)lJoؐX��*      ��vI�ņ�V`�&W���*;���wO_[���f`�ߘ��8�w'z���b�;��*�\����.�	�]���!� ���3����.m�m��!e}�5u�b��B�\L���.`_&����t�x�[;������k�S���#��k��~���;�ߨ��r����K\��/����E�U�um��?|N�'̟�b逮��}����}��	����+Ta��gϞ�޼yC�nݢ~���o���ٵ3�%�޻w�I�/^���O��+\�w����{��{.py����mmmY��v����۷���'��~���ܹ�lq��מ��������������Q��U�k;����~F��\�Y���wS����~�&�	=x�P8'�V����?��E��g����Ee����`n|��A�     ��0�rɘK�Źʎ3�\��n���C��l<�_��j���prt��%np>�������k��}����q` 2?.`F),�
f���5wi���w�?�ײ�+C6�A,�r�WWWN�g�;뻉�L���\��l��L��=wtt�Y��+�~��B�gc��_~M�p�����NzG�q6��ݟά��=�Ɩ^M�=�p����$�?9�Cl�fC򆸫�ܝ�d::M�R�Tܦ�+<�o@��7���䲰]/$_Ԏ=�>��ۓ�m�2~�\�u(QG8'��Rl??���^)$׉֥2_ѷ����e\;-\�)�^���	ۅ��#   @K��"6+L�nV�L����fuu��!n״iz^�^�vq���-(�C�ơ��K��f��      Tѥ'��;C��ĥ1V(4q%:�}��}��O�����o���޾|\��+��/�������S��_�u����������&v�裏��s�U�̜�����������w����>���M.pm�Ča=z���/_�7�.۸|��w,[\p��]'�7ِ-���_������������3c�*����[�f��;��X����湵�>˝mll�8v5?��9�HB�n�J+|�B����S�����^3um7�k\�=R	瓎��]�9��\'l���B�%��'������r���:    H��ti<��]]���*X7����Nʺ�\�՗5/�A%`WɈ��X��0P��0�     �:,3>��0]]
�m�     ��Hl�U�mkm�U���6���5�	��7�p3�Q��(�P)����lʜ-�tmWG��k�(�(ߵ]<�pݒk�J�_�k{�1    ��Zfߓ�\����uum'��*˵�o����n�u���?V��xF�#� ��=      �A;3Α�NoI����V�-b��f���Y     ����Z�{�'�b���!z�����ԃ<;�/pY���k�(ZW���K��S�Ϊ���1wm�w�+���'������4�   � �{����f�;��\ۥ�q0ٲ�m�ķ�/�J������       G�q\C���������   �L���09�D
0�>�#T���		��e�q~Z-����7R�l�0�*;��W���wm���C�rٍ0�I~i�vE^Y��+]�5.��)��
��
���9)�Ay    (��E�smW>������0\Wעk���ނk;_w2(��*gcނ���Z���      �Qχ����G�ik[A��0�aG�Z��!    ��q�=o3��/gl������k�,g��Sz|K'�?Y�B�k��xBŹ�3�O��.	�=OZ@dٵ]hWю�k��^�k;	�H|���Ν7�G   �������3���ZŻ�ӏ����ڮ(]O�q.(���������ߓ�Bz��     ����}2�:$���`�,�;�0�N	Ԙ&�   �e�x��L1εB��������7v����=��C�n�LvL�U�N���:eͳ���@��%P>㫫x�fŵ}Ѩ�	[��Ȯ�|��]�e�k{� >Y�_.��k{Z���Z�y    Ĵ��I��++j���}�z��tuM��Tw2�������z��{�틇p�^��Gm�k��     P3���9���s��C�R��"����?5a    4���\T]�^Dnr�i�<���9uÜa�c������!�@���UR&7xx��Y�ދ� p�T�>۟�e&$_ŵ=<�+[Ƶ�?Gc�v��X�k�HP��vR|�*�a�V�   Z<o�=��k��0���"\�M��Uwm���ʧ��0'{�/�3$����     �����)Ɣc)51X��!yC;La      j�t�q�ʞ�U�<+3�g�?�:������	���{���ү��Upi�P��Ɍ:�Va����K~�z��3]�I�Zn���yU_tK����*�rmO�7���۵�{�Ն�   ��j��yWum��4���k�I��u�]۵���w+4z�f���ew�<�YE}�<      T6>���YJ,�������ք�s�=��0��e��W    ��k�������%�̮3��ɔbv~q�"���!��;bSQ��Lb�&���mHuh=)"����	�a2�P�;�((׵=n[)nW�ծ�|l�ڞ!Z��ڞ���������2S����Uuf3?<\]]    DB�,�ھ>��|]l�m������`� ��ח��!�     @e�r��,S,��s����S�r�=%� gK     PG�7�Cּ������+�Қ�)v���x=	wc���@�N,��Z'���[�*r_�a���A������.ѵ]�6/���ڞ}>*��T���]ۃ�|^�"]ۥ@��j|E����   
�&�pm/I�_�k��x����T>Х�p��ȡ*��|��=!�0gF       �L���m� �fMZ�	�?&��f���Q�V�`�-   �D�Ŗ��l6~@��a޶jn2���Y9q�� g(�9n�m��!WS?vXX������aC�[���L&I!����	q���8��F���ڮ�K���Ο�ޑ��v��j<���:::"    ĴZ���Utmן�y�����L��A�|�U���H�[^�M�     `���@�sR��!���3����s��L�v�?Y�3��LgSj��p0   $677�rxI��`�c�*����M���l.��F>s�gn�;�5#��!���P�xnm���U
9�
�1�{n� ��ڞ&n�]ۥ::���̢Cu������w�X�F���FW#���%    ��NF��'pm_7�v�Jv��E��=D��{{҉!vl�)�=��=0�     ����z��H��}��C�_U��a�i��dB-�޵d0q���S   @�~\\�'l|�P��q3̳�x@"�(�T��L��UC���2��D�>����fl�q@h!6*�2�A0��t:4��b�LBqWp;%]�����e�UD6]��c�'�'�q�Lҵ]��ʮ���O��pD�;;    ����`!O1��\�>�$�v�C����9i��k{�Z]��ءW'���M��u�D)�Nʭ����X�     @e�L�s	>o�\�k�+ա�dU�<;�����d2����>(����   ����w+�y[hh�DLf�������������b��UC<� p7d8���Z܍��N��B���(����`aۣ�-` p/���0����>W���ι��r�G���um�(ص]����S�^�k��T�p�΍[    �����Ǧ�v���~�e�����0��E�:��߯+:1,2:      �>��z��������e�;�u��JN�����mnm�L��c,    ���6�9> PO`�e�:/LNK杧���9�d�����\2���~E�jՄ:q�6��&ĕ��P(S���-C���9kby����
pm'��[tm����v��{��=lgI��4q�*��]sN�y�um����]��C���y   @f�����^�k��/ee�s�4P�k���e\�yF�!;��!�N�N��      ������g��紂v�LSt�j�xeU)7�F8�\�s]w��ԓ����=�1    ���_� PO0������e��������]�Hx�=5j��P>r9aw����/�7��h�Mi(n�E�������0��KKvm����vmO��tm�}�:��=�k�\��j    Dvv����}�3��l�p�jӵ]Ӭ��}Eq���[�k����n5�,�*ωA�$��|��C��       4���F�.!�_�|��w�� U#Sh�|9C{\A T[���&    ��\�@�;?ۡ��Q��5����Y�A��H?��c�*�3F�������o���r����3(Q���R��5��bw�B��8 ����]�CL]�}Eٲ��$ճ����.ӵ]��Z    �^�O�	��Y76W���z�v�����
AH;��Ǚ�s�*9)��*N������Љ�!�*      ցaV�M�ļab���d7��	�,Fа"�3����3C TW��)u��3   �;��!찵��=���F�{�a�#w�q�V�{~4�F�LڝvꪈD����SyTx`j�����%P>���$�.ϵ=��%n���D*q��k�ԗ-����)�^q����!p   ���G�q���y����z�����k��ڮ�:�����N��P_r܃�za|�k�<�-vI���       � 3��[�D��.q�{���I��-wu0q;�(�1@     �F`|k6_�Rް�-e�_ۆ<�V���/��s��|!W�r<�& �{:�*����J,����Q�*��H\(A0��0�.�j�k����ȵ=^���c   �i�ظ�\��x��u���k��
w+���o5h�����Wn����S?*W�������܉aM      4�`���	��屾8�O�V�#|͜dM�ۋ�-���7 p���     4Ƒ��v`:O�d�N�;�d��wf��^�Njr�g�.���B��&���f	7��	q�3)\�(S⪘U�����!�ˮ�ĉ����\�#B�ԎPV�k�ܽ���r]���a�"]��Sl�[�0l�A    �i����"\�M��并��˴�uvm��k4���l��o5��@ռHw�'�+r3Z��Pџh       �`0���X�+�3٢{�A��oo���E��L��g2�1^�?/   �� �^o��nf����C�q�"g��B�Pz.nO�*3<�E1p��=�N����Ѝ!���Rߐ2�_���,k����m�s9^�
J�ȵ=ֶ�����]ۓm9pm���}U�v����3��͛p5   8d'���V74�6i�,�v�x4(�f-HNT��W�$�
2�+R��=4%R     �p5Y��Iqf���u�_�,n�jn0�]cY�5w   @�Ÿ��[;���X�ӭ���A�\_�����34�<b�Ӧ� �{ڭ�i���v⢛;&]���Q��]q�u�w�T���|?(ӵ]�N+��gԉ������=�'h��ӵ=,c�?�t���  �l��x�(µ]�@��4�vCq{IךO�nVw�v�����q᜷N��8F �����zb[r��m��4      ����t���ũ��w$lOI\7E\���yC;\�  �3�ш��~`�   ������@}����{5�j���>��BS��V�9���\ix���I�, �Lp����`X�f�����<��tmg(��M]�5�\�e}��	������U��Y�{�9ђ��a���~B�߻���/�K    �N��Ksm_Aܾ�k{�y���QWI�uu"�������gaA�U:Rcܯ�@��~��'      @���:4�ƻ0��ƄI~V�Z�<R��6�Z��`���C�Uj���}�����k    ��۷����@}]b�g�uA�.�)O�Mf�fX\/	�U9C.���w�)@��ߋ_.�M-�S\�n#�5!4ugpd��r�B��0�h:�R�n]a���9��u�B�k��8U�n�ھ8s�����g;��ג��.����8{<��hk�E   ��������i���sˮ��Z��s;�//n_յ������6��|�,�wU�*��'P��A*V3      �j�j�h:��%T#�D�����)V2��k|�����w+� ՙãCzt�.�   ���wn�/���@}�0����Ύ�����v̷�Kܕs{NG̻���1��a=��Vw��o��r�9*#�&����z���cQ��H�n���-v����,ѵ}�w��]�))_ڵ]rcOз�ڮ>��\ۅ㮋�|�   !7�nқ���B\�U�õݬ#�-�������ŀ@�T5Pe�2U±r���q�U      �-{q�u���0�����'����3dl��
W���r|rB����	    s�wvhpqA���9���@�4i��oڬ[�.�����4"�pݮp�s\��vs��͹�����V�-�M���X䮉L���C�������7Vwm�K�����v]��~Q ^�k���#�jv���L��G,�;�a   ��v�[8Z�v��sm_�����D�1��A��^����!P     @=�Z�x�N�|A7֟��#�	�'U"w]�`�4a�s�ilC�n��xL���I5e6�Q+��    ˏl�:���l��g��k�"ͷ��w?�a�-��-�'c~�9��\i����U���`��������Uڭ�d��`ss����\ t�vQ5N��m_����c�d�vm��z:Az�k�t���I~-�qm�w�   "�H�,��<a0cq{��<�V��4�����&�׉�//.	ء��*mP*�,�D�*u�
�*      ֈp���?�"Uݶ�QZ�����3�r�MI'���ሶw0�-M��      ��C��MY�,�[���LO9V#��UZ�לE����`<kQ�spo.U�j.ZO&��U��ʘ\�UYg����7o��0�2�n�L�vr����EQ�����}M\ۅ��?��n�   4���F�!���k��n�v]��6��_bIk42P�,�>����f�"wYC�	T     �.L�v<~'q�*I'��|nn �S�+A��U<�c,{0!��N3��    h8X�UkF�!;d�������yp<���#H���yY�<���7��=��6��U喃~�+�g�B7fC�}�6�Z���o�����u����}���'n��C�޵]|�tm��WWWt~z�i�'RI��\�Gz$��������Xj�\�������$k��/��d�J�~B}��P������)������jъ�kg�<�q��_^^�;`K��k��9W�O&g}3\�������嵳��3�a��5p���~4����s���ί�#��Za8��6��m'�6���Lo��?8;7vw��_D��˜���Ճ��̺M�<�y�d����ɉ���s�4�<�7n�>�� P�+�T�s������b�8f�;      �c�/v~&1�����7z^h%eq�^�����v��Ԙ�X    �0�LW��h�q�-�0_K���8�ǟ1��v�����%��3���=��G[�`=��O:�II��F\��0��L�/���C�j���_����*�^�\�^&4qտ����1���h�P<(Ҹ�����΄O�oފ7/'�W6�����UH)<9>&6���U��PInvN���oG.;=9���_��ӞuX�P�s'��B�������@�w*,.�����Q`��3�/�����J�����&^����=τήv�py��]���N'�q���[�}��oo����:8:�%�6Ջ_\��{�<|E�vS�{����mj�Z�P(e�zv�{-s�|u��	�ٜ������\��]�-�(�nݺ������t��.o��
�K�7k���     �c�Ue����Ry(1�,˺�ӎ���Juqg;�r���Z</_��j��{W�����7��㓹iE��\pq>�~��9������yS+�p.����>���\���f�k�r��_{����A`�����}�̙�!���Y�.M ]�w,o���������[&���O���_��]��{���kt9��S�c���C�c|vϹ�[�Q�yݹs����*�x��������y�0��MG��ae��Ϩ	@����أ��c���7�ue90�n�Ď����	1����ࠔ����	�\�g���U��O���{�&]�tm�cA�O?��X �s>7rm��3��Vp�Oo^��W�?|R�k��v�Ne�����(�De����O��a;Ͻ[w��l�p��=r�l6�P�M�l�������%��g�����+\�w�lQ�����{.py��g�Cl������l]^;���W�����MP]��g�$���G�Gt:���[7�-���svzJ}�qf]��\'"7;/V���?���Q]�����O��{���R��kN�v�{��)���d��rn�FY�
�h���gM�#:%UIq������0�G�@�/-x      8g<��E_�E��X���(U&�u(�ں�6ff�Pw+K�biL|�0���,D�vߟэ�{V�f���'g���a׽��C�H���֯����g?��~��/��]�.}e�⸮�f0����Y\jww�I߮_{����<�[�����w�q�?��{ޕ9����]3��7���u�i���}��:|W�w��ɩ�1��8#��7��햛�����K�c|��c����Ee�yX��h���D�8@Z��i�C���)�@��8��*e��H�jP)p��P��J%��UpP(��P4���_(�r�i�	ѶFHN�]�ħ	ă�^��=����[ �Nr9a����m露���{�>�ՑNU��|���5������Lq��^����  �n  ��IDAT �mn޼E��pX7��\�j�dX��t�G����<��4&�W;������	�A��`��V�U�/��x=�����_h@�� ���     `]�<�h�������:f;?'g���K�ܽ5�-�y($2�T0������U��3���b�n�k�?�^�G�����;]��>^����G�����v߻�����g�T쳯�������"3csտ�����L����5ؕ����.���{�>Y���>��^�S�wq��v6�`�g�t��X}�c��]�����|���>���<�p��}�a�0-�m:�Ͱ�T��D�0�1��.&5^�.�{�G3�;��q$�WM�6B=u�*!tc�(���^7�2�۷o(�p��u���(�k�P�8a{�@<�k{�?��{��G|���BJ^sY����(�8r�   �D�-n��KD^��� �vMFuWum��u'�??s��aӸ{�n��+��� U2P%
�S�}��Ѥ@      ��ńh;�r�TC�y��� n1��G�r��:��l��3��K�bpA��0��v2    ǃ��v� �s��Ma��2̧�b����
G�P�.�+���1�`ܜ�.�\rp<��A�9^Ȯup���bPkފ6q���=/�!�ځa���dsy��>�L������Z ��W�k��������\ї��]U��r�*   �-����d}�.\%�_M��Sߖ�ڞ�g*n��K��v`�4~���n��'�L��a�j�w�^�xI����@      ��E����M�d�g�^\!s��� �AV�w~f�X�|��r�    ���M�\`\k��H�J��Bm��X~.�#�����1�,�o
��`<����7C�=@|c�7b�����*�;Q�T<{{{�0\��M��.˵}�c��5��'�6qmW
�C!yѮ����Bv�q)�v�8Sa��n�Iާ��A��Ǐ�/�    ��0���l�x�v�)��ȍ�jO�������*ܺu��A"��^��R�┸������`�|�A      T���O���z�O䅯IS,mB\)lg��Bg��"��� ���3#e�   ��t�]��	�6�]	��2�4�"��P��I�C��}~���G��4���z��ጚ�9���4�L�`C�;�}.0��v@ws�V� p����|!p/ɵ������\�E�wm'ѵ���s��g�۽��?E�^�k;W���>��C   �
[�up|�|�a��Y�0��v��e����^�	�S��H�����a0W峎�����(;H�����0��ے��"~�?�      �Z�\^����1}�N讛7H	l�����v���e2��x<�_���;x�pxxH   @y��!�y�O��/.i6k��%��\-��u:�0q��D}Ew�;��	�$�������/��a;D�*������U"v��� �*��A�n������>.ϵ=C ԥ�]��sҜCQ����R��B�
�zX�Ե�/�N����E   @Sy��1�x�J,,A�n*l��5�W׵�Z�{l3h��`}E���9>+� �x\����]�ڼ(��n�`dW4      ��l4��v[X��'�u;?�[��u�V��s��7o�$`�������]W^�yM�<�/���   �&���#��_�;���]���N���<o�;^��*����)9v�K����e;׏O�1@���V�+��P���C�0��Jv���ba��+r��U<����K��������$\ۥ�b]۽ص]#W�{q���N����.p]���i  @s��ؠI��]��=�r��4�v���k�����	ء��4�@�i�J�DQ�8X���ɟE��      �I�z�.��&�I�[���5g��Ur����bp�{�9=;�O=%   ���7�4	�c�c��aY�Ue!��)=g��J���ۻEe��\����S���='�V/Le���8����3X�%+ڋ�W��[����$\�Sw��tAz$���/���mõ]�w��n��v   �(Z������j��F؝K�nV����U��������*����-��MԋHĸ@|�$P��:q�P�S�׬@      �D��[i��x~>gu��ynܸA��՟r�   �3��-�vp9Os�w4���*�h�;QjA6�nw��7��='�3�iHT�spO&��*�����"\<�c�N�����\�v�޲��~���W�߃E�����L]��g/��R��M]�úY"���(p�   ��>dcJJ�W���ʊzza�Q�"��D�Zq��9��+��>���w���|�Yg�>��p/����2~�O\�ɏn�Tq������      ��x����} &�s��崉d7v~����G����)��T#�   �߃�g��5���\���;&�s_Q+�.�R��a�0���R���='�Y�Z�ʈ�{��7n|��a���ʋ� ���N�⾿�O�\޽d��P쮪C���ĵ�Vvm7�Ǯ�gu��M��SM��tm�pՕ$Z_A����"��5�N�3�H   @�w���
e����z"[[�v���	ֳ:��\�u��߿OU�Ѷ�^4V��sٹ����}�֬լ@      �=^�r�X�<o8���pʡ1�r�34���"��t�o՟�hD�.b   �s�>Ů������6`�R]̯th��F"��D���q�K���d���g굩I@����E�aZ�Jn5 mC.܌�Q���~��/�*3�S���9m�A������&�1u�=#�����a��
�v��T�k�ԡҵ�TBrJ�G�'�������+��E�����l8���V��   4��}���j�m��t�
�vsq;��o�������(�~�Ow��u}ne
�{H����~tK��'�O�      �Ʉ�9�IIg"J���ɼ��9.����Y#l7ŵ;{0�{�ӡ1��AP����+�s���5   `�O>�����@��a�������V�l~�v|�pY����DjG��:_�I�1u�c� �99�"�$�@�p�rN!��[�����E�!uP�0w@`���3���m��8�v?�k{��<�_ڵ=!ʷ�ڞ�����ƹ��N��;  �Ʊ��M�W�\c\c�v�~5�:\��]+;�3$^�������0��ڭa��>*�ىRp�
R�Q�JC�Z���,t3#      @�Qgn-l%a</���$�ک-lU����)�e��s��ǳ��|��@�@T����^`�   4��7o��/��@}as����@�<~��z����\�U�st�X\Ԯ�K�ܵ���ߗ3f�5�� �{NNFD��@U�C��=,�׉�V'ǣ'Q)V/�o]T<�����(^UU�k�ؖ"��pm������T�v�8_�Vi��}��ڞ��V+p��F   4�v��kA��\]YQO�7�[	y������h6� ��6�U&�������mpA*��e^O!nWa.��z�       1���1�"�<�3e�ga~`��sx���"��(2��j��y)��3�L���6�6	�f�תЇ   `l�Z{&W�J���f���:oXt�Qg�g�3�����:=q2w�ZH?C�R8�����U�vn�|Ω��rM�*jK+lgTk�Y���m��prtLk��N��<�o���a`9���S���O֑]��kΉ�wm��m8����_��   �&���K�+��]Ʈ���fus֋���ԝ�ھ��}y���芀�Y��^[��G�dT�U\@��(�b��{>���      �����^�+����@7wH5��Y�Y睟a�Um�g�ל����-�q  �����G�1�z3�B��l���T���G}nҜU���9���ỳ�p���v��f-ހ�='��)�6Z�d4C�&:��n\��:煺�Bn߾M��G��U�k���^�k��ܗvm+Ku����\۹��hH>}
�;  ���駟ҫ�oR����\��޵]]���C�Z/�	�l\����6�;��7���0���G��     �t�x�N8�'�b�路�ȹC��Q��2�Z���ݻw	�apvNw�������>~���[   ��G�>�_�ｺ3�B����Eb�P7�����Xa���珇��|ߣn��L>+��~x��oF_���|�g.�ͷ��:�BnݺE���2]��B���@��Ĺ��˩A��B���666   h
��ߣ�����Wwm_M��^D��8�<�}�6!p�GY;lUm��u�J�0F�J.z˓1Y��~�.���       �F0^����$���8����a����'!n/~NT��"v~�����zsxtD���w   ������7���@�����h|�0(ʘǫ4�a�P#�Wc�e��7��}	���jx�8��*.�E��ŉoy����VyE�:��
�f+}����}��k��,Ӻ�+�J���N��|�]ۣs[\e���v�   ��n+˝���[��������.�������m����$W�+�8'�H��	P-:�T쇝��%��      T���)y=/�x'���b�M.T�iq�]���;7�z<v~����ug6�R��%   �)�q(�2�g|��-��7�I�7u��:-q��_H��uixJ��%hw��_^$VG���LZu�'��P:2'r�Q���������|J���4p����#q��k{RE�8.��µ])�V�#��'˔�v�/G��.)�m���\/�ѣG��w�   Pg�R7�L��1�kf��\��ԭ�k;������1�#���-�:�G�91h�T�"���M�C�     @Ua;?��}����j��=�.�͘K�c�~�;?��v��|�;��4L9�TZ%�   �
��	��&0b�g[d-@�s�0�|r����c��9.�����K0i��N�k^��)��!�O��M�
Ri��<iO�k��n{{�<x@/^� P>G�����]��d�U�v��yF�:���ѧ���   j�G}Do��G��ڮy
�/^�^+[�Űv`� ���u
F��p^.�wb�[Q�����\ݻ�M      T���&/.�c�Drz��b� �eeR1��]G�s�,g���������@}9<>�   Pg>|H���	ԛ�xwK�y�a�n���9��4��	ۉ���ߠ���\]�l�H�����Mɉ��χ����C������z��	�8<8��ˇ/\�\����k{X������텺�S���<
���v��N��{'   �χO?����7�ߥ����k�YG���u��tz|L�,�i�W�`T����]��W���NiB�c�q�yN      �^g�z ?H��DD��ryC?�F���w*��]~*m�S���Wm�޽{���Iʅ��g紻w�@}�Ջ��O>��  @�y��3�����@�9=9!`����ޞQݦ�u��E����$f'}!�ݼ�!�K0��i#�"��=d�7e��޼�*���љ��!@������w�R���?]��d[��v�k{���]�)�Ni�틺�\�墍�M8�   �=�~?XإB���L@���q�rD人Uܓ��������nG��9��hn��()~j<@���D���G      �j3]���/VM3Ǌۜȝ���d,�5H�/3%Z��b�ߧ�O��_|A�|N�O p�9���vo�   PwX�pt5"Po���y�X�K����v"}<@#j�bW�B�ǣ�W�ىH�
�����Nت:P%���.�g�&\� �n�a��b;��]�=y/�&����������kT	�UZ��:��A �׿�5   u����ԟ%���j����4��ԣկU>W8�ۃ�U$U۲0�-�������PȞ���~q��s9c��      �ː�ۥ1}�7#9�'M�PN|��yGy������]G�r��w;0��#����#   U��GgT�xT���SvX&o���[Ǽa\7+׭��B�.�-
��5-o������=R'��d5qu�d9���!l7�� �*mC�n��7o]�%7�EY �N���E�*�yY��:Y��j�������+(�n���}��� p  P[~��ҷ�^	ej]�f���`�y>a�j��r������><��ɶx�葲|��Q�m'�!�sX������E����lܼ@      ����M�)�z"��?,�&�bY>�m��e���s����?~L�p�lo�޽{���O   @a$�{��@������W�yC�����=��b��Q��K*?5/o���=��o�R���"ǅ0�-�[��T:�*�Vi�M�����hl��л�K����.	�%q{��z���b��
�e?{�w��   ��r��=��̝���j���P�^D�rD�UܯVW�Z�ˎ��ء����tI~�yT�ށ-�&�3F��Ǫ.a��j      T���G[|Z��V����C!�-΋usa��{��v�1�c,{��!�?_��+����=�  Ԗg�|L�?��@�������~)�V>o���6��#&M�@��~X�ܽ�@����F?3@�'�śS�s�4t�*��*�ȕ�"we���h��ӧ�j�h6k�
WЃ���sm'� ]�72���M��k;���d�2]ۅ��ybM�k{r��ڵ]�<���-��ڢ��   �F�3��uպ��f�u�k�a�e������ת�{�`VW�Z/*��c�����6���Zx��ɽ����X�\]���㓿��u��uq��9�      �ڰ���f�b��o�~� �+TDnqr���y�����J�w��%`���� ?�򴠾�[h~   ԑV��Y�N&t1��P�\�|.K�ބ��J�+�O�J�|{B\���=����o��r��3D�Vn��s���L�L
\��/C�W7o��o޼!P>�����#i{Gc���3�2�1A�^�k{�i/!�^Ƶ}�z��e����^�E������}���   P'����ٙ������8�X�.U<|@�l�ɶ���kB9m�/�$���?<��DN������.��.�      T�w�3j�l��}i~@~���8�ķ2������V��*��p~ZV��0!���ݸ�G��\M'������   �:��΃�%��sr|�9�%�|�ɓ'���a�����J�I�7�ڑ��t:t6j�Bܗ��'��<�bh�U���p�E�*����Si�*�Wm��nӇ~��%޼zE��{�;P�k���òk�\Y��S�k{��]����ڞ�X8��z ���C   ��g?�����X�����nMD��WQpO��f���@�n����Lw�5t	A*�Bt9������ƽ=�$����&��v      �Δ��76h2����� �7$
S��"D7៏r9E�:��[dw�6=	�������o���}����?�9   u������/	ԟ�Cv���-dg����c伡����c��!505���L��^Ȯ
4)n�P�>��!��<J�pZ�\�tW���ӧO����4m�7/_��(ҵݳ�ڮ8�[��]��'���.���܄�	  ����dI�I\��hµ]�Mq���oVq�*���裏���m+����{�q� %��k\?��      փv���3e"��NVS4_P9�e��ù��;(H䮣
�E�������+�s|xDO?~F���{G���o@�  �v0��_��?la&���L�n7z��a�w�$fW�de�۝>5ܗd�w��U���.q]~�Bw"i������Q������vx��5Mg3�[qኮ���`^hյ=������9�F��+�v��{=.//�����   �:�v���_�Za��`=�k�\\�����{}Fm�qm�K p�I�cQi.���=��H�ߩ��ǭ      քv�z�=�'._�����OL�E�T�iO�)PO�ȶY[l�g�� '����	   �l�8#���L`��Jސ���!p98�h;����ȍAvb��A+I�k�� �*�>z􈶷��(x�A۴Z�@|�~�����ǏL�[��[%$O�������뗯�����q᭑�^1��e������~f����Ǥ�ۗ<Y�껗����D&bt�/pš/_|G��W�n������ϩl�A���}���Z�N�Ex<��Ņ��ٵk�W,prr���F�9��嵻���l�.�j�&.�������Eq������eN�p��O��`{���_���kp�x>��<������w�����r�i�S�������ſ�<o��'r}c\W^^����ø0�)$*f�����9�˱=�u�:�</�஢Lׄ4�n�O�����n��M����: -�W��=7ߡ      ��L�^jr�T�)]�Ĺ��%�*2��T-����G�7������ݻ���;   � �^{��5����'�nt!M����@�0��R�0,���z7��`H�9�e�����/����▌D�eǶ��+��~��I����t�s�vEֵ߹���o�(���Έ�M�2&n��?����a�o_�~?y���v�����П�ş�'�<S7�����㿡?�˿�ˮ�{@����Qټy�nݺ]��7�гgϜ�̈́�Lpz��='�����>}J�`BWW����q����=��v��� 8�*���iypy�lA�۷o_�l��ׯ�Ν;��|����g����*E���A]&n�!?6�V��f��/~�o���=�v���� X�q��}�s��3�������5��ؾ*��(���Q�Z[�Ґh.�A<�W��x@�����l�      �>�~�<����'�ùH,lO1ÒY��9��P�W��?�E�1����U<��ڿ����~��89<��̍�����N�N��u#�8=:��_~�of2�����0*��W�������ߖ����9����ܸ̞4ܜ����]��v�9ˮ����I�gggA�M4g
��\�N�y��8_>����Ɖ��y��_.�wt=Ʋ7�G���H�?.���s���]}ޥQ��Rւc�S�S6~qc��ܗ��O����vn5��Ɛtb��ԫ?��w�殐&�b��Ѝ���7o�7�	�"�(�D�J�׉��zi"y�P���|,Y�D}EJv�8Sq��"xR��}�ci5q;�b��9�gp�w�E7o���   �:þC[���`]W/_�UE�y�_}^��ˮk*lW�8�{��=;����,�ܪ�Ӷ4��V��XM�Ȃ�<�����?      jN�Z�g8֏P$�żaXM�FXq�]���jn��Ç�P��ss%<�&�D���k��ݦ�O�c����o���޾|E�7�h˕Q˗_ӳ�����00�x�Dt��?��?��������l�r��3noo�I�M~����igg'0hr�ks&fN�j��/_&*�v{w�ڳ�X6faN�.x����?��?��_��pK���y���{���펽1֋_=ƴ����V�666��})�ua���;_g��V��yãQ3��/����;}����pÆh�]��@��-���>�&LT��W_(�W߽�(\������T�ĵ�O���*)�[�k�'��e���da��=x����o-��������ߧ��o��   �u�g����n�� xl*B_YOe��Wܛ�S��y�~�sUUֿT�g�c{l[�����,�dߑ!yK�v�"�%��]�/�$�g����98      �xޜ�0�'ʄ�v2o��[+���|ar|e����ǇG�	�A������[!   `
ә�_^hǇ�ڂ�?�����������z��W`cs����"w~F�ffdz»�0hR������=�-������Z$�Ƴ]�)ݑ=���]�3��&��K���(����28�r��'��Z�v�̣���H   �����'�������RW0�;�WUpoxR����vm�R��o���G}D���Fu����Ϲ�����#E񀤰E��a����f�      XG�;��g7��{�>o(��!)��3��<OS���U�-2�۷o�{��f&p��g��9��G�E���H   �:�����_��6w����r|tL�O�<1މ��y��Q&yì���=�P������Bo�f��vF� ����58>=*�7h�N�+&� v`� ����{�/7�4��)�hE':�I���TKݚ�3����={�������|؝�}f����}�Lw�{Q��#)�˰��@nP	��HD"��D����f!�EFJ ���c�f]&)�k;�qU�E�x���q�e�.��zX��\�3��������"���� �B���[U�cb��ax�"��	���>�U�~��{��$&������oDG�����`i�}F�\�9 �XEgklnEr�4cqB!�BH�YM	c�f$	��ȍ<�Vdm���e�gA	�n��-���R�|�+���E�hB!q���+��h��1�$�N��Q��P�mM^uC��uк�1Qy�v�XF������ ��,�;�~dn�X�H��AٳgHx�d�Epmr�g�G��X�c;�E�յ��~.J�ڮ�[��3����B)G�;����]�zQD�A����kwC��V<_��k���#���uX2Ѹ��_I+���9q���$Uډ���B!��򢮱���ܽ�kIqU�����X���)�b�{��A|��� �gyis�shmk���-ΧW󛝝!�R�l޼3ss ����4VWVA�a����yM��q[���u��a}�Nա�= s�48�S�*�+p'��Y\I+k����W{��-�;}�8u�L�\۫�O��yl�cP�\�e}����6hӵ���X?>f\"���m�A!��+��ǧ_}�k�!X�k{��Dܮ~�Աc#���d��e�1�T��!�$�u{�j=����RH�������B!��r#UӸv??�]����(n�#��8��P�>VQ�%r/������b�g
�+��~��'�՝; �Bʑ'O��R��p��0��uCE;���qܓܕc}eݰ�
�_�®��(�u��6{�*w���L��xg&J*F|�A�N���X]嬫0��ۭ��u]�AZ.煸������͸|��fl�]�n��һ�;��_۶m�r��B��$uU���݊��][:y�zq�XC��j��=��&c#� �JT��T�W��>�Ȏ��`O\YXYщՍQ[H�tW) �B!��X2괄�m�`/p�
��
�8����z+?�cmq��� �!V��{� ��gqqͭ� �Bʕچ:$	TUW�l|&�s
aP\(�Q7tO'׭fb��z/ݰV�0U���$*
��7���:�c{�vHUr7Y"G���м�ܒW�}b)4��ųg�@J���������T4�v�Ūr���p�XTZ�퐈��v[�W�����XY�[�������3����A!�����*z�}	�K""��)lW�W��u?�y�{�)l�+�SI8�	Ư��
�%FϿ�p#n�ds�H%&������';i^�1�m��5���B!���bj��ƺÚ֊�pL���J�#f�+�_��R\k���+?����8H�03?���LOO�B)'�n݊�	޷Tc���x���e"T/��!�1V��åVˬN,��:���/�P�������WQ���ȴ��擬N~E�P�z1��СC������o�oX�k�LHO�|�؎ߊ�sm�}8c��n�K$�ر�%B!�ƞ�/㇟��u���҉�K%�74�����U��}I��0?7b�������x�у�+��j ��{=^���HD9U)��e`��vB!�Bʍ�y�)]q����,l�'��H�s�)�¸
ԃ�Ӯ]��e��Sx
���ql5�P+���<Ĺ�'p��; �Bʉ�'����wA*�Օ�Nπ�Þ={�c06JMQZ7���t��Z�G�p=��� �U�n
���Ԃ��E��*8�t��Pb)
���0�����p$�1�ߏ��epm�]��pmw��+��um7?c��˞�k{���4Rx饗02BWTB!偘%^U-�7˵ݗ�<��� �T�ך��bGy�*�.i"�JT�,[��p_�j��[|b&� ����|B��w��T�v\$�B!�����$�HL��j��U���bY�V�b��`~�ul��0Ƣ�=�+��O`��m ���e4�4�B)7j�밚H�T½=
�c���M��o��ڻ�u��6W���̵���^E��)pHuCR���v�_��q��zJ�U����[�J8��������W�\��	��q�>Bwm��*׵��66>�3g���w�!�R�8q=�}���CB{P,D�q��ũb��)XW�l�ر�Q���*Q'��ݯ�r43W�Zلu�0E��r�\̤UcS+�����"�B!��YJc�f���ܽ�XN�sl�.r�c'�63X��ݤ�̯���o��$&��(p� �fg�y�fLNN�B)�����H����Hx���+�n��<U�P>�]�9�M--HNUnݐ����޽4�����u�1��:Kc�Ų�>S&N���t�رȒn�HwW��-v���s��[{4�J�ڮ)lõ=ݳC�n�K&ؼcgzyI!�!�B��������E-"�S�T��K���>�~���P2�W�����c�A�����%9n\]�rQ�]w>��K؎�y �7��#�66�B!�R��74aq~6��i�%7xM�d��'���C�r�-�j�J�ё�@*��~ƥ�g��g��B)^;�:>��5H� �IxD1��S�0���&�K��'�L��m��U�(p�\�u��K/aeMRy�ܰ84��.�jx35�Ll�ݻ[�l�r�!�������ع#�k{���q$�k/q��k�뜊����n�K�^����{�����Y����x��!��8#܃�bk�s��5��ب�ŏ5�o��`]q���+�LT����x�ȑ؈�u�wN����Ð��q'����
a��9�M�{���B!���$U״v_?��Ȫ]34��ng�Љ5�`X7�Y�p��&PzN����0Q+���467�|�BHY jյ5H&� ���?��i���JQ7����w��p���� �a���:Wzݐ���Wc�Y��tn�ۭ�n�� .#�/��lm������]��s���I���� ���v�ڙMf����Cr��ҵ�޴����vm��Q��k�����65=�#G�P�N!$��=����wD."W��Ϋt�� �T�����bĮ5��p�������8��r���m�hD9ݰ��'�K��<��7��*^�B!��#KhP��k���-��]�XV�AI	ͱ�Xw4W~nll���H�YZ\������A*�']�i!�ӧOA!�ę׏��_�>��&&��X$��� (i��E�ZU7��)�c�������k2��M�^`)���� ���;a�tb��JD)�W�$��=J�{��tu���鿳�vG]�m��q.q{	\��q��:E���������4!��8"~����HZD."����9��+���Ǫ�U[��8�Xk���0Hx���k�	�&��֞��4�ݞ��cv�DU6��pu]�(p'�B!�,�X�A�b�&]�,U�Њm�(Zk�V����k_KK:��������Do��y��Bbώ]���Jbt�u�0����겏�#Fף����p�=��=�w�a��T���Q��ܺ!��[I�ik#�	������"����3P�h7���<��]�U�\n0\:�>KO�p9�4]ۥbw��Z*l(��\�Q�+�k����s�+�k�3nxl.^��B!$�����\�cu�)L�|�v�� �T��A�P`�?���A����Rn�n��L��}�����yU�������&+7IE!�BH��b6�v�b��G��8�ǲ���!�e�B�z��b~�ū��J�{������� ����Rz2���<!��8"���fi�Xi���IxR7�"�5E[�б���FX.���~�k��B�t��E�����I�D�ډAqa˶�8�C���d����^y����NLL`۶m���]��b���n��\��P]��m��K$ص{Od�[!��|�;����y���pa����b��Vչ��F��w�1%��T�#� ᡚX\N�
��	���cҊʅ!7�ϵio��������S3�B!�R�N�prs��@��zM�������1��@��^XN�W^�X7
�*����gN��/��:!��xr��Y|��]��b|t$<��Y2�6��ۯﺡu��mR�ӭY2C,��]�7^o��o��te�)p/ɚ��jJZ��ve�� ��92gf���� �09K<\^t��������{��[���cG���cB!q���ˉU��܏�=��\%�5�)�rL��=�`
4������b�E������'����7�VM�n�q}�	�I�M\�B!��r&�v_��ڊ����_�,׸���6/�^��V�����	�ŵ�{~n-k�:�����m�BH���55XY]�������*c,ʡ����U��UՍ��j	�%�㦶v����(p/3�z�).8�ŘW����賛K�j�������}���8v����;�p��������æl*�k�zlY��{���mF�8�b�o����|<5=��^{�wB!�����x������\O�n(��/�XC?V%"�=���O�f�y^#C� �!&>�r��$�˶�b��5�Sg�w�,5��k!�B!����o�1?o���4��Z��qG��ݺ�ڇ��Xn�W����W_EMM���^�=LF�F�r���J�yowZ����B!$N[�|�����B�"��8.&V��V7�����{��S����z��KoW:��х*�r\h�|�s��q�ex3���D��
�NzQ�.O��Y�f/ĵ] �gv��<붧�]�]}����˄�A\������
���.�3��󿅁����@!$n467cee%�8L���]u^��������X�K-Lp?��b�c}}}�q98+�"�ב���8�O:����I*�C&a��|R��dB!�R�,��6�Uo�`�p��:k�Yr��b�u8c�(�[�lI��?NaSXAсï�T�{��浛�B�{^~|�	He!&\���X��}6�
�.e�u�mF�qzn��{�d��Y����V�
����)�l�̢(`�A��]'aeub��G��E!�+1+�����"FF��c�N=�v��Ј(����ID�"xw�����*�u���ΰP\۽D��F�}å˗�ч�B�G����P�q�"r�
[�S8�����P� M�z@��y���bl���_!p/&qOtY�Rִ�r�r/�K�]KY��B!��7�+5hi���A�Vl�Κ��swPW�"\�)p���A��c%�@SSS�nL!��a�8�0RY�����Hx#ⰈCMѡgϴ��9 ��N�2c,�6�$�����.�а��^��qq�n�<�r�t�0�C
��'W�|��-� ����Jܵ]��jC"�N����8���cU�v�!�k��+�gc)]ۭm��v����k7����?��BH�>zw�>��R��"��\�b�4�)�+}�
��/5��^$�x/.G�>k2�㞠G�sr&�I�J5�<7n�'P�&�L��E��3Mq;!�B!�Nߌ�W٪My�	ʱ�z2�5ga��k5ȉr�f�P.�򗿀����"f�g���R9|��G�>s_ݹB!$�=w�>��������MJO��q�)�8��_��~��Ms�B�T��ɣ��"��܊��i�������� �*���%�u�t��y�ɑ#G�i�&LMM����'Op����c?��6��C�]��*{c&�p�vg�/�v��8#Pl�:��6C����ə�A�Yܻ{�BH��ر�33J��4۟0\����4����y�Ā��u�8_��4�7 ��88$���0W"t��6��^cxuK����؈�N� �B!���N��M59a��K�f��*�U��F?y��q2�
��Ƶ��Q���_X@k{��!�Ă���6�ayy���{{��q�X1+���a��4ho+�k��f^`�����4Ƣ��X$j��2����)(�e�W�ʌg�K�I���Z�8q��9H8�<�J;z�/�R���+sm�v{<�P=W��r4�]�ak˵�u����#�6��:|��B"���s���GW{iD��*v��^� �c���u��c}��}	�s����Ƕm۰�~đb%�̱��M�y$�;2X������B!�BH��\��onk��kb���"�е��1ctd��k�AꇢfXWWG'���W��T?���O����B���gN��H�120---���͑��P����U��f(5�b�0�Eb>U���pc(l�_��Ȋ�s1*!kT"t?�
������H"�@_��]ǵ=���܏`]*:7�򸶫����~����킢����nH�W���'O�>!����XY���K�NDn脭7_�^
�ZDP����M�󘙚	�ӧO��OL��P|,��R��>�&��ݜ"�d]3!�B!����{Ø�Nn-�f�[^3��#菵�ʤ�h�'rG�U�~	�ѡ���V�y��adl�^}�wB!��y�V|����Bh��G�@���ɓ����>�Sݰ�5E��=7��z���]O�r� Ǻa
܋��Bv���B������a&�T1��C�b�N��K!ɫC�������Y�{9���D��vm�ƹ��7�T���ؠ��p�NNO���S�B��KW.�g����������avX�u?�y��*��yP_"x�dM�� �Zf��LV��s}�=L뻵R:I*�x>Y�vd.�M!�B�F`��q�^?��઻���laݲ�c�O��O\�pq��=<Lq��/�T��}8x� ���@!�D��c<���P%bN�$�!��@duC�x;����˚+X��bR�u
܋ĳ�$v6���0���$�&IV�b2��>�quW�O|��%iV)<}�o����]�a�Q�#X����8���*�A{T��n�W�����Z �{Umv�܉��!B!a"��������j��X=�u���"�b��W���C������=T���Xf�R�%����O��'�e�J{E�u��HT��|&�!�B�L�Ԡ-eX�d���@5��.n�aH�*��A��C�-	���!
�+�g]�x��-
�	!�D�������>�<��Y
�ÇK�����[�P�����uj�NSm��.���X7���H̯h�ֆ��{� ݋TZ,���N���!d-w�'Bl+f�?�$�����,��۳me���n�q.Ѻy���smwoxt/_��?A!����K���I�D�Je��)�=X��k����Ep�X_"x���k�߇��R[[��^{-6���gMPIw�k��=�3Q�˅��3H;���B!�����I'�r+?�c��-JͲ�cG�K'7��B�	'ϸ�47*��8~�H�11=�m۶all�BH��ڵÃ ���"�W�P7�����a�I61ݭ�Ͷ���m+�Y��'(nP�^Dj�Z��<f��dK
�Kz�`��q;A�~VK��+�ŝ�p�|։�����.�������j"l�vm�r}��pmw�� �D������bnn�BH�ߠ����������@�v���� ��<�`]3Nլ+lwƎ�`yi	$<��ݖ-[���\*�>�X��ĐW@R�ř3him��4U�B!�lg���RCV�n-T�����c˄���y&�
�!M~�С��vtt$&�'����ƦF��⧟�֥���Ï@!��ɉS�����T�󘙚	��{���_�FB���[k� $cv��]U3T����1ɺa
܋�bU�t6���ݙ����Y����P
]��P�}���3Hx<��g�;.�wV�g�vC!x)�k;����Nq{�]��{7<6�kׯ��w�!��N�Bw��5��\���4E-X�ӿ�|=���ՍU�u����~�p9y�$*���1v�gfC5d�:r5�m �B!�l,[ڱ8;��甬 n/������fX���=&z�XUU�W?���8q}D�mX��~� �RY�ﶕd---���!�����P�4�>/X7Q���Ƣ6�*�>7��a���;#�5򜑵s\�e��J����Y74����/Vc�5Ie��N)��.�[���YŴ�>�ŕ���_G[��u]]����}�D[}�}�}���OP]S�~\��������O?����&V����;3�����ӣy<�gD"(W���U�{�������̿r|��Z�~��)�����<Z�[��ۛ�.�p}[T�������#�{uu+++XXX���ړɤ���1�����_Zw����f���Td�]�u/�w�{#�(���W��.�HDҿ�[\�Q}�}݉����aK�Z���]������Y�}��>�G�����ޡ;�:���8�������Z(�?��%�����<�W5�w��7�"Y>���%Q�����:v옴����V�}�q�z�{R�鞨?�ݖ�&�ֶ4��PB!�BH�HԴ��&�c �)��v���	��M�����n3���Cq�c�X����>�_jjj"�_���k��� }����=�
z�xݢ�����(X]Y���rd5�d"�k_^{������ĩ������~��[-E�r���Gտ��ﰨ���������BT��(�;�]������wͺ�$l����5�{��>�gΝ�W�~�D26�}�om���D��X+���k��}+��t�[���7�O��ߋB�a<,����k��}�nN��g<��v�4�r�E�ruH��}�ʘΉ������Y�nVq��b7����*k��mSUU�$���]�+�T~�r6�����ňn$���w�ٍ�G��$��P�����_����q��vm7����϶�rmw���$���I}�ɧ�q�Vd��}�	n���3%�g���~�ڽr��o���!l޼�!�<p�@$}����,v��I�bB¾}�Q��B`.~CĵQ����� 777k	SKA��]$����#[�kpp0�sT�����mC[+6@��\�Ų�{��)�Ւ��}� ���N�W���"�z�O��#���k�`jb2�����v�yyT�^������Ͽ�.Q;E��ԩ��y�pp/��Ai	z��P:��Dn�U����R��|�{J21~lI�gVA!�B�8L�֡�HI��~W�2�2I��	��5i/��Za�r����bbLU>M�M#�(��E^H/r���\ZX����`a~>�y�J�%���'VX���os[�&�~bGQÉ
!8�����{V,�~��_�3Ң����Q�k7E�Q�����wET�u�yT�]�-��Q���|�b^��~���c##Z�������B��'#��[Z��q�!�wĵ_,R�f�g��[���7��Q]w^��[�P�ɟ���&����.���6�,�;�n(����L.�м�	Ʉ{v���E�R^��͒���L��M�t���=}�tAn�p�>~��+D׆D8-�{�U�3q��*��<��nt!�W��V�~w$q�;���+����m�v�s��)l��󾯬���={�B����B*��������0�X=�u���"�����s��С@7��?]a�:6�6�$\�d�W^)|I����y��ڱ�S&�MHώٝ��+���f���d4MB!�BH����]�ِ��c���:�q���Xq���w��ق�4B��1��[1@~(�k����K�v�\����=�qʹm�@sDF-bUĨ^��Zߵu���O�V���ĝ/��z�<��Y�5S���znڴ)��+���w���i��(��s&��!�0�پ}{d"o�;�k&4bb�x�Q�k7�/�u�7������$����}��h�o��cwa�ܔ{����E|߶����Ezr�n�Q�ۛ��,F�ޯ���"��
Y�pV/�>�k��f��ayk�5��֟�5�	QA�{��oj��̤ˑ���>�%������rbv�s6�-�*iu��)
�C�������븶kŭ�۵]W܎*�Ъ
���^q�P\W؞nUL p�i�3{���;�F&�p��M|��� �BJ�,��y��v�����S���k���\�׵�J_��p9��kr��r�gx\��M��Rmv1Jʐ��S)�s��[�'��"�B!d��;��k�k������]�.���1F2��������ҫ?��� �1��_����7B����Bc,B!%���		#K�0	����p9w�\�Ϥ��<k�^�r�l9֚!�f������������c�P�^d����.�q��
��w�Ju�g?$�f�ʗ���*��
s��������Ȉm�����.(o�v�ݩ'�'Z׉�OѦ-n��2�v�+E�.�7	�=;v2YE!�d�;x ��p���GX�+l�4_�4��q���v?�������9���'I����WɈ��zq�J�a[�{�aMd�T��Ĺ����B!���Gr�~����s9C,Պ�V�6e��^X7q	��Ͱc�{q���N�{���σT&_}�-�_��/���BH)�|�
��p�r��=l��pe`�f���(Y�ݡ��S�S^� ��X�H
܋��J-�,�jg�ZZ�NɒUގq&2�9��t>=A���A��>}:=[O,�C��ɣ�i�����ϵ=�l�s�R��pm�ŕ�k�3ntr��x��!��br��I���ݻ�����}��Op���U�k`���1}	�5�T}A�~���L$<��މ'B�/�}����=�?^�u`0ۗ��Y�B!��-H�����]1nH�
้��L�l�w3���se�6q��s�pp�1V����afz�� ��pӭk�Gcc#���@!����,'Wi�X�L��c����#�U2�P�+�>Ǆr��Z��~��c�o���d��DMH
܋���NVIfWH�U�6庸��*+�6I�*��7��y(N�J��Ϝ9�/��$<���#nܾ�%:7��m"s3n������ڵ��~��u���θ��U��s���9��BH��Q{����g\���w�avp���ؠ"�u�8U�Z�����{��A�e���8v��\
�O༗7]�w�:I*��==q�>�����ZOT���@�B!����L��)y�0�����2�aH�t�C�^�z�}�fXSS�D�c�0|ч���A*�o�����.�O?!�RL.]��/�}R���L.b�0���*�ڠΊ��ڡ�nh(�#����87����.�N�ցu�����.lopϮ��#Y%��B]ˇ�p:0YA�I�M�B,�A�{���crr[�l�4d�rq���B]ۑ��µ]7�0T�b�����[��_�B!��>s�=]�u��X��ZҤ/�Kخ�U��
�u��Kp�>p��/�K�bYk*/^Dmm.E��RP��v�N�q����*^�&�$B1Q�B!��1y1W�����c���X�%z��q��l8��ȭ[��'q?|�$<�zzq������jkh�E!�����bae	+�� �K��p�����$�_�P�;|�y�v���=>�������v,�NggZ����\�:2�Uָx
�K�� 	��??��פ�s�k{�ܹf���l,�k���һ���S�i���z�`]ߵ���.�Ov�܅��6��΂B	���ڵg7����"B&���g����µ]}�c}	�5c5�Bܾ��De�qHJO4!sa�?&�wU�� �y����Q�N!�B�F�s"��Ȏ�u�|�g�c�<c�9��YV\j}A�99{�,�!39>���9�X�0�������|�">��B!��ҕ����; ����4f����ӧO�8q2�r���G��5C�����sʜ��m������Jd��I������ֵn2���ǒ�̝�D��!����KKK ����?���ktm��C66��w��K��nA�ܮ���������_�
B!$�ϟǳu�v;*�^A�P>_�W�X��\S��)"Wӗ�^3N՗</�z@�E�?~����>kj
J�v_����w��{s�`�B!���j�@s{V�uC���ڡ�.���Y����ns�8	�i��1������_�L�W���ʸ���́B	B{{;f��Ƌ�r���y�U�=}UU�����j���f(�*r�MH���朼�Y;\ۚ�:����@T
�����:tH
�Ra{�����]X�aKT�	��pI��9���'p��]��x�ۋ�il�ؔ~l
�]��R����������W�c7�k{����õ�~@2�D��m������4!��B����܁�.�v�[!��\�+U��Y�v�SRח`]3֧�^���_􁄋H���	���t�槠vbp?G1.�LTW
U��z�ru�}�	!�B!eGCR�sҺ�z�g��!nי��^ ȞBf��ĝ 5L��.�M��A£����
��{���K���A!�A��t�s�ʦ��H���ק�Sq�񕂜P�ږgܭ��j���1V����%��x�kSҋP~�z�܀��aG���Ǥ��,���r��=|���8}c�ϵ�&{+��u�ܮ����.:w����,�k;4��;��z��@!���k���E!�V��]M��K[5�J�\����c�����..\@]]]�q9'���!+j7���*���Dx"�ԮJT-���*!�B!��d��˙-��������1VX�Z�c�ر�'O@�cblK��hlj�LV	�$Wӆ
333 �B
a�֭����d�
gnv�SS �"�Ž�IX��(�κavlI��f��S�񾗸]l�+�k=r�
+����Zv� ��p]��V}q;g|T�wy���q�e���jߙ3gBs�'9��.]�\|�v��Mi%���%lW�mD�vY�vmw�'D=5u�8p� ���A!������M��<�:�h
ƃ�K#���+Ϡ y��Ԃ{�� ����>�Ν��3a��{�1�u,m}N^��c/[�-;���֘�!�B!���*u��X��.zOIk�^�XY�B��1�}w\j}A�9�)p�ߦ���z�r���{x��u|�� �B
���Kx�A*���^��9��vl���B�9��.� U�;_��Hyc)Vx{:Iͫ
�KDMSV�G�3.d"w�s{Jq�{$��[VPk(��a�$xQ�����mmm���,Hxt>}��5�ڶ�L�!�ѐ�����;�%n�ĕڵ��f������v��\�u����;cG'�p�����p�	!�_�z�6����"r��Z�d���ǪE䚂��"x_�{?�����h����Muuuz�W�u�Iw�ò�]��6s�nNBw����Đ�����nY?M��}�B!���N��*�o��Z�9;�P��������X�:FPs�BS�~��i����	�ߡ����i}�C�`?z�ihA!�G�����ԝ���n6bl%�U������k��K��9��ݜ�w�1��f(�mni�� �N(p/�h#7���\��}9��L�?G��)�r�~���>-����A�嗇?���˱wm]�q��������g��ݻ �Btعk��f����ڧ��������XC#������=b}	�5c�7SZOW����A,--��ˮ�ϠH{Q~I)�~2������`D�[*�R�k�T7v�B!���1�*4�n��씭^�9vȎ5�.�	�y�f��H�ެ����F���]�t	����7���������R�<�|�߾�z{z)P$���0�9x����G ����&�'@�E��~��ٲ���ϡǵ��}O6W������ؼ��%��\5�(�!�.;`���R��UI)�D���6��e�&�T��Ν��=�~�-.]��h���+��ݍ�8�g�v�k�@��θ��9=v��	+++ �B�q��E|q�kW���Ї0�8�u�8�X��{��vu���իWm��qHX����r�݉�֖w�+���8r3)Q�!�B!��rM��X`B��Tܞ�j����9\�ӕI�PF�k�^X���с�'O��o�	��������@*�����3g���߃B��¥���ӏ �EW7H����M�Y����vh�*�堮%Z5�*lU�P�/Cmg\�����D<M`oG���t^�v'����r�qHh�x1���O_����a�m��qrm�	��Bt��%�vq���|�����]�!�+��oxl�n����B!ċ��N��}�Z彟�`����u�0E�rm� ��^36��[c���zzA§���X�ڧ�^��&��x�D�غg�q� �B!�D��r6)��ұ�ȇ�P�\�Y>f�b�w2[��Xs��,��p���w���7:���^K��Nc,B!�hjjBcs3&&��M��'�{@�G��k�^X���v�p�to�ku��T�5k�K�ء��D����v,/�ۖ�9�e/h�,_��DUF�.v�~�A���^{�5�޽ �������mM7���{����3t�
tm��IK������ۛ�smwƮ��b�Νزe&&8� �"���/�ۋ����m���f�J�.��F��US��WDD�P���ɮ�Z�_�!��{؈�����c���8���xں��8���.�[��ּ@MM5:�WQ�	�B!��x�h,������%�mL�{�|�Y\�X���`���\#T�;}�4H����anv�mm �͝{����+��OA!�xq��5|~�k259���i��Qǳ���L��V�j���������N-�@��
�K��Ў�ܬbօ�蝛ɑ���)��־d�*�{��R�S]]�^.��#H�|��7����6�h�p���@۷k�K`noL��Qe_� ��|m�4N!�7�?����~b�q�øy�6����B!D���7���/鿕�����RN�
[I����
=�] �s��q�ر�3&�	+���'���8���U�b���}3��B!�R)L-&Ѽ��+�9�+����v����w�=��y�2�	.l/A�hlڴ	SSS �"\�_;u��Y\\�J2Ac,B!�l߾�s�\��}�>�v�±c�bQ�Y��RS,���*c,������S�ˠ�����ԣ�Zȶ�eEoC� ��eq%�r�&��qHh��@�{����ap`�v��
�%�k�F�[�^t��u7vC3�}<�bvmw�K' �vmw��NJ���j�iU:���NB!V���Q[_���y�}�R��`=�of��ͥrm�=Cf �����~��˴[٨	+�3'%sb�?�˽]�(�Kr��- �B!�T5M�XYQ.I.K����O�0�a��uuu�x�"�{�=�p�������������[x�wA!��8����C"���	�+W��W6���U�}&�ڡ�fX��۩�U��,�4p�+����)�uñ��b�A�����5�U�{��z�~�K����˨��E"� 	��~�	;w�;E�R�q��=�k{�/k\Vd�+X�'lw����\���a;�1��A��;&&'q��%tuue�S!�B�o\���?h���ڮ��{��]������j������B�.v�}^�+d_X���=�[-�U�Jm�I�#�k=��B!�R9���v��b]c
����cK�gѻ�R�>��3���Ħ-�A*��=�Gc,B!R�;�_:�M�Fʛ����̓�ϙ3g��q��AZ;t�3M^cn�~���i��z��;��D�Z�Թʠ����M'p��iA[v[gpd.�TZ�.�px�JTY�K��`1����;w��ѣ���A�廻w�߾��˵��h��rm�;.�k��|1��a�yč��.k�����7��'��B9z��H&��J��߬�߂�f����q��k;�b���ݝ�A§���ϟ/k�=8��ck��)�ߪD�s»�:�I�B!�T���ؗJ���e+>\�Y 3�rcdk&q�r�����_D��=��4O;���7ޤ1!�b��}����>!q�H�G8�_�t�,�����ܣ�@5Ô�_�8����p��9����ж�S�v�l����B�������ڵk�G���4�?��GC��.C%n�=���[�@�n	v�����
�!�X��%�)�o��Kس{�mۆ��!B�l���q��Q|�ݷ���������O�k���Bjo������0H�\�z�����~I喰�`q1���%�rb��t�dv�+csk+F�� �B!�TO�8���=!VR���+?��1N\m���n.�o��E��A�F�ݻ��� ����'Ξ.�$zR�|u�[\�v_|�9!������o@�@����y����*v�����❃E]�z���\+?Kk����\��P�U�9f�A�{��C�R�YQ{\��~w���]�*����%Ո>���G�	���j
�ڮ�]�.��G̸����ѵ�y���!��7��ÇA!�����m����\�R�]�߬�ڮ/�WtԵ�G�����g � �K2���P�c9�R��3�N��D��q�,Q�MR������M �B!�T��ܱ�3�Rw���l�m����i�%0�@:ò�8����7o�w��H�,.,bx`;��!3��X1رs'���A!��ٽg&g���� B�}XY^	�7n�ǽ����Cg���果�Q3����Ա�(��*(p/1�S�x%�t�u��-c������nXE��$��+��rHZ�9s&�=::
.�����G����R�q�v���a��[cumw?W!�7J��.i*����ﶉ�)<x��� �R��y�e�,�aii)Ӡ)��-B��TDnh�>�+4���⸶ku�!6���>b�A��U�L��G��\P�-HU�})k�,a�tfL%1���tp'�B!�Y�i[Lz���&�X�9����Z3��I�_C���/\��������!š��9�$����۷��7_B!���g;y����bҽv�H�G|/^�����<����O��v�f�|�ܭz_��˹��|U�Z�)9���g�xu[�2Q����3:���[��������|���U�sP(V?����~�:���?��K2����p���k��ն\۝q��yqum�[��mn~[�oC"����
!�T���8s�Lf�A���L\�3�
q{�#��5�_k9����a~n$|�?�ݻw{Ɣ��]�a��[�{���g�9(����<@2���q�0B!�R�����%�[�9�P��5C���j���1�#[�0�[��".��+W����333 �������hhh !�s�݃�k'=BH%s��U|��=b�Y�g$|�oߎS�Nž��2�Eǘ�! ��VTKY��)�ڡ� �g�������F�:�8=�JT�_�ܾl�5a�w�A��;2�X3��ﳾ�D��O�SђpD�����KW���umO���t����� �v�u&��Xw�8���>sS�Ӹ~�>��CB�,nܼ���vu�V1\�u�TD�K����
���E��N�h��V6��=_�E�a<T����2��}.Y��҂��!�B!�Ƀ�$~�^%��*~K���J�n��r�X&z����uㅸZ���}�]�p�q_w;
B�cc���CGG���A!��زe�U&��@�I�����E�͛7�F�&~kva����׏EU�f#��z�1�}R�uºs|�to����ӱUHœ$�!�Pպvq��MRً�)�Ca��+cm�&���FLZ	�HX---��K_?���c���cma{���[��pmw�\۝�b��rr�O�Ə?�B!��֭[�Z�ᚙu;u�Ƶ�_���Jqm�s^��p���++����1X����p���f؝�������e]K:Vqkh�B!�BH岚4�ھ��Z�v��ʶ�y�C�9��V(#��C?�/^��="��>����x1Џ����x�o�BHeq��U����A����.�h(�n�7>NuFk��Y3���녩u�j���c��6�oEr��v/(p���Z���Đ�[���%�Rz$[�ʐ�z���(��զM�p��y|�� ����������Eumϴ���~�9�D�n����#��ڮ�ƾ\�3�rq����,N�8�G����$����cW�_×�~mk7J��U&��~b�	�5�T}iƩb��p
��=G2�	�;v��2�A����ջ�d�-9eMbI�S�Ñam�2��z��;!�B!��r]���`���f8����s?"�,ֱ��6��ʵ~(��jjj������	LON�c3'~������c�8y��!����ܹs���O�����gld��3 ���؈K�.EZ,E�Q����=w荵���c{���U-��#��=������2J�7ð'�d����55;U�����F��^�~���)p��o�|����ۨ��˶�@\n��\���vC�\����hS��u��>���;��zWKP�OA�^$�?4��׮�?��?�B��F�={b�E(�k{i�tm�3�Z��=��A��\�,N?�e�$��{tD�V�H6����u`�nI<�`��B!��Jgp�[�IW�Pe���:W~N��-�-�1��0݉�
΅k׮]8y�$~�����~��/�!&��8z�&�;���� B!���4��a��b��Y'H4�U�6oޜ}\��A=�5�t�Ϛ�l�m�S��貚�������sB�Kc,/(p��Q��-X��T^�r�7�C��ڮ��.ITم��s�HI��W��~=�8�D�p�3��T��Va��;�urW��%m
a���zn�q���nm���Rk/��S���O ��1ٶ};[�1�ە~L�v"r_�u�8U_�q�X?��f���xz#�Pi�
�q�fқ�c�9+���Z���M��K !�B!�΃�q��*i�P9�VQ4wn�X�B�cE��^�c	w
ܣ��yN�;�jO7Ri|��W�}��{�]B��ܸ}��1�������^�h�|��vlj��9�e�l'{���:&�kcFzu�ǣ����X�nY�8��I*���ʍ!�pf���	,G��I&�.��ڀI�W^yǎCWW�������%������Ghjj��MMN���3WlZ�G�n����&q�����]]Y���:mq;4�MNL�ɣG�P�y�N���_����S5��u��&#C����M͙�aۖ�X\\͑aii	��ш�V֮7�:�n�a"�+�򽟟����F��ƣz�(����9�����!
�|�b����Ey�WWWG��#����I:|���ct>���E���	�ڃ��/�/`d`H+�Ϗ���}a�����K�a�����|<��q��E����C�*��U__�.����7�����Q�13����)t���M�Ei�ʑ��6mںvSB!�BH����Bk�&,�Ϲ��b��]�9e]�\��ܬ�X�T$�1S�!W���6���?��?�����e�����W����U<�|�S�O�i�E!�s����_�uTB��vu!�J�o��ѕ+Wʪ6����Cg�����83^wX��ElK�f�N����虯�n�l����� b��'�����������^Du�7n��Ӿ��� ���³������[�nͶ��ա���'��m����U�׺\����l��D|
۝m��%�F!*��ԑ7.=�U�q:�?ѿx�U�����֖Ʀ&4�����5�g%��_��&>x��P�QN*�OM����;*�{�ｘ\ ��('4E)x��q�E=�,���D�������x���������GCs�4F{▲����g^�[�N�R>[[D��x}�ucSc�X?��oU�����ٿ�`��u��j�
�T������U�^4�{�8���y^b�������R'��Z�0so�qiQ��wmw�mIT+�I�YC|7��:!�B!��O��}m�0#]�YV7�������k�"5�Xg[k
�8��\h���ɓ8p�@��D�ӢB�R�9G���w=y��E�&�{MOLF�W������,j뢑MLON��i'�@����I������ً���qP(�OO���Q &{���"�?��u�hff&2��(_�����f���龣�WG�ދ��0UQ�ϼ����o�78j��KKi��dD�
G�;u��l�~r�+��mog7ZZZ������{N��G�}��}ٿ�8؋r�z�ˌ�UR7�cV����I�)k��CО[�-�x��$?���/ëػ�Z����ڐ�1�OPْU�$U&�S��:]���V¥����m�ė����s�AT����;�=ë�_�����'himŎ�;��Tn�ra;l���vK��z�f�]���wm�~����Giq���һ�[�����?{z���!l߱��}ss3�������_�ԈH��+LĄ�(����Ć�6DE��H��6��>��Q��"	->�����k��bBUT��$��;��؎;��ц��zt4�ɺ�m����Ԧ�o�7m���� �����Ɔ��;Ա��k5|(��؆�����v�4O@�ZU���d
ɵ�����yU��_�de�(���п
�y]�~]��qpf~��o�xٺ��_g'�����	�2���9U
�	!�B!���:t��d�>����+J��C[�P���a�%����V��K�-ꆿ���\qQ	�L�IT�CAX�]�s��lڲ9���م}�"
��ж�#m�Btv�ȡH�^^\���8v��'����]|6������o��_������NOv�Sؾ)���(_{��������UD��E�xtt�w���~�ܹ3mQ���OL.ؾ}{$�G��������_�/���q�5�߼��	TUW�csD߷��G����pZ����}�5>:�񱱒�CT��B��ؘ�����"�EV6FmP���U/��f�w��f��f�����༐ns��|P���ܾ��S��v�f�ܽ�� O����_G�&�N�>��_~/^� 	���|�����.'[�v�8/a{�5�Nw�_a���=q�?|����	������/`�� zϞ=�A-!��򦩩	5uux��ܵ����ԋU��5���}	�5�T}iƩb�ܛ{�>�$D��֭[%wS�S��:�0Q�:�e.=�tWt����B���d��9vB!�B���X7!�����e��k��TW{�����Zfxe����ʋ���~��߇"�%n��>���A��y�s�\�r_ݹB!�}���o��}����S��qㆴ�k�������s��V�,E��1����h$?���bM��:�d�-I%)��
����$��%���P�Ф����7����˿���X���O?���\�*s������jm����S�i��%q�#g�İl�R���
����ڮ�?4��7o���?�g�B)_~�֛����E۶�Bq�ր���rm�o�!��:��ˏ�}?�5�V024�^�D��˗�u����%���������/nwO@WNZ_���&��6m�1Jq;!�B!$��������0/]J9�Eu���=~mrg��~�������uD��s��u��El۶-�dK§�yN�=���hV�$�ejz�+Kطoz{{A!��9x� ��3�fg@����e����}T�ݻ'O����|�j��14T�y�8����LB��z�]۷�M[�<ŉ?:P�"�ӵ؟JJT��;���0h��q:��?�z��R;5���n�G��|���~���Ɋ��^<a{fO�v�c��vm׋�o�~��_A!�<�p���v#�v�j��-�����#��=�N,]�����ڱ�̠;�LP鎩�"vU��S�nYfp"%�=�dNB!�BH����fg��C��f���E�.�D|��nh��+�������o������I�&��;B����!޾�&������B!�X���#���矢eKq���y�,�DÛo������i��ceƀcP��W��2>�2�2Rr��bm���������k�ASخv���l��s�����V.\��]�088>�}�x����ۛm�k���@��|�����*�X]]EuK+^�u���� �R^lݶ�mx��'�8L�zԮ�b}	�5c�
��k߷��--.��.�QWW��7o%U�u���+D��ڲD���������B!����xI6�+B��6���E�O����X^��KL��=::?���(����՟?��CB)On޾���|BTt=}*c�����;g�e#[�����5��
k��W��{Zȶ ���=D�
�[�05�Y�v?^OT9f|�$�,�KTb�������I�1���+H4|��g����o�um��!�ǵ=ۮ-l��	��.?����m���x{���$N�>��1;;B!偸Ǻv�>��N�!��[>b�ڮ��^�O�(Z�,��$\Μ9����E�$��ߩe������ͱy.Qe��&�Z��0�GB!�B���ë���5Jw�����nuz/h��y�s\j~����իغu+���A�gzj
c##���K ����2���������CB)/Ξ=���aeu����uAQ!j��s�Qj�:}[k�~D����c򹟚������d�uC](p��T�SC6�|38La{ʲ���̑A�~�q�.,�T.I�k׮�����|�M��������H�mO�V�k��+X,��!�S.J �W�w�������Ep�R&���_��?��T���ȧh����+c}	�5c�
�彗D�n�k:?��[�n�����_�eշ�vջ�:s%���}=Q���%������@!�B!NkÅfa�53�rpW�-EtS��^�e}|d�V�1�������?�D��_S�N�t�t���k�Կ	SSS �Rl߾����	JD͓��D�[o��6�3��8��c9J��;�LW9����ִi��Ԯ�B�{�<3p�:���N�LA����vd��m�~0-��/�rJZ勿|�2�mۆ�Q�����;hinɶ���n\O�f��P=�4����u��T�����K ��+����1��w����� �oΜ=����-,J���;b�R��5�AE�J��d}�_�_
a�5��y��@�A$����	��V��eX6KBʺG��Jم�9�v���t�Lb7���Ƶ^�TC!�Bq3W���3c�՟�"w�)�Ic,/�"Tҷ0Ƣ�=:z�07;BT�UC��[x�w�H$@!$��������x��@��ٙ���;�16�r�r�N��>����^3L�h�U��\�а���wo٦�ֵ�yo��!34�ĵ=�XY^�[w:���⬮r)�\�D�awc��r�|��5i�/^�Lݾ}��@��O>�[o���\�e}躶G��36����{��^�����M8w����!�ē={����]�~��-��N\�����Jsm�B�h9y�$����������n����}�� _UM'I%�?�$!�B!DΓ�j�:�����=���Rr��1���Q.B�B�oܸ���v��̀���o���Sl�ĕψq�|��x�W����B!��7������� �<��n)��ҥK�5���߷e|l{ _[W}N���-�6�8�ч�0�6#�8���n�۝��P�9���n��#I�8��ݹ�5i%�U�G���"����Y鸶[�T�sW�D�n1,����u����	�}��NNM���C�@?!�ċ��f�:{_��ƱGo2S.��R���`]a��X��y���KÊ/l�Ŏ���OOr	�(�կ~e{���x�ee�?N��a��%��ֺi様�'�B!���H���F$��������3�R�k\����]���j���؈�7o�?��?@���Y'N�=BT,,.���'8��ݽB!���ի���/XZ抾D���
z�w�D�����$�q���S6�i�wp�isU�>k�ܓI���a��w?P��ˍhO%��\nP5�C+A��潅�^D��7^,7�s�N��΂DC���5]]UE�vG�b�J ���b��n������B��m|��o�νo{��;��G�.?@P��f�����їD�n�_퓇2����oF�V��>v�O��;Q��-Έ)G{�M�0,ն��ۄB!�BPײ���y��mm��J�)˖�TW�W�U���v�a�%���_@�aue��$/C�xi�6�ۿ�== �/<���E��/�?~�D���F����h�홱��9�E�����؆u�mY�ُ1�7�����q8��MU�Y:Eq���r�Z"ws�92����{$��
~��,$!��ӟ�����|�G��\�%vmw��+˵]���}���������?������B)b9���!�v/�!��#���E��+�8ߗ�^Va�G���,��@���ٳسg�g��tfȿ̠�s�}����h�zgj�zc��B!��f,ьF��[���m������].�Uó^hi+c�B�V�߾}�6mJ�I�h[���He�������701>���9B����x��~|��� �1��|�$:�n݊˗/��Ԫ������0Z�����f
ߝ�*���c�?�Ը��*�>�G�����ݛ�8;c������w!>���vdȄٓqKZ+��7ޠ�=b>��c9z4�8�����rm�����@p�:f�?�z9>=�S~�� �-Ǐ���,��MW%����!��*V) n�%"�9qK+��{ih�����<|�	j#��V�;�s��i+t������p�#;�=<C� �7�f����{�^�VK��ƽ�ݍ݉�vbw^̾x���b&B3!͓v�Q�>�eZ�k�&	z$  A�{W�ŭBUefݬʬ����/�jԭy��Js���s�)�d�HK*U�x��!�B!�D�^�6e�H�z㏀k܈�5δ)�R�m-&�1�'7���,�1���C��>����悐H���%�ُ��}�w�$��(iiiرk'N^���D������8ǁ|���4�2o�.@U?����^1���|,�K�W�Ⱥ�Y(pw����/n{ج����e�C_|�"wu�*�Ɛ���'�P=��6`Μ9����0�xX^�ڗ/1g�ܘ��]�M����Ǉk��\�Ip�v-=�=�^X�7�x��� ���EE(�5%e�Z���H��vӱFk���<c�v3�{Y��v#���x���9���}{��i!a�FLL����Jj���dc�IS����I�B!��ȴ�� w^��8����l�K5�W����A���a�%&���g �QQ��wa�u��U�ܽ�_ !�gٷ?.^/�#b�G�C��v�ޭ���6'�#!����7����}?+j���h+�)��)��z��Y(pw�Gi�E�>�c���Y� T��Ǥ��$�$I*' j�|̉X0Q��g��@����;����o���=�M"n���Ʀx�˖B�k{<b����b�Z[�|�
446�it#��X&M���;w�ҵb��>bM�nFDnu�V"��v�ۍ�	�vQp"αc�_��l��xc��n���i�*�2���v�����m$o��aB!�BH4��S���6\�O�5'rW�cy�5ƊD<��֭[1c�<}�����Ԍ���@H$:��PS_�U�V���� ��k׭E��j���h4�֡���9/^�իW;*\7�����:��"R�P=����V}����fL1��y�fL�}yUKF�B�*u�* tO��v�!�U	�U�b����`6~׮]����o*)F�˝��p��1LKV%µ]���wm�k�ŵ=<ބ�τ Oߵ=vQ���*�ݘ�]���<t������!��� �<|�.߼&�>'�>�8a�nl�&nE۩)��4,��v3�CCC���q�<+����is2>�9�f�T�d��2�Q��1����HB!�B�1��fb��|u(�)�b�(�+���C%F���˒��=�>���}����q���rl߷�D���gشn=�͛�/^�BHbBٔ�t<�k01�x�#�r�С�չ��x;]���5�Mj =J��q�F7X?�"j�{T�{�:�T��Xf���!��d����^����Ny���U�N�}j���B'�ڑ�mn�>�+V���r�D�����W���9��=�M"n���#��wm?�!��C�jU�gY�� 1�����<~��N�'���O<G!�~<���]w���X����ܛ���8����}V?��}�arrr|�&�p�j���w�M�,�h�v�k��e���-�`*��S�N!�B1FI� �e�M����\�C�?��?+�*7��K;̚�Xb����T�ėښ�l���) $7�����{|��mmm �����0w�\�^B���܂���d���2�j�ڹܡv���Z&V�q�WeN�4˒k|÷��l<l�s�&_
��v #����-�*JVE�K�G��{Ff�8���}�h>�}�(pw������������E�Y�|_����JodZ'�P�=��F�tc-�l�[v�5�i׼�ux띷}"w&�	!�^v�ٍG5Ot�>"�[�{��3u�Y�����0���KkS�ڱA{Ճ
gٿ���k��?>���KR��c��̩ ��J!�B1�Ǜ�I����d�f8������?Gͱ��3Ɗ���֬Y�%K�����9*�`��� ��._ġ=������!�{�:�G�ӟq����γz�j,_��Q!��}��Ǫ����FK�~�K'��D�pR�,x)n�
��N��姨�۵bwY�<��A��H�j<�1���ѣG��}��\��)����K8z��qm7gBЦ��.�í���b����q�C�h�hÑ#G��矃B�=�]���him�%r�]ۭNr���| �Y�c����(���z������ ��\߆�v��]�n[Ǿ�`eG�� !�B!��ù����3��&�1�7���R�n�^D9���1�[�F������a�?~��׬BNn.��8�]������>�]	!��CZZ��ۋ�Ιz�"���N�*=�Y�1�'��v�e�ƾ�q���h�X���$����I`�06(pw����lޔi��lS�u���4#�d�li���Zwc����&��Ν�6�ڵk ����w�>Lʞ�j��k�,����7k�=6bl�����"� ;v��M� �_���
&M�Cy��`������=ǲ0�L���=��d,�X��	�c�?W�=q�iӦaǎI�l�z�����1���&�F�I�op�m��={R6*�� !�B!�%�#؜y�(�&���ci�o�d�e4> p���7�d$�:����A����p�z1:��'O�BH��I�:{��e�ST�>���IOO��s�U�n&^YT��֬�l�^�m3j����,��vǘ�B���t��#u�%���jS��91Dsc���?��b9�ÇS��0����z�
�8�{�k�,.~��&D�m��H����v�z7�'tlooÌiӱr�J����BH|�>}:�/^�;�K|�������o�F��ٯ7�,K�v˓��$J����sb �r��1ddd_�A�K��c�*6�I*�x���fܭ��Ҹ0�e3
f�[Oq;!�B!�m}#ȟY���Ni�P6&��C�X�E��z�@���y�E���F�\�t)V�^��w�8Ǔ�GX�j%2��@�zzzp���m߆�+� �_�a坲���
���x��	��l޼�gώ����p�5Cm�r�^�6�6b�fl��o��"��Q�+�;LIS
֤Jfo踸�;a��B;1xn n�|N2�1Ĳ!p���'tR��(�??��۷#''�� ���!�iwm�d"�x�}����D�eA�M�{�n�6�*���	K_]�;kjj@!��yyشu.߸�{����?҂0�L���=����cEK��g �"��9�����h�7��D%�Bz��Q-�P�^�:$
Q����0���lp�AB!�BH,��OW���:bw�R顱����^�Okw��.#-��X%%%��$�exh���ƺ5 �(ͭ���?k׭��;w@!$>lظO^֠�����q�#����=�z�pݙZ�dRw�=�,�dq=c,��#�!v"�G��B����wy�}�d���9�EZrP{�Dr����KB$֍��DVnn.8�O>��9���q�����.����n�/c���gM�k�� ^��a���>y
mmm ����8p� .]/��`��}���/�"�޳L	����k�o@Ow7���Y�+V��K����H���m�)$j(��*!�HH�r[����sa��aޭg��B!�[S�T��+?G�zC.��0gw��X^�9�w�cEBoǏ�w��]�#4q�G+���אEwb��Ϟb��7�l�2TUU�B�5�����A<}N�#b���A�|��Y


|�H��zN�e����za�M9��d���7깷��}yW}��.��=#��E�a'���=�8/uc�$���~'����᷿���c$����Sضc������V\��qtm7ؽ�X3�?KBAo��*V�����>CGG!��#--��A���Ȅ����X���k�õ��q�χ�.B�+V����	��h�����>��M��
�V|w�%�����~Λ:��B!�Bb��u���ahpP:�Э#*k���X��|�L$�R4�l�<y2��ۇO?��9����X�v51ý�R�ش��ݨ��!��ؘ�`>�f���;7A�Y�^��{���&M
�v���>���s���wc�B�����xQ��
�]��L�1�� u��;1h��nwc�s�7oƒ%KP]]��=��z�
����{�W��k�_-�nr�k�?Ԙ�ݺ�0��?�q: ;��ϟ���c��>�%�!�CL�<r�(n������$"Q�k�p3�^��Y�I/��L3�q̿|V��.��_���q��!G\ⱏX��$�cb�CȉA�Z�4I%�{��e	!�B!V�)�H�tըH.��0w�)�̓��^n���)xx�P�j�u��A
�]@��]�<I�.߸�};v�r6� �b�3f`��E�2z=%�,�}}h��q1�uC��bm�5>�0����y�D���K5��[�m8�������a,����aT�\B]�@����
f�!~��Ē��YN~��➥qq�cݵݪ�ݲ�\1#,�o���=�|�u��4'�/!r띷�O~���^B��o��'p�����5�&�>b|��X���@��p�/qQ|/,%I��Jt��?�?�T����f��B�v����&N� �B!�X��/EQ�H���jbn`,6�	�uV~��'�1֎;�`�<��9��|.YB�r��>���!����B�1�M��U�����AH,<,-�{�x�W�n�:�E���G<�5�Wcmх�����h�KV7�����އ@b�w���gLG_k��ҥG����$V����7'���}�{q��{1��ߧyG_�K]�#�=�?y�a�����u���c�x�M��w���� !�����>|w����G�n��#ք�fb훸eQp/uV�nf�/�>GG[;222@�C��B�n&�H�����S��L�J����x�"����=/� u/�� !�B!�%u�845͜)�v<3��F'�P��l�e6�ic���4_�����>��T=x�e+�#�.�$�_��;��z�Utvv�BHd�L�����Q�NbF��?��FF:%�Ns��	��-L�b_�YG��S�z�\?Ԏ���\]w����t��S�j^M\B��$LI*�L���.�7e���n��G<Y��s�b���x�"�����slݱ�Yِ���F]�ÿá��c��ܲ��&��8pm��3����A'��!΄#���GœG���R�Z����d'3A3"r�����'����`Μ9�����S�$��D���&vW����\F4c���"D��B!�B�!�F��)����lX�*Əh�����,3�R�b7�J�(�f�������~���.�Utq'1"��/._���{q��	3z!� ??��n��ۉ*J�3<L���dff�СCq���p�j��6��=l�x�`�P�f�j7P7̙:�&��«�K��rG
�ͻ1��F�n��T2�����#��D��}9r�w ��.\����7[��ь�{��%����>�X˂6;��E���_(��^���o��6~��o��&�����h��P�&�>�lTn&־�[�?~��f�����>�v�<!]�,��6�x6��2�����ɕ�k�����t�U����L'B!�B�u���=Ҡr��C"�%K�kW�JM5n�����i�������vK�,��͛Q\\�,B���k�"3+��E\��~yGĹ3g���B!j&M���w�ԅ/b�"��+�@�g׮]�={v�'��ݧR���Z[�Yo���=��ڃ��9`��:����0�`:zۛ�UV�Ė�j܍A��/N$����;�����A���>����|�D��܍ݨk{�
~l�[��$�wܵ]�5~�fD�C�x�X������o@!���;��--c-�����eYDn��e�����In���@�;�н��eӏ;f)�V�v�x�b3���%�ԛ7�jZ'���$wt�R��I*B!�BH|�Y7�]�)���?�OQ,�_c,_@�^	���=��N������V�_BbA\7??w�����@!�Ovv6:��ϟ�=?+�%�i>�Ę��ѣam��cmsbZ���u
ջs���5C��g1��vχx@�����E��^Z,��Eqc�o���ɛ��S^3�ѝ�H�X�����/~�؉��	!������$F���O~�W������>&O���P[G��e���g0'�3AA[ͳ�x�|������Y�������756���I���Ϫ=�����:;;���S8�p�ɲ��>G��]U�H0���I��Ku�p�;ݿpA����mN��g�ZWW���w���n��_<kh�;w.N�>���n���L%ikknAEY�$��5Ȉ�|hh�����}Í������*M���������6<�|d|��M�ZZ}c���\�k�}�aY9i�k�S�ց��B��-\�0b�[� ��>B9)�#c&Q5���DLR�%��\<���B!�B�E����NGog�����M��#c�~
c2��ݯ���?�3���@�%��>)'�Ă�}q�<�3�N�B�_����~����cuM2>�����G�A�gƌ>�d���ǘ�v�x�`�Pk���F7�R��s���@�3���.�F�0�MN�]�<Qnj9��DKq��B<����7�|?�яl�U�����8%v����I�����~�k(�2E�.���/���g~���@�x��x���A����Bܾ{�^��5]#�Bܾs�n��j�k�����.^����	v���:�����N�BS!v�9s&�����X�`�B��-Z�H�����m�ԩ����gw����&���ů����.�5�7o�#����aڴia�۝�����������U�����"��r��@OW�o2��ysUǤs��&Y�qq�㇕X�|Y�8�n�=ߚy~\Q�E˖�}�ZĽ�l����z��7�|=88'�'�o��_�ͅ{��-R|<���86��KT��+]�ck]a�d���]�WX  �B!�ďo>2=M�b������*V���b%&�[1�
_E�}�V��ǤI���[o�׿�5�D�E�NM�w�K����6�G.�~��Ήk�=]����Bz�3����v<��v�o�����C_�#�;�مA���|u;�͙�ǌ��D7g�`��N~vq��ߩ�8�D�fE���ɿ}�ϩ��g�E-�����}δOC��N��ă�0�r'?{�������@<�4�N�1���8u�{��T���T�eJ�kH
kn�g���rc,��WR7l����.��;�;u:��[�&�B'�|v��p/��Tcn)c'����b�,I(��b�m۶�ҥK �"�O~v�'r�㕈\�nx�b-��M�����-�M<D��_7&�[p��ߏ��|��������'>%���Ğ�{Q�܈��F$�>bM�n4־�H���f9v��#�T��J�N�c֬Yؽ{wB�Opy�"1h����OTI\%����1�x�����Z&�!�B!��v�5�q��fp�S;�[5�R�����D0�:q�>��c[�s�D��Dw��n�8@��\���'ǭ����ȟR0:�wȨ��ڰaE���G[Kf)�B���=-3�֯GZjjPl�H��)��D1�͙����3hr�͙�9՜9�(d��/_��ٲՇ��{q���O��H���.����/�c��E�'���-�H��Lu�z��gOd�BH��uճ�0��/�Vp�K����}��~�1V���s�=�w.T3T�Q��1�2c�%3��w�>���
�]F�'�<���'�70{D2�Ŀpc��%n�#ل���w
��A�����0s��O�H�����kT�gYDnB�������Po��E�v������x��i��W>� ���7�$�!$шg�����Z�Z�1V'3���X[�#���m����H�W�> q��+]��7�|T@خ}#4&6����0�N4׌ս9�@!�B!�σ��������A4Escu�ݱ��v��}�c-[�7nĵk�@�E|��K�cˮ �
���y����|q�#4Bq
1�c��=8y���Pz�$.5Hba�5��q�ڳ>��-��c������H�ʺ��u���i�9/(pw�j�ؙݍ!|�A���	-Q�h���<�"�1�p����}�۷s����"%�"�ϟ�G|���"������n��ܲ���=]�#�
��Gϟ��w��~�{��;!��W���#ǎ���J�����o��C�v�N��Tzx��Q71B�0?~ܶD�'\*7A��U�1��2�è�K����B!�:S� ���0�
M�U��KV��#�B�X��"�����
c,
��A͓gX��uL)�
B� ���;��{����/���B����cۮ8}񼭫Ӑ�CKc�^P[��F��mf�k[<�kfjC�P�ި�=d�%[���0��z��n�Q��=y`�0~P��2�G�7w:�:[�KHg�x�Dd'�4Y�I��<��#���}lB,"�U����@��֍�س-^�x���k<֨�]���U���vƙ��*�4k�%�?�����?2aE��g��G��~E9:���޷�>a�n�ν���ͪ�^'�i�z<��}�}x����I���͋�f���LK�GNRi7�n�J6F��3	����Ƽ=!�B!�D�f��2�jW8��]5~�*�6c�hE~c� ���1����x��СC��w����z�)�[������k���p`�\�r ����ԩS�e�6��������xp�v	�;5�]�v9^L�˻�
}�f�*ǵͱ�c��� n��O(pw!m��O��.�r����'�dN�D�:��U]D����h����\��%|�_�?��'��݌��M��M��]۽�8����nQ�nU�3� ��{����'x�����Ą!d\!���@ɃR�h�V�zIv�v�����Ǔk{�����3���n@�W�;�fv��ٽ_�{����х�z�*��^�|<e�A�Cj��}Q�N!�B�����/,B_wG�^u�g��MV�OM�P3��� l�ceff��Eݐ8O݋Z4��c��Y �*�y��8�{/n_����fB�x���k7����gm������5hnlqo��6��CR�d�Z96�dm��@�z��,���Z]7ND�����	��wr�ދ�Y��=�|�"x��$��41#t�_(�N��O�$�Ѿ�Ν�={��̙3 ����c�޻�UkV�^�um���ܲ��h_&�tm������̇�U8|�(Μ<���6BH�#�m+W�����>�{�#��!a�{��i������6���,\�;w�t<�����;�skfPjQڄ�j�\fp,6�2��Nè��핓�	!�B!�ѝ^ xZC�Bc,�8�;6�78�	:�k7��ϒz!����X?��}���)�y�<fZ�C�q}<}��n߉���h�X�2�����kW�&�/Ľ���� �@h�1V�k~n]��?F7Y�ea� K��sPgn�%�`��|>��m���������>�f���=����y��jڵ'�p�Ԟ�A�g0����,nLB�9^��:{�3��o~�+�����sF�&D�m6	�-����(t�*�7k������I5>��KW���KBH������������g�DVV��ݾ�����5'��X����:+X����[|&v!---���.�ݯ�$KBA?I��믄a�A�ds�2�YY�(m���B!�b/��S�.-4>���YR]1�״)�F�>���-Z�l~��y��hk���O�p�����>�{z�C��ւB���3�\x��2�'�+����<�9s�D��K�ﾌ�{��G0�VL�����by|����zz���ݥ��NA��Ew�G��tI�~1��+^+/����$�ō�-I(3���%K�����yZ�[p���ڳG�M"r��6���{\���&�k��}���'��q�fL��B��RBH�1}�tlܲ�����s�(X�	��X;~�X;D�n�|K6е�-��������`u�������n<Q%GZf0l�-sb�oƔY�42QE!�B�������K5>��_���Һ�̥��XƏ���ޢ��Eܿ]�� =��?�_��m7#7/U�U ��de��#� G�k��-!�bhp���jS�6���g[<���pիmP��c���jc,o�q��n�?�mOG@�G{.�����A�l��B����8�\VA��6Y%�I��%�G_a��I(#m����{����m��᷿������h5#"7kB�'�n�#X��+ݣU�[��b�~O�?��EQ0� �/s3!$yX�t)�,[��7�����9f]���l�-�,
�a����"n�������(,,�N��]����*�P��u�J_�.KRyu��a��&����Q�)Vʠ�;!�B!�~z2��v����Fc,+�ݽ{�����ӧ ���ׇʲx}�*O�o^����M[6�Ƶ� ��dc�ƍ���͒; $ޔ��bp` ����زe���D�C�S�G^�Y� +�S�Q����q;�q�w��50�ܹ3��������_^=5���C���\\���$2	e�~�ڄ;�~�����8O_?N�:�w�v���0'h3#�7�=��{]�-�e�g�����ô�"���[�㧟rb!���Y�ٹ9�~�V�ͨ���}Ą`�L�����{���!����_��a{ .1�.��DL�5ow�]��:	j�T��������^�8Z7IHP)��9��(��r8!�B!��ō:`c�W�����>''�]���4�fcb\���|�T��c�+K1)7�ē҇�X89�M�fHI�s˶;PS�5�/AH����FuE%�{��W�6�X��5?{D�!�,���ߩ=\'nY�&l���7j= �w�8��O����_|?��N�HM�8����)^���T��3����D�{����<ߒ�?��A���3g�}�v̘1C�nYDnP�����x_�tm�EDn���ٵ]Fsk�s����C���;�B�Ȗ�[�34���I��#���'�eJp/�G��6q��� ���;v`Ŋ�LDّ�
806u�1�иX�̠�Z+
�h&������ENCB!�B���;�ɋ����]��.��V~��yB�T�X�7FSN2�1����w���Cttt�8���������[AH�yV��=�8v�8N�<Ś!!��ddd`߁��q����A�ܿu�7V �@��,V~o�W�⵲V��������(3���L�u'�KVV�+���j�ws�փ����ur����OXɜ��5#��&��PF�I�v���~�A�K�����_����#�fYDnY�����{]ۥ�1�#��u����C���W?���)��\Kq�Q���C�z�-�-�6{�#��D�v�G����:\���.��� �;����1����!a{�g���e���#��x����=c�8>$�B!�$�o2=-Q��'�j�򕮴�v��Ke�%q��7Oc���|������A����'X��2N+!񦥵�/���c8w�,zzz@!n#77����]����A�4����������#''��Q"�����ۯL�ѸeE�!���F��ZS��Yu��~h2X7�
�]����Sg���>b�J���'���a�����8�zÖ�H�$�D����o�>�:u
�<,����X���w����ƃk{X�)�[���iFh�?�wE>��	���@!N������.-AOo������{�(����#Bw�����OU����K�b���I��2ۗ@��
��D��I߽=4��q�,c+&���
����I*B!�BHb�V;��y)a�LE3����+]	S�ڡ�M�E��<����������A�G�ݹv��1=�#����/N�о}�}�Y3$����ӧc͆u8u��y�;ㄒ��A�Cvv�ou)N��}Lr$ZW��C��[��Ħ�𦥥�z-�vA���y�7	Eڂ�$Aeĝ����I��Q&q��dIBY�_�N�>�Pa�̯~�,��ː���h5!"�,h3ڗ5�^,]ۍ��*���
l߹�e��� !�8�̙3�q�f߼���g?����k�E��)���XcǤ;�\�ܽ~�Ͻ.C�*%���̉(#}�Ƨ�ve�JyA���uAol�ua��2�G!�B!��3�E�ԙ�io
��[�9��;��"#�/^�={���ٳ �����% ����乳صe;�rs���cB�ӈg������� �N�+*����:�9s�8^�K���\���\+��:4.�7�RQ+4�J��I��0�b���;���%-�k����w��ܣ%�����;Q��x�NBE�j_[�l��5kp��]w��ڊ���Б#0-"�$n�&X��ںQD�V����x�={���,��чC����hV�\��sg��kWl��X��3u\��Y^M��'��cǋ��i�c476�����;v̱���ɱ`ZJ-l�:Q��k��v���ݣ3�\=��nc�h�t�!�B!�$���y���'=]];4,r���2�:�{���z!��Bm���.����p>222@��k�ū����X7u
�ܢ�-!�96oٌ�����b'��(�{�=����h�dqf�kw�����M!n�]��v�&�����b{֗3�+��w��=�2
f���eXaݣsb	W?�C]��#:1(^+/�����b䶄S�m������?���QTT�j7%��E����`݌ͭ"r{�����g��x����yy��W?���)���@!v#��v�ٍ��N�,�c�c�>���wjJDn��-3�e��!Bw��]044��;% ������ɓ���$t�ǅAo�_^0R�J������T��&Q�?u�R�N!�Bq�/�p�0#�=NwL��*ꆱc�j���Ac�H$��=Rێ;|�eee �  �Z�i=��;��0w�<|��~��BH����ۇ��>!v#&��!q6l��u�\&>�_���S�5\�e�ʺ�n�Pn�5�̬,ܩD`lL��I@EG&�y�GO��,c�Ɛ�
$�:��׏�,3�&{�6����uuu �@<D}�?�����l�~�,ڌ�]��n&�k���ѵ��n�а��=��8�֛�|�2�jkA!v�������Ni	�::u���V��-��V���#�c�*�wZ�]P^r}����&D�Z�e�I��D�ڳ9 nW)��^mJ#b�}DW"KT��v�N��	!�B!N14dO����z���Rǹ�t��HĦ�b6Ƃ�f�+�E�ь��x�wwQ]Q�E˖�`�b'/�j��юc'��ʥ�hmm!���ԩS�e�6\�z��|$!����Y�w���������g��иT�0 n����uEO��u`��B��]8�F����$��q���axpP:$�r��U�%!qf�z�'��Z�$��"�Hm����dտ�˿����wKP��._.0(h���n&֭"r�5a�u�'�mW\oVWa�����b&�ܾB�7���Ǫ��q��˄�V�#�'~Y�'�e0N/v����l�@��Jwq��!��&�M&�H�{ ���:7�cTqr14N��kU�uΞ��B!��7�=ãc�C�X�՟哂�b��i�u��q|�{�CSS�;��;Wob�у �nz{{�ǳ��e�F�44���
�b+V��܅�q��Y��Idb �gw�����e,X� ���O��_|�
d����B��x��[h��0*��G��+�	�I�H�tx����$Kss����. ���6�̠�cPaJ�'���}��_��������|�����_��A,ڌ��ڮ�}�D�H������>m9�3�O�����o؀Iy9�t�N�U�E���8�f�\ۍ��t6��nHݾz��3�!�_�����dqF�b�?�m�ra���"'�d	�@�*�p��!�B!�8˝�A�3k����-����X�6co�����'���+�{hnlD͓g��x!�q=�z�V��;v�ĕ˗]��%��ĳ��m���݁3σ�D���- ���?DzzH��&�{��d�uC�M-n�b�*�Fwo�7�
bi&�O��Ei��vC�{�PҒ��F<a'ˈ���������� �r�^��()1h&RR�/b��VPP�w�y?��A�CkK+Ξ9�c'N�tm�V�C���#p��ܪP�L_��S/��Ѹ��fL���WG ���?����+b �w�>�l�CՃ��s"�k���_�E䉼g�ӋuZ��b���Ghn�ۘ�عs'V�\�x�I�����jq{a����D�J9�V%���8\0z� �B!�'�򔼙�4ר풉�ac��B~d�h�X�#S�<���~򓟰>�2Jn�¬�����	B���
L/���o����g���B���L'j�7��AKk+I�}���.��(**��o��*��5G�bӠ�*k�Z��Y�v�)�:�Rڔ� �C�{��m����S��nԉA~�z��jf�A�����῀(�S\�p����׾�5�����e���$V�]��s愽g\�f\<h�>�"rsBI#���M�k�n1�3��ׇ�G8t�0J��Gee%!�,�f���-�p��m�Ȟ/��Gd����b�pm�߅��J�v?(�S�.ĸ㣏>
k��9�	;]��*�vu�*z�J�ܮ�T�������B!�B����t,Q
�u�a���f��]%nW���| ֕�RR�/b��6e����������e�)��-�@H��Xg����޹y��� ��X�3w.V�zg/]��0s�$��ɂC�� �BL�����vS������B�H�uB���R�Ľ}dă��i�={@��$�=m*�=m:'Md���M���*��ܕG漰�,V��={6�?����7 �A|������_����k3'h�C��V����wZh��߽�Ǐ0o�"��lN~���zL!FX�a��B�ɻV�#&��c���g���uZ��a{���o�D��]�Y�[�nE�8KDYuaP�ݵB�p7�do�I+ɘ;�p6�A!�B!��Q�kLEO��K�V(_�9��]��]�f�ө�j�,7�#�Y!0A�W����\Ɠ�GX�x�fL!�b`p 'ϟ��u�`�ܼy�b�l�i�f�>O��x�$���:�<y�.rss����#%e|�ڍcƠ���b�L��;�G2�ҚQ�O��gO�K�'�/F�'/E�̠�Q.������BȍAv���Ag�1*�3�L.9��.����1̙����ӧ�y�:�l��Z�v+�v��:�	����õ�(VcM�������|_^����zB��y�سw/TW���$ª�ܠ0�L��ޖ��E���+W�G����5O���1�Њ�$c�����̱�0�O��{,5(OT��#{�g��!�B!�;�)��$]�Z�W]3��*q�3o�%�xʜ�̗,��xc=z���oA܃���}��8꫃�H�߹���g���c��aOO!$y��]�UZ��f:���#�w�qr�y�w0mڴ����b� ˨�=��9�{u�J��l�g��VL���IDϠ�
g���^:3DZ�OKsn�w��KR��D�(��jwu�j<��#�-[����ǩS�@��'��5��X���U�Dqm׏�*�4�+y�D�N����(�|��֣��/^!�hY�|9�,{Wnݐ��`�>�3���NM��w����>�$�y��� ��W^�5ܓ8���=.���.pa�*I��P��_��/(n'�B!����^��AX�=�)�gtKS��,Ky��*1�(�!c,_%1�'�1֧�~Jc,���֎��X��� $�445����m�&�44��� �=����-�]7�Z<q��J����.233�կ~U����2��ޮ�!d��F�*Ǹ���X�U�[jj
�׺��?^��=�x�3	3��qcО�"i����|/��.]zP�:D
��qɐp�������Ӯ,Md��������ڨ��+m5g.6a��^㟕���c�}�׾@���x�+��_�]BFIOO��{��ՁKׯJ"��G
���&�>bQp�����(/����Nw!��(����j�ō϶`jʰ�]-r�sb��̠*Q�k�d	G�B!�B����"w�,��5�L�t��v�1���?&x_+� +P;L�G`�4Ǣ1���bϞ=8{�,��9�� /?�$q���W�,ŁCq��yB�Qغmj�p��y����,�d,7"V�Z�p!R\^���z!��+��������^2��G+L�m ���u�DA�{�q�n������`����L��=�DMU�R	&���v��]y���q��h0�%����_�[�nEqq1���u�&�oڈ�sd�.Xw��܍�{��;-44��>����щήnlݱ7�]�s!�Y�fa�捸y�.z��4�Z��X�����>bQp/u�}��*&�܉�V�8qnOR%ąA!n&�"�۵n��=����6Q%^�}\�!�B!������(R
�5�X�L�B����J�fGc,sm}����W�&"�\�s�v�B���q5j�j���A�=u-�� ��ٳgc�����������ϯ��������HKKsĽ�i�{�`�P�!�]=���y=��a+>k�uO���DA�{24i<��ԅw:��6z�S��cnju�*��+�,�"%%�NVڄ��իW��r!?��O�������3�bM�l&�����E�����~ݚ�эn��L���g/j�_P��[���3!d� ���m�oz*.^�M��*"�����5�v�2x z�f7�G܂�7ݸ|�I*�"�����׉H 9���B{�
���#v�NbJ7Y5�^^��V�\!�B!���[�CxgV���B�B��\4�{�A�ܹ��X��6l؀͛7�ڵk �O=ƢW������é�_`ڴ"̜1uuu��#B�C<7�۰i�8y����y��-M�|�F�*Q+W�tA-Ͼ6-�1�N�*Ff�5���>�[[7�5���srsq�nJ�,�
ܓ�[�X�ꑞDF��*���RS� xe	+�ɪNb��$g�hۮ]��v�Zܹs�]tuv����~�#����(��(׏�*�4g&VGi�H�v�ۧ��]�mj���D�Ç(/+!d�3{�lظ%�eh��м�ዛ��`�����@�^_�"�:)nO���������V�1m�4�����9 ��;����1�9��O ,Y�NP��T�x��)y�J5�k���<��!�B!č�:�7w<-�U�QE2����M��KE�ʣ�8�B�1���ד"G4�(�y3��¤�1!���I5�L���Ǐ�ڕb����2q(**¦�[p��6ZX�!.���ew1��Di�dq�-d�eDܮ�#�̟euC��6l��6�L�z���$��˃������=l�H�tr��	���0�wJHuLX�/.�3��III��S�m��o~�����W�`���X��rU�U��u�]�qfbM���n<6>!�o���
3f��{�_��S��=:X ��?����];����W�H"��G
���&�>bQp/�ݕ����щ���d�V����#///�:Q�[���GPЮ�h�*܅!���ޘY���2��p�Xy�.�B!��r�)+��|�l<$��׮�po7c���Lc�`�pX\�f�޽�.�q���ؿ�8M{{�ϵy�u�N���K���&!����͛����;����D&���cxh�}�U�7n��"���m�q%$��fo�ڡ|�T7���s�(K�jo6���$qP���4x� ��<z����KT�%���w�M<X��*g���X�7��T��$g�h�޽{�~�z�ɪ��U����ɾ����?���dggc����&��ScF�,i5(�.�}�}�b�pmׂ��^C}�[/������4CǪG�BC�g�}��8�&7����{���1=�y�������A������>4����N���=d:��D�ۋ��w�'?�ܹs�_0eU���^w,^[}oD|�~�G��zrL�"�'3��x|�|˂{���H��Y�C����^�v1���;y�{��\sF���嫾���YL�Ϸ����|�AR���+���x�0xF�v�dU`l�5e6<��B!�B�͋�al]8}�ac�Hc�HYF����BE�04�U&�1����K<��,!N#�7��F����� ���������B>v�n�D[G;q��h��qb\�o}+�M7�ڼ�-$nW*��Q��d�MS/��#�b��?�O���'�'
ܓ���L������4�D���:2DXrP�.�I#P��ĻM�ɪo|�����D��p��X�����I����_��~��_a՚5h[⩽�c�]�BCsar�_cC#���W4Y���s>�&�(�_}�&�F���C_���Ի5�_3����f<,`h���f*�;�|b_%��1);3f�D��G�������a���)�K�S�&�����	Ŀ�D�ۋ�wuu9ҿ�]|�E��e}?~�i3fh"L\Ǥ��~����������1ԻQ��{fwW7�^�F�ܙ��V��������z75�J�w���A��I�^q��_ i�o@��uю簀��)��8��dF��G�½=???�z<��cuaк�k���y�0q���0�f�]K!�B!�5e
2=��q͈'�_Q�
�+��cj��zZ@�~�n��ٶo�>������a�W��\��_[�I$⻘�����Cff&2�2�������K̩��յ65;ҷ0g���v�'?������ ��.��I�c,�� s��CYi��n�f�:V3w'����)����S�]|n'��-��N���N|ޙ�f���?�����z�"����;��u�H������<������N��N>ߊgz����/�v7mڄ����ihk���HY���u@U=�#��j��U�Eݰ~� �&
ܓ�!�Sfb��VZ��s�S%�Kj��nR�;��ɇ�9�M��G��x��/]���݋ڿ����i��x��C'It��e�{`?fΜ�{�p�"X6�b����q�f�XSn���vE��7o��˲k{�����X�h!�Ƅ[�:��;8���nX5N�l-�����X��5�~�5dێ���_8w>�I+��y���)D�ĩ�����z�ԩ����gw����&��� 77ב���W��/]��[70���",ze�"��}D��:q�l���T��
潦�C�8q���xa�����X�u\$j��;0s����K�DQh΂�p
���E��uut���b�@�ĳ����IN ��k�X"�/**»�;!D��mr�2{h���'����n�:��'NC�S&�!�B!���쟜�.�덁d��ʓ���ͱ�c!4nK�1�Q�0����QRRb���b'p�o'��K�V�j�:ߪ���af!�"55ͱ���=-}b~v���v���E}����i�V4���EM�-����+8�����E.۩��^g���2�q�ϙ;��ǵ���ى�ӊ��{���D6��n�\�T�n��G�ו�ܷ��W8��}������ʱUJJ2��bkS�P��Ɵ��a�X^hM�e��X�U���6=�^�n��'1�Z��J���*wo�IpcP^ �\��v�z�.�nqO�c����g�g>7�Xl�^~��?�G��3_b������L��Gp5֦�jE<hW�����YEL��'���ǻￇ[7n�ٳg �����BlݶO^<Å�˒�����ucm���\�����	���ĳ����:}�


��'B�J�_m�%#�0����ܽ=����PlM��x�B!�B���a`R�l���E�J�4�X�X��5�Dc�KoGmr���X�r%�޽k�����@��8�w@ ����
��.Ƥ�I���C�CF-�Uu�8�@_?������t��<�^�U�cŲ�غu+.^�w�q�b=y�d8������0fMN��g�Y����_��,V0u��9�{����[P�Ԉ��!=+٣my��������t�ã�����	�����ֽ�<��F}����V�x�v�=_�����m`B����s��͛�����o�&l��K5cY=c��cfM1�h.�[�aBC�{S�:�����6sDof�Ȉ��.�!U�Ơ��f����2��҃���-vɪ5k�JV����щ+/a���v���Ċ�-
%%����֦3�N����	֍��r�]�](�|�ů��UkV�����܄�!�;v�@Jz.߼��9o�>bP�mUDnq2�~l������du�n���R�6���1Q���ߟ���^Ŧ@������ubso�_�L������B!�B��Ҏl,��)�cV~3��q��1��6����׾�sqO֜�x�v�u�߲	���Ux��)��ځ��V����B܍xذqr��q��u�ĵ�D����n�q/v���k?���ǔjc�`;�S#��)�>c,Ot��h5Ļ͙�GAw'��=�iB!�=m�Y##U�qii~��r��W�Ƞ��KP�(]��	�ɽ�*;X"(���r/�X�t1.^�{m\�,�]ۍ�o攰Ghh��5���j�}�����a���ϝ� �� ���׮��ٳp����$Q�Ms���u3���gY����d}�kkiEEi9�{㇩S�_O�v%�a�D��P�,I%OV�h�T�IޢM6N��܇�U8�.�B!�����i����KU7�3�
��\��c�Tc��v��A���?���L܇��<yT����A����_bƴ�8r�*<���O@q.����v�=4��p����z��U�O\�ƍ�}��q)j�ަ6����m�0�s�Dm�f���N
��O.,'�;�I��a��)]R]�D��=#�H�%�RG�Ґ�ٍ!,qHP��B�<�@'9�U�L`�d���d��9��[�S�H�u��<��{3��pm7J"ŋ���b���E\k+?BvV�|�-�|�ׯ]!�9DrJ�ۅsJ��:QV�#�����w1.X7k��j|B�D�{��q��˾{
q'B���$q�)����R��Lܮ��
�޵������� ^2VV���vK��@!�BIFZS
��i������\�}uDci��������!i�K����<y��o�!n���	��;�W_Y��Ǐ�Zq1���@q���l޺/�kq��9�v�)VSC#�;c�?��?��V,��D[�f��B��@c����f�W}����"9�k��aTƺ�SP���� ��ga��f�J�
ڥ��90|'pj��؄�])lW%�?�x�2'�V}�))�#v��wĤ�o~�����{w280�_����O���(n�n��Qpo�7������X{>��(���e�1etp��{����[���!$q��Ԧ-���َW/���"ߟ]���$�>b���b�xI&Jn�Awg�{E�)�I�ͽ=� ��ݱ=��gD#^� ��}t+(��gta �B!�$)�^xpdj�aS��C�HZ��+m�}/���$v?t�~򓟠��ĝ<,}����a��f*U���jlX���Y�Z\L^B"337m}�J���i4D����6��Ь��lذ۶m����6�b��$j �K^?Ԏc�v�J�Q��cY��8��uC'��}p�1�R�'�T�|!l�.3>���M[nP����]x���0^I�8MV	w�d�͛7A�I僇�z��vlGB]�-�!�7�k�^�9���X[��h��@���ڪ�X�f.^���.�	�������� -7���v�;���nE�nQ�oJp/s�}$�h����*�2c�|��I�|�2�`{�}E�JW��˪6�z��h�v�6��b���B!���dpH�2-/#�ڕ㣴�13��1V�+�1�J�.�zi�%����o������K�����ߋ7#��7��ANNv�ۋ��6ܺu+��ل$��j�*M���wn����$����bN�p1�����Ͱ�TW4ڦ���	M�0�qU�֯*��ca#���0�
�c�	�A(p�vc����l3��.��������P@W�.���$�HII�dU,�/~K�p0�n~��O�ʲW0}��`�;D�	�K�Z��vut�H�k{��Ok����{�CO._�ā3!q&==��؞_0%奾s���ĺ�[8&��7q��}��n��$��y�*�������k7$��a��L܎��֍Aw���pQ{$�B�{�Yٸ�bJ�!�B!�$��2�W1މ0�W�b�f�Km�%��+���X����5�@H2��ۋ/.]��Y�q��Q��/�
Є���ŋ���[v����d����hkq/;w����S�f �NUU/���V}6�ޮ��5	y��9(p'�����M>A�'w�̔��7-$r�:1h��&�$ɪP�&$�NII�dU��۷o�m�/_q'bɶ������w�Y��.�[J���`��X78���%�:�o,��1i��E����:^�
��{p?<�����E
�	���<�n�:L�9����QE���H��b(6A�,��6��G�!n���=��,\����+�O����\����bw��zS/3�	�q=х���[�y�4��� !�B!d��݃M�����ݔ1�����Jc,=���X���c�X���h��r��}֜�(�>�$��u�mū�qh��(�w��� �ď���c�����EN]��$�u�x��Ľ��poW2Q��k������aX�F�nt���E3��1��NC��8���a�5+�C��ɪ���tq���a"��;C��]�'�+�N~qJI��*�HV]�z���&���'��޻a�%��\*��Kpo����=�v�;c-�<�`��ء�!<z���w� ��|B���~B�#�߫׬���p�A*�?�[� �X���G�������H�RU�u/^��q��������lU���D�%>a�Ulc��["�ܮ��
X��#rU��p��]8:�hːs�F!�BI~�S��i���@Q�c�4��=c,��n�cź�-[�����r��K8��qdff��d�Ae�o{u�+8�~J��E�K�	���ٳ�z�4�4���s $�>߸\<�j��C�a�ڵIch����Q����]o�g#��hbv�6<:��(=�ag��}��=a=���iyfj���+_�A/9�"��.�ިX%�!Y%n>��S�@�˗�/`٫˰b�J�k���5��5Ｘ�a�-V�W#�|��B�~� �zzp��e_;!D߽z�:,X���Kq񪿸�k���ݢ^�����c��@?����K��ĉ��۹�p�v٦��$���1���fUy�3QGB!�B�8��fǦeE_�Yf����3��h�5����ŭ�kضgIF*���q5^u9�X��ܺ���&B�3s�L�Z�Mm�>a�x�#��W}v?>c,%�ahe�-D�KV3��N�Y�ꘞ1�Q�vaTv�Vh��k]�=P�>��Z��^��*�I�����'�ҍA�Ȑ���C���_��z�>Q��dIV��_�%Ο?���A�����	���?(�2%�M�D�Ƅ��q�5k⳺�m׺(U/���E�,nPݟT��N��&:;;�克 ����o��������.����^�b��ڮmM�k���v�`7���d@�"��y�s�&�����}ɪ ��۹��m^�B&`�sc����핊�#�6¶����@>��@!�B/� ��gc��ቿҚ!��h�5y��O���x�R����OY�C�WV`Պױn�zܾy��� �������Qn�g��Sd��M�Ҿ��eY�,;�c���q��/���؎�؝8��L���d��93���{���Ξt:�N:��vbY��K�}-IU*�JU��J��\.?�  � ����"���G�x����� 9���b�����D��+ݽ��<���X�z�Gk�ۥEvn�3�Ҋ�C)��)�v�g3�/D��� �D�H5+�`��ۢ��OZ0��!_l�A�f����]7i%��e�{<q����*7�G���UW]%94��7��_�����/��u�"�D��BGG�e2�Bl>8�����N	�������8�4����*|�s����7TTT`l�O�⦴�7�xf46���Vl߳+���2���Vbszq��JG>�z���br�T�;r!�M�7�X��vBj��Z��tdJS0����b��jZ�х�B!�R`���z�~!?�����X� v�1Vas`Of5�c�D�s��1����u�a��p�i���@I��؈�7nD�`?>ڽ� kH���뽂�˗A�a^���O��y��g_l�6�R�墢�^o�g��a0h<�sZS�@@�W�{w���������Z,vE��R�����E^�	��)��JrcHra�
�%y��d�Sɣ\o�_�*�{�=�K�3g���͸��{���Jڋ�����|ݹ&�bm
��Mn]?��W���0F�Fq��	����?�2_)v�څ˼�!E��1���P?�ǚO���3��v�1���,��NM��4b2�(6_�#^���ε�Emm-H�"��P�B,���gv��y�Z��yq�F�v�k�z^�ae�E0M�*���'1��T�"WB!�B)$����]2��I���=G�X���2�J���X�.�!��o�=}F��!ċ�~����|���108�y���BG)f�,]�U��r�@?>ܹU:V)S�ٺ#�@��	�=��.]Z&WV>�o�fR�����M������jf�C���
������z����ۓU���=��'� &79i��&�Dǥ|��.�v׳h�"|�_��~�3����?���˖a�����������.�wYh�/�ҍ�y��m�%���k�E_��rF*6�Y-n����Çp��,)d����K�Q�O���q�rk��E��[����O�]���sy)��������[o�m�����Ė5�v�䔁�=�aKK���Q��!�B!����bv��Xq7w8c���gܮ
c������ ��`� 7��7�B
���{��sX�z�}�~\�Љcǎl��-��f��¢%Kp��6m���Rp�Q��i������eŽ]�|�'�C�,���0]?4Y;*�u��818-�� H~@�{�S2U���ɪ�"w1\�_$��;C7�&�c�)�zB)[�qbݲ[�pq����_�o�'��!�|�[�����9��`�����m׬�Ӛ�զ�^?0�.ȩ�/>��y���a�����ށ��tRP��J�>\��Z�;zXz*W��d�?�d��"r��#�ꯌ6��9�k���]m���H~#�^z�%Kb��K4e6/q���:�%�ԓ����h�*���LRi��E���aFz
�� �B!�7�xtQ=�GG�`��wFc�L�#c���?�oZ�O�q�L,^���mg�i��y���{11:�=�w3�L
�sڸq�ԧ=ul�B
��3-8�J�C/��SOa��ٞ2���z:vŔ��a�����ڡ���F5���8v���|��d{{ ͪ0��.�~�	_0&f�%	��4�*u�F�ae+Y�̈́�S�L�>]z�����	���?�^x�%�a�
�ӵݮ>�{��$`��}����̮K��a�|�{�MMM��� !^D���֭����y��؇#'�&�Y{��(�\�o�x��yā�#?�#�ā]{�����<���X�~��	�|po�'��H)� Q��o�>�-���a�RI��I��h���e�!�B!�����Fy�%�X�s;���G�~���������߽�PW_B
�ή.i����ͷ�
�M{�bdd���ո���ر}Z:۱��QR������} �Ϝ9s��/9ku�L>�^�1���C�	ݓ5�r�0&ne6곘.���a~A�{�ڹ�������ك����$�Bw��2tc�qdH�dU6���O�w��Ο?�ߴ�9�?��>>�3-�����vD�^wm���[�y���Mo�l�,�Rm���¾ҙ���'M�Խ�FEY9N�l�ɓ'A��5k�4AiyN�mAk�^�X��Xy���J-��{�)�}�ۂ�B�ZO�A[K+H�#�h�$�	�l�Ǯ{{bJ$��F�����0�1���$UM�\t�0IE!�B)l���4�ʫu�1�3�<������oS��x����(-���&�CCضg�T/��ƍ�,+G��f\�� !^d���Xy�U�Ǟ��z�K+� �P#p�ڲM�	��G��\[[oWD�]�v��G@U+L]?��M�1S,�1��}��{{Ee%>��1�o��@�~��[�J�)��~_�''��&��a�
�'A����K�4Y���TF:B!n����?��?�?؄EKc�k-���
%��R��v�kW�����Ѷ̶ɰBQ+�f�oZ��-�^<*^��S�-R�왳���##ؽk]H�!��֯��s18<�ǏH7)Q�>�bi�Ϸ{�g�<b��e�v%�N��m7�����^:0x��|�+X�p!�ە��H����FCjTI�vy���:1�LP"�������<*��v�B!�R�L�����)^?������Oc, �q�v��͟��2�^�c�n��Z�x	n�󓈜p�������|F�q�o����8�u�wn-
C$BM�wahp$�Y�v�4�"�|��煡'h�Ӛ��S�b����b)F��/D ��F�A�{��7´�0v�KW�ʉ��rP� B�ɧۡ�MV�א���BHV-��g>#%�:�������o|�hll�ϳ�ڮZT��6E�&������oI�j3V����Qj,�rO�4U���O݅����̩Ӓ�;� �M�P]�\�Vzr���f��k�Dd�'��Vb�;�d�oˇ�H1�Qa疏�kz���~멧�r�y!��dc{�c:S8Iܮ��R�ۓ�[�a�:���%Q�<E�k��p���vB!�BHq��Ӈ�+@c�,�;��1��h?{�����V��BG�S��ڤiZU���:4�O���V�ٝ�|bѢEX�j�aߑC4o#EG���p�����˪Q�����^���d�ڞT;Tc�9�����n��7G�A�
������*�9(�$��~�b�A�4�A�/6䠺c��t�tD�2�:�|KV9���M$����
$����c|���QVVf۵]��]�M��p쿤�6E�N�����ܛl@:y�X�vZ����ON����zά���#���� <���>��M��u��cz�t���a��#:Ǉ3�Xqm7� K"rf�C}[>�G
�=[w`xh$�� /����c��̼L>�{{��<!.h����)�d���B(�<Ġ)E���?LRB!�B��+�!L�/��.�˥������_2�jjj��i�i"�XÞ�E�_���G:����D!1q���*i����h�8�ͻ���b�Jw�<�>��O���ow�������{�D�PF�h��aXs/��j�����z�B�.�����?ͺa>B�{s�/�����`�5�����!��SJ'M���&:�������7�x�t����~��t�w�׿��x��O&/4-�Ά�n��4�u[hh("�)J5���.�V�m��-�+���%iz�p�M���;48$��@H6�E�֭���p��N�=cm�7����c�"�/�k�<bS�o���z)T�:��� ���k�Ib�̈́����:��x�ڹ]/I��*���!ɪ��rl:�$!�B!��8�W��{�<0�.�F���`h�+c������?����m��s�Ayy9)6�;;�I��7�p=�**q�B'���9�(q�x�f�̚3#�c8t�(�'�AH�2>6�[�J�'$�Zqݟ�v����2�A�0�+��>y4h�+�,d79譈�" �P�^�Oգ>�-]�V~�4i�x�Jvb�L>�r�A��EONViV�dU����J
 Ye�3�=�6mڄ��Q��g��&,Z���~{t�a�N�VbÆ�����Z�����.C��~�ɭ�/�&����NMM����uY��r�ףzZ5�FF��>��L7t��^��ƙ��%Q�����2kǻ�Xk"rz�{1X1]�!l?q�(�wx饗��M�M�{&����b����KR���A'��.'�􅘺\\}!�B!��������+c,@NI%jl�f��q�F�w�}4��#�Ò���{>%��	)F��ư�i�����7�r�UT���'��؝d��.]�s�χ��ͭ�q���;�Cwo�D��<�裒9����ro�ͱ���o�����C�(�iͰ4��u��p����|��gWG ��Sc�3 Rz���!C1р/�qc�%%��	+�EiE��e�7Y��g�E�c�=���� ��w��-�̙��+�'-�&�4g%������m�R��wuL�jr���N����T��܅�p*����PYV.9��kj���I�~^��j�_��RN�jF�Ʉ�׹�^�"�:����t�<����h�;�2C��سmgQ~w��O}
w�q�#I�|pYH�n9A��t��5I�ԉ�p�~U�k�UVU�g�~A�[!�B!���zMcISd>����
7�>�@����r�E;x�6n !�N�+�$�7g.��.�����y'���؝XF�/[����I�X�ζb��= �$8��	=�.�x���z<��3�y^�f=�@�cEEs�C͈ϲ)VP6�ү4�vy�ى�VL��'�C�P:�
i�$j�k���C����pc�I�>��/)Y�JX��(�udP�.�UNF�ɪ?��O�x�"H�#~�?����7�BccC|�%���tm7۬\�������ܺ�X�����
�m�A����Ϝ��WVV��O��Or2���!2��m�5kP[W�`�s�l�؛gW�n�rʵ=�eC�  ��IDATl"�hvV\�m��<��I�����9c疭�����<��+��M()�U"�M�v��
a��>2]�Jf0jPzm��ALU��w��uB!�B��=<<����$S,=c,�h��1���W�sh����vyޒ%K��O��?�!�7h>z\�s/]���(]�.J�@��o��NT�����?v\:��8.[���,FYE9ZεQ�N�mgZ�z��wx��g1o�<�_e۽]y�'n�d��%c�`B�nb��f�������3������C����>�H6�Tn�"wݡ#�/�$��am�V��*A]]^|�E|�{���9�?����k�c�tm׏�Q�F��3��)�76k{�Y�Zm��a�R��Ǎ����S�k��0k&���g$q�`� �;&Ő�@\#,\��W�@�*������V��m����\�Qlѻ�[�͇�H1"����;���x�'�|�V�ʻ�T&�ɖ{{b�:Yeֹ]5Ġ҅!�A1%����"��FB!�B�a81V9%�jc�tu�lc�j���C����\��ψ��=���������ދ��1Ca�E���/^�w~�S@(���}ӦM���(HqSSS������u�>�9׊-���b̕���Ň?�Ċ+��SOeT�K��u�Qc,����P[;L��:�X��1c,��Z����%�-@�
܋��ȕ`�z>BWΩ�L#t���nꄕ։AvqW���ɪ\~�G�������&o��ى_��Wx�+_V��s)X�"t�G�]�����iQ��uc͋E-�+K\��b8���A��	ާ���{�/�������L��ۋV�Z���֢��.r���.@{�<yL�wξ`��1�k��Xܛ�u�o���H�p��atu\ �s�Ε\����5�v(��:�v�ACq{.*�{䚤n�|�k���B!�R�l>�e�c�k�4�Jz-���o��oA��8>���<� **+A����i\�-���k�P�󣵵g#S1��q�[�h.^���
L�p�T3���3���a�G[9���>W*������;��.�굆X�{D�ڡa-Pa�7�
�`V�.^WT�c�y���
܋�-�{��k}��bP3̠R �n��$$Mʄ�ϧqbP$������gD���^�VBtA���� r���;��[�����m����ܦ(|W��&�oI��qk�@�4	J��X�b��n�����/_�bD�+WbF����bht��OCkg�&:���E���?�u�iIpo2�h[0�dl��G�����8q���I��ӧ;�(��N;�ɚ{�2)�K��6NVYua�'�8:X�0B!�B����mQ�n��c�4bw��'̱lc����5G��z��v��	�FGF$�����#���LNN�����kq�,�7��q*��11>��ǎa`���BA���\�e���O��`?�> ][B�#��w}�U��p�w���]�˧z��y	�XZ#,����X�L��)��Xf���~���H�C�{�02F�����@ii��`��L�������3�E�Ps`)��%IN�a�d�ӟ1Z~�u��/��/�_�
�;��CcC#�\{M�B��D���y���T¾��q{NE�ľ9�m�n�z^ @[������r���jl�č��sg���҂��)���q�L,_�\ri���111��p�+*f���)TTVi>�}���:��z}���Z�����C/و-D�z��i�.o�O|>���u7�ү'����{����A�.r�J���k����B!�B����YS�?��K��X�:���$��{���2�L>c�������̋{����8�w?���FB�#��:�IP[S���\��i�G�J�X��� �`ƌX�b���H紡��<s
m�1� �����	�w�Aow�w#U����5�\��ݪ+&���Xr��ԵC���|ߙ��M���c��p@��-�cK;���C������t��M9�pc�]܃A��#����� '�r���g�NV�Y�׾�5lٲ��� ��?�9���k�7^t��E�n���: l7h@6D��m���m
X�ؤ^7���b_��p�#!x畹����U�#G�_S��u�--�����K�`��E��������L�'X�=��Ll�]�5�F�k��u*�ccر�#���1�}�po��XIy!���v�$U($�0Ӻ0�I��f^���H( �B!���D�b��]�˰f��a)̱����V(�˥vqW�3"z�Hc�������_�"�����;�4�Bm}V^}!�14<��C��kkj�d�Rlhh�F�LM�|�9�;w��y���Ι3K�.EeU�8�a`x'[[1<2BHv8y��ZZA��3�<#�`�f���:�նd�X��XH�������+��~����aY�bwӽ�P�^Dt�Q5o>ƮtYrP\�����J=�bP9��t/��;�3�5k�{�9������4eee�6m�B�%��ɢ��,>���w�ug䦭Jg��{^�x	�� �F��H�~�/]���oɒx1��]]FEe%�	Xu�f�M���˗q��XŬ�5��vll�CCL�-�w-��ݗ��|�8�n��� �`��=�h>~2�J�D�'q\�~Z�8���A��zD�]�s������0��!��Abߋv��@����n19��n_�����1}�tL��������t3���v��.��1��T���+ǻ�d�F�.r�oE�n�M��K��S��>�om3�����,�@���Orw*-+��Nd�os���������GǤb�@|���?�-n�O�8)��������[�xN\cY���K�#�<�6�Ny[�VL0�ޮ~V	ۣ��p!��
���$UM�t���vB!�BQ��˟�1V�>-�1VT�l��́1�a{�c}��4�����CuM5�-\ B�}���p�d�V(t�.��w}Rʣ�ĥ��R-lpp�Y���1�|̚3%����.vb߱C��i!� j���s���W���<7D�N_��gǽ]Y7L)L�%ʦXAS�v���B;���i	�^��"cwO�Er��/'�R��eG��|����&��uqϕ�SɬG}���=
'���q�����+���9���.M{����Gy�Z`$������5W���wm7�֡�!�Z��T�i�]�N��c�����I+�9�6��
���V�]���4�DOw7��\��Z�V:���(��X�����]m�R�F�G"�_[�����1P?��lX���Zi��l ��K�q��qId..n ���&�����ݾ���*��+�G������}�s�Wr��Z��~����xי'��kkPSW����$��X�Yc����H��`�KǠz��T@����`����+�3}�F@�̊���M����F8�Ϟ?ב�&c��nth�sg�&��1k���>�{��Bߕ���/�;���DaA\c��8����ˆH�h&I�n�ׄ�2V������\�ɨPP9Ԡ~�*>_����` 13�X!�B!DI�H��K�Rc	w�ce�|�����/������4�8�-�wy%��v�m1i�s�p�� �PQY�6Vĵ�n���Y������S&9n}w��?�c����������TK�!��E�cU��,zr�ꄢ�%ȔN�b�h!�w˨e` r̷���m�ω�o&�/j�������_�W���n�ik�h�`�
C�Ҷ��Ν��߽y@4	3@7(��V<�������~w���3��[�}�%�n����[�Ш8Q�sω=7��z�B��]i���KU/L̯l��+g(n�
��AܺbF�.K���T�ܣb�`d�:2(;���KVes�����ꫯJ��'y�o����������+�����'��O@���N�f���"rk�o�?:<X�8+�L��+�{EE%*++��f�j^�S4��k�v���(�&3��+ȸMz����{yE�鄁�}�m��ݕ��'r�����G��6��:=rðj��(���W�Z����@�#�@� zzz�iddN!@e�_r�����pK��{����>�E���A��1�\���]����>k�D����uY;��ņ��w�l_�=:�a��5۷� ���K�.-�l�,e\t�v��dD��lr8��vA ��t�	�cI��>�w?:�;l���k,�z߭�y})�ͳg�v5�de�v>cڽ=6���$��*Ɂ!:iE��$��������vWL!�B!z����1V V7LU?�c	a{�����(F�{��wq��������<y*���+��/r��K)��-�N��>��&'DoKW������^�u�m�������{�H�Nolpe�Ű�+*���5�7{�T/��9v��%��E��!n_�t)�@�ubT��.SUU%�g͞���ӥ���y2�y�"�"�R_YU���d���f~B0�c��ݏK�p���qe�mE�ߊ�]���l��w�b���d�)�Z��k,�n�n}�[n���w����|5�J���ͱd���$Kq���$+j���1Ɗ�����`�>X�8X;�
�!G�����!���?���p�Q��r�HJ��r`�M7݄�~���oA���#G���������z�E���X'�Vb�������� *5n�Ia�c�{�";�s�վ�7u�Ŀ}���|�t�;�Pŉ���͑\�++*�s��	G��ztt��C����G� ��B�E�_r���	Q��|�+���ҿ�����$�q�t3��i6x�������]e�x7����oؤ��n���y�jl��z�N�8	�=6l؀/|��8+�[�[�:Ie��Ҿ�s`�wb��C��z�Ae�J*T�-A0L�vB!�B���@7/�����1V��$9���1�$nE33�ʤ�X5�z�W�)�l�,�##���|�{]sR̈z^��sҤdxh K�.�5�VH�A	)�	����w�=�������n!j�bD1�W���ɓ��7�O�c����Ckg��������f[�v���}�פ��e�ŝ��:���/IȮ���'O�eqa{L�n��5{�BL������{+/���"�dw �.�����dG�ȁ,:Y1iQG�����&�|YMV	��^�Un��|7q�۹s'._��->ڴӧ��M��lQ�h2�����+J�C�����[��Tp�Dl�ž�D��/�b��e�J)�5��
3������ʊJ���J�!�B�'}V��"���yrrb�X��A�?��>��3:6*=�,����P^8��ϕ��I���p]�c%�)v���X&M������@/�.v(D���a|b"i߄��kD���Έ������;�~��|<�3]�8��	�{������R��g3I���Ʉ��%����u�$����=��r���$F��t�I*B!�BIő�,	^�7�ҩJSd�/�c�����X�e�&�oN����!�7Z~�7JN����A�E_��ݱ��y!��0�j��@o_�2���^?���쪕(�N)�F�����X�(FF�1<4�9*�ΝB� ����	VuM�+�dX�_q�E�+D��}�҃��˸�y�4!$�׃��n�@_?��xꩧ�v�ڜ��-�n=0�g�?�V$�+m�Pg�gف]6Ē��)D��I1�`u�%<z	
܋�։�莊�S82h��"	��dU\�HV�fC)�2���7�l�s�̙x饗�_������_Gn&k��ڵ����I���R�l>֒`��\G���`s�Y���W9�g�:6Wb_��2g���H=*T�S�Z;�E��P�1S���`�[k��m�d����k�q�̮Լ��j�N
���H1#�\��n�����x��'�~�zǓT�*t�&���q�*[����uA3Ġ��_��K�w!�B!$�k��F�$cɓ�'��V����"�U=(�������،�v�؁�/�x����8R} �n����F��z��JS*D-D��b��Ƃ�3���e�ҹQ�ʅ)���d�%�#1���wq�'����K|UU��'&Y�xr*�y����Fϗ�u�q��(zGq��Kzo�w%��?��CW��x�b<��s�y�VC���V�ە�X!�)�~�Pֹ*G|���5���V�۽�E���)<��cÃI����{�{�Mwe��D�yA��Rw����7�)^7�͛7c��� ��?�9^��KX�d��ޒX7G�vg������x\+���%v�&"�����V�j���k��U������w�&X7[د9�ۋ�W�v[��l�uC��<R�g1L�f�x��z���U�vNp­��gI'a�����J��Jvo73̠<�`ii��� E�N!�B!$F�T=�Q��9V:S�`��/sw�c\�1Ɗ.J��9e���.�3f���/��������h>v�Ӫ�j�� �x�Oˮ�@���^�ԅ���B�8q�(Z�O�xq���o|uuu�����=.`���R�ci����J����X��@�ܣ��)��i�������i4�1p���INFn�v]�u�U@R�J�ٕx>��r��_�u�߿ccc �B�����_ŬY��L�Js)V6�S��6g=ָ�&��C��
X͋}aK�k�]�q��H�wq@�������e�x�V~W�`Wnk�7�k{rX~�G����	l۴�c� �C\����zWD����J$���̹��vaH��-���3�k\����@!�B!f�{Ac5`lx(!P�b)���^�1��ϸe����cӦMضm��8�t UUӰp�bB!�hi?ۆc�x�x w�}���Vn�e���bv�~/3�v�1��k��KY3���f����{
܋��<�d����+�U�F< �۳�������U������իW��_�2����{����G���x��WQ[[�i��͑�=lO�l_�k뀸=�"r���V�����>����M��h����T�:�ry���3��W�v��k;���?�ÃC ����ý�ޛ�$��I,{�ǧ�=�F��MN�IV��T:�Z��f�A���� �B!�b�󁙘���͚bY1�*)�E�U�Cc�_.��p��X��� �B��lہ��
̞;�B!2��.b��] �D�����+����!�S��S,e��h��t��F5De�P�ό� �۽	�E���*�5���]$O����:�g��R���v��L���~�����q��i���ׇ�|��x��PQQ����\ۓ�s)V6��-"7������������žV�e.ΚX8sa��X�������a��ߕ��6����V~�6����aa���k���#���Jw�7����kI�܈�3qoONRe$l��Q�$U
a�ֽ=���oX��n��B!�B��H.�Qc,�!V@�⮬�5�*)��W
�i�em�ʕ+���O�����A�����ܲ��̽��>�B!}����6�:�x��^z	�-r�F�d1�g�k�Ɏ����F~N�O�ޞ�n(���x���v�B�{��LVŇ����]ϑ�L�J�R%�����&��I����
N��h���Ւ#�[o�%�{�=:;.�g?�1�~���;#l��،u@��h��ľ��Y���m��0ڼ��l�V���	������^lA��[i�����ۍٷs:�;@��8����X�x1���J�<���0�k�U�Ĕ�}P��
��������~l�aF!�B!�lD}�+�)�9�d�{t~v��
]خ\�����1�ɓ'A����$�o��~�~TVU�B!����0�m�,]o�a�<��cyU#tG螬�1W+�^KN��XA���ں���L6���ޅw�JV�\܅�ƍ���=�^���&�R$�"�O��dUt�ۉ''�if�m�݆�~������MZϴ��?�',[���\۝���X-lߴ�7��{{�v��ۮ�F����&���kr�s"r'��v�wk��Q6��Vb�濫�!r�_�gl1rd��E��wY�v-���/�U*�I�D
�Iߍ��{�*e0Ġi�����fD!�B!���#�G���Ȑ�+��{�ߘ)V�+��9Z7L���XJ�,�C�	����䋉U&�4����*����9�>����>������B!�����}�c�c ޤ��o��&�������۔8m\�Y���a8�di�g�1V(�� ��
�I,Y5�#��.��d*Y�%����LV9��ufs�x-�U�w�Fww7�79y�8�&&q�'oW] �V�l>֎(�86�bes��D��������m��:m����(6����m�B��F�����Z��-�.,	��g��[���z!	N>��c'@��HN���ۨ����s:I�ny���$�R�0�JR�b�ȅA<����/�Z�	!�B!$S.c�ܗ�5�`�y���9Vd��+1�s�1��}�b~��4�~趉�NlS+��y���7��&��ضi�._B!�±}�bhpĻ<�����,�����ν=q��5���5ŊNA�Xto/\(p'�3Q��MV�M%�"��KViUJQ�V�+pqRˌ��9ud�d��ٳ��o���.�w�|�������?�c���X���D�v�f�i��L�+��ޮ�c�~W����uLD��_s��n�3�tm��`�����4�Ʊ��A�ͳ�>�����4I�F+�:�T�\�U&.V�TF.��K0�Mq;!�B!��a�cc,��{�f�_���{��`d�'��5C;�X����5�c��{����ě\��EYi��Z9^� �BH�#��?��W�@��ҥK��/���F�fQ��W�g�eT;jꅉ���a-��
܉D��*����bSP�̴�*�2Q�x��,�>�Kɪt��A�ne�C=��۷�����.���@MM-��.S�/:#`ͥX�^�~[-�+�����V�����LG~+�`�X������n��vm����$X7g�].?�b%��vs��m��=M �檫��W��U�$��I�l���[���J�����	�S	ܭ$��\��~|�B!�B!Y�+<��X��XA��(F{���BP��McA�WU椊�kƌ��7��w�yĻ���`���q�]wH�!�B
q���m�|Ļ�7��M��չ^t���&��R��bI�B�u0>�s|h���3"�
�x
�Ie����]�*7!|ɪHg�����i:��{�D�^�J���U���Ӊ#���t������Ž��	��� ����ǴiU���cr)^tB�k�]��{��&l6�}�ޜ
���/J5�]mÍb�z¬�݁�꜈܊�^g�#�{`WD�����4-�7�<]ۉ�K�]ػ}����;o��v�m���&��-7^g"A�c"A���R��HRI��{Ҁ�{�H7�7B!�B�;ڧLc��
c���Q����'p�d����K���{�̱���?�x����۱7�~K�\!�B����۳m.^��6�>�(�㎼��Z螸oӘc)�!��hv�g��=�R
��5�3��y��
�Im�J���6Q%'��	�H����d����OV%92@-p����J2���ϟ�W_}����@�Ϳ��_QVV��6nHZ朰9sq�mn�v�[�q��[��Tp�Dl.žf�d�N��ڦ8��wuFDn�����|Ws�����r�8ЏP�m��]�c���u.�6O?�4n��Fx)	��$�n�*�dօANRE]�e���I��PZ�Öv��!�B!�;t�g�.�1��n�o�ҭz��n�1�ۗ����ۇ�/�x�s�gQQY��7n!�B
������<��Y�p!^z�%ռ��«�_�O�ꆖj�s���=1i�i��ۂ��{{a@�;Q������:�{�2Y�OVE�4��Һ1@�Z�O�OV�M,�˂��Gy[�nŖ-[@�Ϳ��/Q�+���I�s)lvB�k�]Fq�Xu��ir_Ym���vY��|�iC�����pm�ݼM���X��p��|�� �"r�ǻ�8� G�Wa��}���:��;��=ر�c�:�x�U�V�^P�s:�dkv�sI��bBJ9A�LV��T3��UtJ���qo��%�B!��Mv�O�E��a��{�W3�����;i��+�l�o���x�����~�9<�s��I�����ցB!���}�z�������ַ��А�5�t˳UCL���̛b����X�b��a����D��� ����Ã�d�*Qe 4�&�CJ����U�ӑ�L��� �K$'�F�*%�$\7��L����W�C���������%%��\���gl����R�l/V�����\>�`�fŵ]3ۑ�J4X�Uf��ι�g.87�Wf�oi[0 ��y'\ۭ�Zܛ�3ږ�8������I���1jڏ�o���x�W\o����4I�+g{I��ܓE�	�3�*���b*+�cS;!�B!�8���#��qwq_��c�
����h�Pi�U��7�
��c�Q��*� \�E}�h��>(c��O�6����k�_B!�x����Ա �G���y�y[#�E�j�PO�.&=S��#{�����t�b:;E��B�w�ĩ��\��ڵBw=�A���/����dUII����ua���P	ܕI��]۩�p=��F��-�׿�u�����@������?Ǔ�|�פ����t��D���;�M�5�"rb_�X��]q=���?�"�,�9���J��n�9q���ݠ�s�A��{�M9"Bw*� �W��~�SSS �����-����$��$���'N*�ۍ�T"9��T	*Iܮ^0_@�aF��N!�B!��4�R9�+G�N���A?|¡=�F~����X%P>�4�����(���Wu1a{���HUK|��7%c�K�.�x�cK�?_}�ZB!Ļt_��s�gA�ς��+��լ��ܮګ!����(5���Za{jS,1�s(a�%Mi�Iu� �f������$up�����R%�dwI�KT��jGw���&��bw��aMG*w��y�L,��f��_���Ȱm�6o#��_���x�٧q�իuc�
s&��Ю�X�f��ka_e��ᤰ\�R�׬���j��:m��m
֭��M���C#������k{�D���\�S�n���~|��QV�۫B`ٲex饗T�
=I��<!\�bJ/nO���VJ9I%����k�������gB!�B��D��zMc�uÄ9��K9�s�K[/�k��$���6ƚ7o�d�����f~� n���Zk~�gB!����N���e�#��_�u̚5��̰�����L�Rdc��4#>��
c�c#3"��!]!A���`�/G��D�2Y%��+�Vqa{ܑAt8%�$UB�LV�"�'�d�{�d�]a����pQ��\�Z�-�y��8q��� �F��ӟ�+�=��+V����;&`�)��6�u������V��K��������oC��9�v�+p"���*�ǻ����o���$C����������� ������QWWWTI*�r�	*��[rp���bw�[{��������1YN!�B!�9�1֪es06xEe���i��^����!���	��XJS,�1��^�c�|�+���L�6m��}�; _��Zy�U �B�w8}�$�D����� �������_�fX֖�SlN�{:S�ĨωZa(6iGz6����6���V��*0�.�zX�b.F��S:2(��j7B�`<i%:�D�x-��:2��hE1R���9%����ƺ�b.\��^{����(J+ ĉ�g?�q\�n[D�+��v9&`5�}K^'�������)��+�ς�ּX�¶��n@��k8���`�ǻ�:���-���m����h�ُ�5Df����� ��3�<�[n��I*��4WG�n�y!�����`�A�}մj|p��vB!�B����,p9�K3��n菊��џ�I%nO�9I�Y�V�n��i�,�j������-;v/^�>�4I�,[��B�Μhơ�� �����曖�J���Ś]nv��{0�Y��!idg���Jc,i��K%rW�cB���5��@

܉!�z����r�SP:2�ĕ,f�
��Mv0�uc�%%���:�*ّA+p�]4�*iN�U��`%q��#����	��A��,r�`�U�����-�mp-ę+��t�Y�w�x�岀�8.�b_+�2km_; ���k��v9�]ͭ���n�̩k��88�������ׇ�� ���5k�}M5/���F��Zn���6Ġ�켠�'�0��I�v����{������@!�B!�@�K;��v�g�1���}��?� ˧�WL���W/E&�|��!
���Fbw�c�
����*�r�عs�⭷�¿�w��0طs�t\�XM'wB!$�ii>��{���G<<:s�̼���V���Q�c���P
���c��1�^�P;�s�h9Cq{!B�;1��?��W��ؕ.]G�N$���qd��yr�*1�`A+t7���Q�N5_���l���7��<x��� �G�|����K_yk��F7�PD�+�ѧD����E���C�{���W�u��p�v��3�[�+V6�x.E��(�7g�K�s�u���n��X'z1ؼ�u5}�W���͘���`����_��_cڴi�'����̓X�$�4�t�Jx�T.�@za�2IUS[���'at?H!�B!$�$cE�ϔ�C��=n��u����c��d�1��պ��>�ܹ���oA
����cb՚�A!������q��px�'p�]w���Jl��'��4�X�eP����c�ҍ��c�%�p8���@��w��m+pCyX��
7m'"'���x�*�Ŝ�J�z�DבA%r�Z�''��dU>&���,X��={6���oKO���G���;��g���O>���U-���R�k!Ζ��b�Y�w�x�eUpos��ͥ��l�>n{_g_�O�v��լ�����>�um��_e�d,Q��݃m�6cj��х��/��k���I*�$���~�Am�*�HN�sa�'��΅fE��c�B!�Br��+3Ē'�{:�n(��*S,�B�����tE�P������r~!���Ki�u��9�������I��ukA!�������c���R�PI.�~n���k녲9��ڡ�^�1�
&j�1c��|�)&z�&y~��E�<Mq{�B�;Iɥ� *V-�xO{\Ԯus׊ەw��Ȑpc�&��Wrr*���:����qd��i�l:6�����;��c�ᗿ�%Ha ���L}�Ql�x�����be�dEDn���^�������|��}mM�6g�ޜ>4����޶ۇе�|�ۂu
���s�2�o�SS�7�t�|�ɬ$����R#'����ҭ]��JNV�D�DSHG؞�ĠMRń�u�x�,�AB!�Bq�1V��K�n��
��_g�gq��5�J�F�!�S}��^W]C�Wa���Ϙ1���|�M��A
�c!9��n!��>��&R8���I����Ei��~��f�6�
��^����>�cik�w��β��� �	�$-�;JqG�/1�b�Ay�A����/��Tn�!�*��]ב�DUX���I��7�M��qdx�Wp���>}�p��_���w"w%9�Z�sB�nMDn �5)nwFp���v�ľf�d�q�b�����n����k>`�_0����k;1I�������X,$�O���|�;(//�]^Lnj�:Ae͉!�vl�b0*r���%��)�o���wB!�Bq#c,��]�n�0�
J#?�����F�P��k��O˳{뭷⩧��O~���A���q�n�B!�=ăg'�),��ylܸ�hͰ�u�dQ{�z�~�P�gu��ص]�*k���a e���}���B�w���� J,B���:I��jWԍAv0(�3�UQg����]�l��G֯MT�'�	�BsY�[__�o}�[x�7�.Z`��������ƛo��;#`ͥX�\�Q�Y���j=/`5�]��S$���Zi�~��6~���bs�Ј�{{�tm7�`��v�tu\����I׺���u/[�,��'+�NmK;�t�
�e��^�*�����$�ERJ���k�K�vB!�Bq�$c,�)�_�K��Q�ea���]k�%���
c,m�P�0(c�+��n��Ċ�/���d�u��Q�¡��q��s���@!���spOΜ<RXlذ�>�����/��-+��"we�PY/L�9$��
��k���:bd~ii)6��"�
�.�S|p��5T�9�+n�:2$����z��%�����h+w����\����zo��&��_�%�������o�ѱ1|�t�: ��爀�R,xs&�7�|���Ή}Ͷ������y��.m͆�=��u��+�����ݬ����Vb��o�>�϶�i�.隔��?>�����a!�I�t�R��k�JP�qbH��S1��ƠLRE&��4PiGQ �B!�7Ic�%��1�{@��T7�w�)�v�gu�Pk����'r`�#@;e���u9e�%�����o�����)N=���Il��ƴ�"B!�dq��o���i),jkk�Q����t�Z�0�1�y��u�䑟�\�U��ͱ�
a�4?0�����f�С���bl*��i�Q��j8�V�.�W��ew�h�Jv0��'%��ve�
��]�ɪ\
���v2�������СCػw/Ha��O`|l�>p�o-�D�+�ͥXY'>+"r��\��Nۣ�z�vžV�e>�����~�Nã��'���9�v�v�}��v��S�n�ph�>��dѢEҨG�>E�n�\�q�Jߵ=�HR�9190(RF�ve�JρA̯��g�P�N!�B!�����x�1a��4Ŋ����XZS,�޸n�4�sd����+��v������/����RX�4����>q�-�<!�B���.ݳu:Ν)<^�u�^�:oͰ��fo[	х�V����k��uG}����+놱��beU~�RP�NL�Q[��c�#�"w�$����/;�xMR9h(r��EJ^A+�R�28�Ȑ/ɨtɳ��r������y����;�n���y��O���-��gE�j�bs�4l�M��6��V�����8�؜>aAp����ᰅ��S���u��������o��\�aA\O�������.a֬Y'��rc�e��ȁ�8A��� '�B�2��/�HT���-��!	!�B!$? CUQ��b�+�+����퉺a��ݠf�CΡ�1��"y�mx��gq��alݺ��h?ۆ��n����#�BH�ײ;�lť�.��C���裏:V4�L���rum��K�~�5��3ƒ��Q��ͱ�������%�
������&�Z�0+0 i�4Ԡ$lW$��L�����rP��Ҿ�R1���{ul�����B��n��Δ����WU�������S�o���\پ�nuuuV�u�L~���5׮M�ʐ��t^�DӮݖ4�ר]`��+���뽒r�[��Z�|t��ȍƁ�}iV`e�fE�����FG1<4�.f�"l�t�PX����a�m����i�im���4:2*��=�=o����	���<r��:��M4�Jd��GO�ޘ����H��^�S�2+}~�n�/E�r�Tl��N�Z��u���`�+�b����z��0>:�����vڝa��M���D������]����9��k�l^gX��k,+�^to�����э�n�J߭�ع]��ҋܵ����%�롸�B!�B������z�������Jc��џCIuô�Xr]L!vO��X�XW����"g����hmmEW�Z�%�=�@n�[ۗn��gc�Bl��͸���#ksy��t��S汝��m��}ї��}�������&���}����u���nQ��;����oK���?55��[������y��k,e���k,+�~�x���9k�z����5C$��qm7�9�9V0f���W�����Sp�Br���������MRi�Ը2�_!|(jP)r7rP�����EC4f�+C��*+�n�,XIb=��طo��_�E����/���}Y�499�����>��]�����?��+*5K�_B�~��7�^�i'n�߲r�'�`�B]�ё����x��v���7���k��� z{z�l���Z`��TN�G������P��l���S�V��}���`�X�OXqm�zq��3on��n�l�Ѿ:q�(��vmR��m�h[��B�~��5�Ӟ��ŎNT�֠���DK��6���i��/�z����+þajr
]X�|���M[��]��9g������/]�m���J̞?� ��};v�|۹����5V��3� ���<��5���w���%���S��1�KR�3�q_HNVA����MV�0TTV��y(�B!�BH��%8=5������]���9��9�P��n(f)k~��X���&��9���K���s�J��~��q�����UUUp�Wrk�⻋I�?r��l}����ܼ˯Ziz
�{�q뻋<nW���P��k��藄I����]��pd��cc��OF�\��B�.�P�P���y���Hn��&&091��b>���vdx�"FI9{����-��ݾ�rs�b����)�73�7���=˿���3g�̉x=_j�Fˣ�Sl�A�P[7T��
�{0.n���H�4�slY����v��^,P�N,��W����h�#r�&��	�`l����];�`ԕAߍA�����G;^�s��s�@�溲!���|�M477��ѣ ��pr��?� O=�4jjd!�� �쵣ia{4�\���2k��7)̵)`�&��<.ulvž��F��]������n,�"�p�^���� ��+�;�Ě�m�A���m�9�sK�7Ļ?ކ��N�¤����***t��C���Z�`$hW��]�b�����T���0IE!�B!�ȡ�SX�|Ƅ1���]�k���~1O������亡Rخ�
i�Os/%yh#c,%�P��.�m�뮻��#��?���3n�&���_YY���)���NcMNM��ލiiFz���h�.\ 7���K�-��~�i���]�~1��˝QSW�i5��w�L�/a�Ⅾl_ț�.��;257���Z<P4k�W�`�q;<4���lK _��X�K�󸅙���+�ছn�k�s5B��DM��+]�PL����>k����55CQG�m���-��˜���U1�ۙHRiD�r�J��roW���C&;2$�1�ܣ�&�2h�UN%��-�E���jjj��|/��2FG�y�8���.|���{<��3�5{V�r�BIkbes��D�������Vž%ڇt���V���m2��"xgD��*��kǵ�(�����dlV���~�@a�;ǖ�~���+ ���&��e˖e%�TxI*��	q{����=�Z��J����B!��Q�^��5%=�{=IخqqOvr�Gk�:"�Ľ��nhd�%>�}X[�g�%)o�sQ�溲e�%�<'O�DSSH�!�r?��p�=wazC!�b�+=�R�pb|�0���[�r�g+��Z�\/���OV��ʚ���];�sP��rr�N��zv�L��͝�S�;P�N2bsG��E�Qr�J�ZύA9�V�.'���jG=7��]�.|Њ�ԮF�^wY����k���^�����0������ɧ���K�H�r+V�k�V�bߜ
�3�K��7�6.u���������pm7/X7�!��|g�0�������i������N2B�/l�`��/)\�x�	�{�YO6���l���H��3IR�LP����TCtU�` '�9� !�B!��;����a��˧c��4��5Ŋ������Fu�0QKT����ʆY����+z�\��X���*|��ߖ�����A
a���p˝w`�� �B�y�:.`���%CR��Q��~���9�fX�c��v(���^�P�KYC��S�c鹷����q���b�w�}c�Nh�B���K$��!	+��]��Ҋܕ�Ɏ�"w��+������1q����&����СCؾ};Ha21>�������_�UW�6�9���,��͋E-�}=/`5/Vv��<�Bd��F�Έȭ	�Э�߆�ݡ�Ftc-	��f�os�o���=z�{�c�G���.�AO�LfՁ�knV�T�T"A�.I�/xOva���Ӹ.���uU���p�CB!�B�'�X�����u:"wm�P�'L�*��N�rmP9����]4FQ7L�?�Xn	۵�W�Z�7�x����@
��T ;6��o���ZB!����L+���#]k��D�S��=���Vb�yz�v�	�z���=Q3L����Z0�Ҋ���~ljRg���$c�|.��ά�7�qq�KX%�%��q��,nOvd�{-�,����NTIsJ�;2�C���甯���s����R����?�'����q����/V�k��6)��"�Չ7ܺbSU����}�����.&�Ypm7�k"�|�� ��+�����Z����ݢ������B�SWW�����AmmmVSVב�X+m��3����+�Uz��PH� O!}Q{�vщnﮎ���B!�B��d��`½g�5Ø)����]��=^/L���X%I�v�~5��a>ce;�����/H�X�6m)L��o�n�����ցB!�?tD�Ha#�a�ﾜ��|.����Ê)6GY+Lc���#&�#?�������u�)�f,��e�ۋ
�I�L����?�HRe��.%���VF"w�9�SB�r��$�WFu�%���Ƞ]�f�w��믿���1��������Q�uϧ�cS�}���Xk"rb�|�ڊ͡��t���Z��I�$V6k,�\pn��r&��k�w��������e�:�7P��.gN6����ܷ���׽�W��zb*�r��JvbP:�+]B��v#���{{E�"t����B!�B�ğφ�9�059���c)E����h�P�9�1�@�.������9�����&���p��a��E��FGF��OH�!�B�k���p�������ǫ��j��M-�Ͱ���A�9V���ܕ5�T��t�XA��]���V�k���X����b˹ ����Ã��+V%�����=��23�`8��F_G;�h�N^e#�n���(3�'l1����������6t_����(*�˥yFb>G��a��w3�̱��^���J�v��	��	�ai[�b-}W�������[�׹��3��G��C{����S �ϓO>��~��y��2�l�!�I*�����Cl*++æv?8� !�B!�x��`���P5r���ݴ1VL�.�eq�c�D�Mm����Lb�~�h{b���|�;x�W088R���i���(n��(+/!�B"װSS���v\��	R�̜9S����:�uA��p+V;O]3��6�֥]׹=ͨ�qQ�A�P�=K��X��������^�t*�����\��{ّ!��J$�tE�vHI*��=�z�A�d��$�2��x-�\9}�4~�߀6�O6�'��<���t�[+���&"� ������w�/�5�&�u���Ní������[����r�x���,<a�m����{����w���� R�lܸ���ZV���в�^��&���ۃ
q�����
�������1t9B!�B!����|i�L�����6���}�Q��N�F"�T�X��f9�m�+۱�4�J��5k���������2/Y�\�Ѕ-����.�}~B!����0v|��|ȯ��b��e˖e���K3,+����R-��#��L�5ĠB�n\?L��{]�8�R�^�P�Nls�7��V.�ؕ.��=#w)a��ۃ
'�dq�*a%�MZ�eRՉ�آ8��`�Y��累�z�-���p��"�bg��������U��X-��M��mǰ]y+`5�]�tmOw��5�Z�}mW�l.�9y>
�a���U��w�߅��p�\ۣ��
�YD�>#�����G� )|�����i�\ML�C�l%��\���r�jjJ5��n:�?'�T�Y!�B!����f`U�7zߧuq5B!x7��^�pq��C��aJ�;27��D�^�X=��?�_�� ��@_?6��'�x�- �B���������s�<����h�{���Ųe�5n��n'��۱c�]����q'�7{��&q��-�Mb'��E��"�V�3��f4]���$H |A���_?��_�8$p�������E[k+H���_�:.��Ҵ��n�ͱɞ������fuC�`,���v�>��m���u�4�g34�Wx�X�/͕�U�Rܵ���Ƞ�T�X��Q��-��`p�V8�PY��;c��Rm�o߾X�r��v����w��Ԅ훷b��Q�>sf‴��m�}�2�[��X��,>V6ҩ�W~LV_B����#s�C���+2�po�`�}��������{ة9��^쌥���@����U6 �=V�Z�4���	SV�K���"���=E�����,�=�\;��t��B!�Bz.�;0w���W�}ƚa��^h������#���ڡi0�keU�ĤC���lƺ��;QQQ�6��nZ�[��;�0m�t�3�BH6q��!l\�!:C�&��w�y�ַ��[���`�a����OP���bi���������G��8PFs{�C�;q�ږN������D�J#H%�&�q��,�A��h�*%�A|�
�{�w8!�!6���Q2��7}�t�X��>�(�uY��{y���ŗ_��˗şH��ܢ6��{9�M������u�Z���������mwbnw�p�}ú;�y�������/,�Mv�Fs�&t����8�M��|�������&.���#Luw=�"U���^2�R�TS{<�!Uz{�wc���!c����vB!�B��~$�S��Tc{P��97e���f��S����y�u%��4����R��ѓj����x衇p뭷����w#L}��+wx�5o!��l`���ʃd�F�>���BW����o��V��J�JR7�q���Nmb{����F�{A���k�s���B�܉k�q�7�돖3g�b��ԟ������}�V����U�
�J��"�����.#�����g�g�������Z�:N?����


���Dn� �7}�t�}���6����]1�K�:1��l6�x_0����1��ذ�����o�I�X۽A�^wlފ�;v�d˗/WZ:����nû��P����<���Š��=77o+�:NތB!�B!��ƶN4�����xr���.��Zab�0�3���@ch3�{��`,�8k�XZ��	vw=��9a�<���(�TӬ@���46b��s��SB!�7�b���ء# �A~~>V�^��cǦ% ��6����x]PolO�e�On������n�ţ�t<�ڙ�Nhp'.�� ��:�C��D����hnO�ȠMqק1$3�KD��ஊVF�JY�"��e��]c�v��;�@YY6n���ޱ�+�p�>��*˜���ߣ6̾v����nS����gSj{d�3c�7&�L4���&r�72Xg�8�R��p��:�����B剓 ��ȑ#�r�J%�A�Fw'��c�w"����Bz{G���`B'����vB!�B�M�q�7��֦F]�P<�њa���њa(��J���܍uC�`,q���3��Z��'B~��_�d�fC]=λ����B!�7!n�����P_[�=�~��X�ti���UO�_&���2b��j����ϝ��B;�v�(�? ?$�>'�!���U������#�\{���nLb��U�D��`��McP�`%�	k�*�e63m�Ay"C&�QN��2����~����ѣGA����J<��_��[nI�86��0�z`����n>6�f_��d�M�fa������Æq�o.�lX�3��k55�{pӈt�N��n��K�/���g�$�hll��-�PWG�*�())Q������0ee=#����w�z��L�
�E�N�@��Tک�QR�9 �(RB!=����Ĥ��<�~Mc3�����e!��<�� ����Pm�����Is7�ۭ���]��)�f&�ȱ$�Rki�e~�e�QK��o��ػw/�{�=�젮�o��*ιp9��B!�7P_[���>A[kH�p��_���Z��uA���f�6�*�e��l%K��cu&7�'3�wv�����1��D�����;'���(�w1�Z��)w��n�b����Λ%2�1���99�Q�Fa͚5��������4�����w��EX~��'���XG�v��v_�|�S����6���ڃ����v;c�,�_��~�aYr���s\q;�q��&t��{=x�?ژR4 ���}�=�`��i�������*.T�E�pT��=$-�*�Z�23��$���0�� �BH�c՗.�]7/�|?�'���_�B�;!��@v�`�)��RsR�wY���n���)����F(3����w�6�ҭ�QMЭP+7B������#�(ɗ�4���ڰ���0k�\L�}!���̉��Q�g���F���3g��{�E^���������_���z!j�F��ՎϑyC0���Vh���â�c����v�w�:UM!�G�C���������X7����V�J0���ј���^�R���Cvƺ����c�/V��x�	���7�F]m-���ӊpiĺQԹ)U���{/��1�¡���1�lӱYءa=#L�����3�1��X�n�ph���װNc�w�����۰g�N�|S�Fz/_�җp�7����%�)N�����T:3�{"����G��r��	!���H���o\u�r���/��N!=�7�by�x����n��9�f��uj���,��=!K\�F�A��}�Xɶ7d�<��c����ǎ�Y������4��c��%��+!�ғ��:���Í8~�(Hv1x�`<��8p���@7�v���}�5���p,�P,m0V(V?L�eZ7��H0�����c]G!*4�OX{�׎*E[KK��`�`pO��I�*c���@%��2t-�Q?��I>�����2]�rc��믿^i;��?�$�ؾy+N?�>w����g�a��!�ސ�.=V�0�ߵ3ú�q^��~_a��6���������a����F��{��=1�3�=3��{_��"�����q�m��fn�4a��zFTS{�'$�T&�,���He�����ݿ(RB!=��?a���*_��b�����yI�y	!���Z;=�>�7�Gk��g��Ě���,�][3��@��H�0��n��il�n�k3�ټH�|���z��X]�d�*�Lc#ν�|��B�	4�i�o����Z�d"�}ժU�:uj�jz^m�ͱ��`�?#�2�	�?˂�B��ϝ���p�Q?4u�Lo'zhp'����cx���C(� Ms��U�D�@@op��4���(X���+�����l���]w݅cǎa��� �E�J<��_��ǔi��w�d��4�:4�:4����q���N��f���Dnq�w���o�ll:Sϥ۴�[g�/�����mX���[j�k��;�)B�>&L���+W����u�(S�����#R��ۥ"U�4��؞�ܮ�0x"��in'�Bz��~��/�e�_�|!�]�&�+��	!���ZE׍ꋶ�f��ݐ䮭ƌ��Rj��`(ftWk���������;@�c����ow=/��b��+�@YY�}�Y�좺�4^�e�s�29�BH&s��1l\����A�q�*B�.��b��~l�;ce����aX�B����`�`��,�=e��~����Dhp'���D7M����q��!�A+V��Uc{ "TE�E�$m�{��nfrW�*%�A+Z)�*eI��D��y!@Y5ډ����x��q����� �E[k����������/�T�{X5|���z������qfc��ߵ������{a��s\޼V���x���3�xKž2lٰ��QYJII	y��92m�t��)��H��,}!��S�J�0Oo�U��E*C���~���
!R%��B!$�)꫾t����+#/�I������1c��Xfwy�� rB9�za V3��U�j0VHW'hk����X�]��ڟ��X���wp��!���� م����[�9w��H�qB!�F���޶Cy����\~�����Z�ϫ ,��pg���]b�2��)�j=��eLm��
M����a(�Ζ�]׍Lo'���N<卣�8�_^L�2�2�&24���P��Z�*��b��`k9���4.^��Ȑ�t��lo���X�f��4515���G8q�8����������J�6lX�([���jl����t�n~\��)B}�`k�dr\��n�ܞ^ý�qfc{\j��qf��	Ǧ���8
'�!R�?��n:z�0Hv"�'z�!,X��w1�+q�;�ӟj�E*�$Y�Q�2m-hG��=/D�!�!��Ƨϙ�}�*d"�=�ƃ��x�E!=���A̘2-5'�>�5DmV��.�՚a@�HLqצ��b������h�{�D���X�XK������h2ǏǮ]�@���صu��U���KQPP B!$7bmX�>N?��̝;W9O��Km��DӻW��k��p,+u�x��������X�Q<tv�gݐȡ��xJ]k'�F�EA]������VB�2U9�e�XZC bp�ъU�R�J&X�ZF�*dP"COHg�7o��^<��� ����G��/��u7߈q�G��0�z`�M��5�f_��d����:�8�d����&����{;��a>m��fc���Ә���F�t�%�i�o�＇��z��E�/\}�����NaJ?��7�T	���ʘ�.�%�H���`�͠V��Η��e�!�����1C��)N�*kϠ����>EJ���M��ꕋ�)M�ҳX{� �W��]�U�{b�{��ܣY���|(v�,ȂX?������ ���[���ӠA����"���$�8q�^���8���<t!�?9]Y��Y�֖��d�СJ������Rt�.hwɞ��!�j6��k����ΤuC+�X����	3;�94��y�`�L��z]��\���\�J4�kS܍b��`�&2h[&&2º�{J���H6�u��ȑ#x��h��R�����������/����V/��}�=��jݬ�ɩ��֎�dޤ��7b�D���o����W&���_��ƍ�2��mX�w���8��nT�I�r����[oU�T�0��-tuwV�K��� TI�)Yz��0�D�Z{8�!���C�����Ϣ�8uJ�_����?!w���|�R|��L�&wqJ���O�;!���:�P4E��	]��5D}�{0�f���F�?�dŮ����o"W	(�1f��=���t{3f�P2W�ZE�.Kiij�;��^��ӧ�B�};wc���9�N
�f�L�<��Z�W����/~��<���&wY�P̧LoOQ7�.��b�Gu��q!,��^hp'iaC�@��Ztt}@i�۵FwU��&3��4����V�2&1Ėu���I���ԽD���2�2����w�m����/��H���{�D���p���g^<41��-�S�&M���}��i�������홅�7��D���{'۴�z��n:֖���X�oz�3֫�b�����O>ڀ#�d7���H`���8�M�N��۵g[��s��`\����IA��v���"!����ɭW+	�xm�~W�����2Mfr���$w��	!����� n�4��5�:��nh4��ꆁP�~��#m�0bt7��wH�z�{dU{�XZzc-��K/�ѣG�_�$;W�?ڈ�'��slkv�BHwikkæ�*]EHvs�]waٲe[t�.hoښ`<+fj��eu�����v�h��n��>��W�Y7$ɡ����C�A̛2Շ$i�C�hpWD*!V)�Z�J��`4��S�-U�
G?�ӑ�`w=?��V���Ã>�S�NaӦM �ˑC�������3�2}��I��^�#ce#�}-���k5ݗ�C-�����5��ȭ�����o}loHm�o�}s~zozq�M�=jNWc�{�q��Hv3z�h��?��|�2C�21�kE*�8��Vf-�Ȕ*�!�
V�����!��^�.���/��r����q�Ϟw�ܮ"L��<��뗚�&w1��y�&wB�!|P�s��E�����=Z�D��ω)����ƚ��XWR7�c4�{���6�3�կ~'O���������#����9矇!Æ�B�ʓ��������݈s��}�s�������6d�ˌ�aX&uCuj��?'��Z2s{��]�%y]e�����d��N��+�kF����-1�A�v01�!bj���S�U�p�ܵ-�P�2E��z?���J{�;���^Z[Z���	�/�%�]���|O��5����k��LVwlvnX�4f�C��pg�|�u��5la���s;�צ�-���arw��c���w�:���S�g/�m�̶�%%%x��G1a������D*c{A���(X�ZS�۵"�jt���!���ŤQ��䷮L9���_�8���ٱ<��k�V{�u�&�/_�P���N!=���!̟2A5KS7��Le&w��5���H0���Y��vHk���ab0V ��"�r�&�F�/fv�*�����Ǐcݺu �KKS3�]�&f̙��sg���!����=�wb����\|�Ÿ��L�9�0����2�^A�SQñ��C����˳4+h^743�ñ&�D9�$54����
�@�H��Z�Rڵ��JIm�ܓ�UZ�J[�5���T��Ƞ[;�(7��8?f�<�����;�����l��	�9�kn���=�.����X�H�f_���V�k�fe�c�3�g����؞��ng�s������;��=���l\����@�8�衇�hѢ�	PZ�����خ~j&3���0��
f	F�J�fP*Ti��(RB!=����ˊѧ� �����%%��k��k"��^w����	!�g�jE׍.U8���ܤ�X��a �Zu��U�;�u�x�0~���nOW�΍mtw?��Y\\�tݻ�s�N��E�}�ںU�*�d�y(.)!���MM���Q]YB�̙��~��kZ2����mĉ��5�N��C�����3VC4{XMn���S��uC�IRC�;I+�Ot�)��RsR���L[�)Q�{ fpW��D�J+X�S�]"CT����	&w��Tx!n���s��G��ի�/��T���s��k��EX|�����wFSk�v�f�LNmO=z�ޘ�3�p�d�f�k�72�`����Fg�o6֋��3�c����7(�~���~;���j����2���==Zc{�ܞ*}A+X�j�Amk�Dc�Q��ۃ�!���g/���SG����o���lG���o�*��^���~��?��w@!$�	v{ۇaL�AC��\������E��0��H����ƚ���VX��9Z7�c=+k�^�E���'�?�:�Њl���)�����xٹ9f4!�'=xX�v�{�5��F���{��^��`��񚠾fh��n���vh��nflW�C� v�C(L�!��$�y���(\���L��	V�x���&�!�X%H�Ȁ�K�D�G�S�exe`�2饗��ѣ��/~B���ۯ����e����A����O�0�ה�.���X��պ��� d�2�D�ý��N_�ߩ�ˡ9ߖ�^:�:��CG{����@����_��~��ʹ��_F�t���T�Jan�	Vj�A}�A}kA5�=e���k��H��u(B� !��sҿO�1"�}կ^A�Y��4��}Ҩ� ��3�q*��SFG��D��^����jpW놱���y�g�����b�BE��1������<K��D�ꊓ'OV��x�477�d7mmmX��;?y",9y���B�k��HII	֬Y�	&��������Y���u�XH^C4��uB㼾n�t6�
�������C�a�~�ۉux5A�NmK'ꇍGq}��Š*T��d&�@�����rbI�r�J+R�%2h���8Kd�� 姙�l��_�2�;���<����Y|��q��Y�1�X���{Cj���+����p������ՙaݹ	^��f7=��nnp�p/��g�홅h'�q�8�x��,[���{�r]�=��nu2c���l�����a�մ�&0����S{L�����D��!㱻��vB!�����w�y-m����}��;y$!��|�8V���Eꁚ��1�]\�����X7T��dݟ��B�k*OrWǨZ�{�XN�ᗙ�l����Ê+��SOQW%
�����J,^�C�!�b��Q/\�z5�>�l�k~^���-��BM1Z������e���a0�v(��l�vD���x퐰+w����N|�CA�2y8��N�����hnOl;Mtb�X%0�ݵ��
VP��Q�y"��Ft���"N"��>466��7ߴ�^^�??�Qʯ����_���w���/���;w��硸�HY��Ԅ��:�����[7��8���6���X�n�wf��t�II-����d�������[�^{C]�=s~�m�ؽ���vԛ�߳���T��ĉ{C}}�}Y;.{���D�������jٰn�D]*�nolhH�	;7BX;.����52�N9��X۽�x�g�����YGE�P�yK{{;�|^ڻ�曻>w���i�'.VS�vq�V�w?�U(?���$���>���χ_�y�������O��$~�$�L��-L���꒰������ۓ�jRۃ�-�UQq	^>�[��B�<�ob��S�Cs��!��P�B�б(�/ӥ��?�S�՚���5�Kꅪ�]`���ؖ4�=Ffc��=7�o��F?~�=�M�DA���]�&Ϙ����5B!Z:���vnݎ};w�<�����q�W�fnO����z�>�hjצ�'�ڵݝk��a01 ˬ���VN��vjz�4��x�D	���E(Y�A�ԮNc�U@Me�Ls�D!V���Q�h��D�`%�����*��vaa!V�Z���zlݺ��~�4����k�~��t���#8������a�СhinAcC�b�غ$�qc�~fӆz���|�E[��ܬ�M��O�e����mm�kO<9vh"���"�Q���v��ܺ����[��wb�M����l������ar>sƅ�s;{��{�޳u#��}%?~apW���3��kMv���Hji��õ%������;���?݈�w񹓗��Z�\�쵋���=�����w�Z���{ޭ�����M|Nn��9�?�8�����}v�X�"T�J�� KaH&TS۵U*QJL�F�c���dz;!��ۨoj�/��!�7Y8��'�@sm�i�gY�gm(����
h�?G��dwy�P�v�!�]yN+qfO0��y��q�m����/��2� ���������EO�?��뵧SG=v�0j*�0a�d��(�DHʉ#���n������D�o���߽��o��Wj"A��|�	�Ų����c�9>�PD�د߽�Ջ0��OzyO�����OIQQ�k��s�}�W�N��D�������������կ~Uw�\&�۽4�[݆�^h��YR7��e�Xj�gY���ܮ���aHq�3d^-���؇w��͝83l,
�*t"U�wm���堚��$��*B$�=�S�Z"�T*�����5k��������S�8�i�&��!T	����ɛ_�]��߽��[���Y��`�ĉ=v,����e~�:�|\dy]m-�M+e�Xm�ߵ3����_����������ʏK�5cƍ���:|���%��uu5vL��zj����/�W>뇍�r,\x�F�k>Z�2����7ld��m��-��Ò%}�����Ү��\"�Ю�w/>oR�!.��;0d�?mW;:�1x�Ю��/�����.���ڃ�[�)�^�
%~}��y������]|�t�������Į��"@���d���0���5"��X�����^�Ҷ���^2d6���N!��FN�4*��B�ۼq����S�3�ݟS���X��������o��ѥd5C�*\��n�R��\��]�Q�K�9�-����{�Euu5�}�]K��K���������kW�~�ڿ�϶O�`��0i�d��=h�����oȫS���e����j���(��p�|�o�]h��ί����]�ep�h~����&�����3�o>�D���طk�'�Cu��v��{�ﺡ_��<S�u�K.�w�u�'`��9����)|X�0��6�ai뇪��X;������A��Y�Pch�.���Û���e�xH�w�+o�IC�\_�`l�ލBUlL@�r0'�N"�*X�q�v0]BS:�.�H�|�'��ɓ'A��J���#K3fʹ��sS�u��s���c2٦U�sdp��ɍ�V��vƆ��c�پ,�ȅ��S��/���a��zeBw~�qq�Ѧ������{�1̛7/#��~������Gj\��='�&�P%K_�����4wM�BP�jдŠ$�]��=,9(RB!���:UB��Զt�a�X՗'��w�Fh�j�ܕZa4�],�u��j�9�5��녑e=�ޗ
7�)�Wy��X�۶mK�_�W���j&~���ӹ��������cJ(Va�?)ڂ����/~����������p ��������������}��w�����w�~���`,��멯���|���՞�[=?��6�1�~�����z�j�������L�3Ʊ���3l�ޞ�vhLmO��9����kK&w]�1�t܉�W�g�FL쪩]�~P"T��wE�Jh9h����^5�kJ����w~E���D\�R�%F����jf7��6m�br��{���B���[���E�(�ŗ^��b��Rn�����F94���=0���-�Ӝ�niG�&�ݹ�&8}_9����8[�e�F���oc�ݱ�>�奸�i����])�8}�}��.��ߦws"�v�H�
O	I�a��v�@%�Zs�����TA3�*:=�?g�)RB!���&���!��~�>�-�����>��$K;��5�Xj-Q��Y��Ko�LE�P���Y0�nK=��ne~���x��'���!Z��N+uC�C͘3˓dVB!�I::>��͔)S����[�n�'�����YV7ԇb�������X8�y��I-Q���2���3q ��wN6��2t�j*�,��'��Jd�?کN����U\�
�?��63����E����+�����f׶8PV��.�g͙�{ι)5�f_��d�M�fa;�ou�W&rٸ��M�ĥc���LHm�tL&vlη�Z�0��؞Y�"Ŧ�?Dc}�!�o��V�x�aV�D��R��A�J�ޮ����������JLK���'�!��^Ms�>B!���,�5�'��j���&�='����푀�x0V�T�'j�T硽v�h�ᰶ~hnrWɶZ�1c��SO��;�Du�w鬤g"��vE;@���\4�Bz7"�}�����6l�r�8r�Ȍ�����iq{?�uCՖ�։��u�X&�C�#�v(���t�vc����y��x�?��,����N2��+B�e�`47�%��R�c����]�Ȑ��.P�c�0�T�ct/���Pv�/��2�t�����?!2Z����__ā�r\t٧Ч��k�̾��_��fa��{��[v�;}����.h�ؚ9���;1�{eX���[:�.|7�	���wM�r�-��k_��o	M~�^���aӇ�{���P�Mk�	U]���B���h�̿{B!�7��ƛ�!�xKus'����ri �Hs7���X�I�w�#!�=Z/D�(�cuM#:�ZgT��Sk �ZK�1c���):�577�#�����k1���5.��	!�":>�ٱ{��dj;1E$�?���J�{&��Q����6����X74N���ꆲ0,i�0��0�7����*j��4���ლ���WI[P[��IdHl;�(V	T�K��������YKd�$�������,N�>����74�S��ڍ�r,���_�0�ɚ��d��]���3�[k��J����X��+���m���9�����	�������c�ؿu�u $W\qV�X�ܮ�|-~M�<�d�L��`4��MR�թ\��TRڃ&	Ʉ��`%�����DWB!������{B!���� n�<�u5�za�a�N���`,s���8�%�#�n��XV��=�\�Y�F��,��1"���;v����X�t	B!���&���W�����Ĝ��B<��#�?~F��3����J���Jr{b�3��9Yr{Bz��9�t�!��*�>���dG�C�=y<B���S��G�D��0%7�dSm�{\�
 2Dk.	@fr�᷁=���'��z�����������ގ�־���wⲫ���a�Ƹ��nѰ�Yj��͚���:6`\�Ny&�a�S�����u\�n�����a��voiin����p������$cٲeX�z�"Ve���Ix=���Pe�ª�=�<�]�b�3�b0
�[����1�3d^-�ٍB�Z�Y�"���U������V�0!�=����cm'�$)����	D��\�gc�{���/GUU~��S�%�����W�b�䉘�x��1�BH�D�@�����@SS1C�������K2�>���c�����>S��k�C����P����ܜ\�}BxB �)4�����!�4~Z�MM��$U�R1�*�R�܍b��^�\�Ҧ�k��[�N�W$r�}�ݨ����/�B�q��	����a�ًp��磠�@Y.�H��W�{�Z�x{f�$�u+cM���2��-����nB��ku~#�Cýt���uK�E�7U�ۏ���)���b�x��PZZ�"��x7��4�Am1�1�*�T��)z�*3�u	R�J�4�b�_P�7��"!��t��O!$=�h�}�x��V���k�j�0jn7���v��l냱������ֺ?���f�.����466◿�%Iơ�8u�$�,���&�BH��P�l��	�Z��ERr�w��n�vm�+2�Ψ�@2S{�$K��k���ڡ�n��c�C�L:?�@k�ɨ�bHq�IF!ğ������r"�~��ܞ�"w�M��T|��փ�yDl#*X�q��`*�)L�ݙ���W:�����o��d���'6�l�~\z��?Q&ZY3�:6���uh��gvjV�6�;����1܇-��oמ�ܡa��8��Non����>aܤ�&x�=��N�7����Xa֬Y���A�e�A=M��H�{��d����Θ@����a"T�.�����B!�dy�9 �B�����e����IjpO��D�9�wM`���] ��D녝b��Z/T-2�NЛC��!~����wp����3�[��֖l\��U`��g�o�~ ���45���n@剓 $������(�V�I׼�b�Z/t��Z�Ϋu���Iz�����ax���v�4���C$24���Z�*�U�����.��VF�*jt�<9ֈ�b-�!��f����X�fZZZ���T4�����#&N���.���ڀ��l?�M�VM�^��XwL��q�o.��/���kej���*�\`�W��,�xG{{;vmݎ�=��{&�?~<�|�I><#��~`��vui�.%S�*�@��"�v�P�
T��Z�W�hn'�B����|B!�Bc�U���iP�G��`n���a�v���?�L����Ѯ�j�PS7��]0Vo�+
�������܌���/ $�'O��_�Ysgc�Y3,�!��q�w�.�پS9w"�
��r����&|�gBm�����y}0Vb�g��]�ʦ��>��X)j�2s{^׵�ۧD�~����d$o�)��T{�R"�V�R���=�⮊U�&w񝠊LF�J����6��4u����Z2APJ�|߾}����������A��W���CX�d1�,]���x�c��X�\{fa�fe��v}>�c�1�;�?��p篵G����O�9�Oc�ݱ����`Yvlފ��6b��#G�駟VL� 8e¼9�B��؞L����#˂��`t�^�2
Vf�����|0�B�.�YR ��^��B�<��m�c�C����eqC��6F��.P��S%�=�^����j�^��熁]K����������T��֮]BR������T�/���a�� ���8z[6|��3g@�U���Z�s�=�ya&����ߞ��.��l|���[�Mo%�
��Fs����}�����X�]�F����%X�7/��`��`0&E����F�{�!0N���ӸȤMo��,'S�#�����z
=��m�B� N�6~���܅>u	�͘��W��S�u��Cs���ꉉܡ��޾`�U�S��������8����?7��l�߆u۽��T%�l؄��:bq����ӧOO�8�&��R%0Ȧ֓�5˂���Xr{�ւ&BU(ԁ���d�AB!$�`�;!�?Xw�7O��S�k�Zs�����e	��j��!�`�Ȑ�F�e1�|���?�0Z[[����+45���7�Q���^�Ҿ� ��g�e��8y�8�ç>�)<��(((�S��x�j��ݮ�qs{0I�дv(3�w��a�g�4������'����2t$Id�&1hS�uFw��=�� �M��b��*Nz������c1b{�1���C�@�U�.�^���`��	���K0h�`e9S����D�v�f�����X{&r�&zc�֏�����{�4�`��-8T~ �إ��T��3w�\WM�~Mn���Pe.N��������v!P�+��B����<;�hn'�B���B�	!����#��dP�r}����ż4�]ol��H��x=���YL�`,��]��;@3+�|�>}�f��\�6l !Vi�������S1{�<����B!�B�o�۹{��T΍�Ò%K��KJJ2�p�	����$��$ݞ��w}�P��������;L��E�x�H>��g�6<�'͆c�i�h�ԜH�)Z�"UL�
h�+��]�� ����U���"ȉJU.�쮁�O}w�;~�x%�S��9y�$������>�y�`�ҥ(*)���Ooj�4]ܡa=#L�����3�1��X{�{����eq��X��4�{�*N��z���L�Aqq1�x�	�w�y�o2APJ��;	�*��=>Ml/��خM`0�����?����'U�B!�ҿ��B�4��q�1<X&OpOR3T��j��Z7Tky�:!b�X�r�l���j�PS7��o0VO�8p��%j��w�!VZX��8~�(�.^�1�ǁB���@,�%��˜9s��O���Q���ym �6+�1�ǌ횺�ݮ�AC�0h��Y�vDk�ښ�:�`�ژ�N��w��|� W+FG[��؞��`�^�JLq_�JkrH�*�4���$���w��Ϙ1?���p�}��ĉ ��k�Ə�s�v,X���,A^A^��[4�{dl�l��e"�s��e��a	{&r���vƆ���!��{�Ą��Xb�{=v��}��MM �;��GŅ^h�$�X�ռ��@�.��+�F�T���"���Ik�L�jz�Y�����#�L�Ǎ�
��B!$[ط�B�_l>с��Ek���@,Y�P_3L��9��92�k��`,h�2�қ`,;5F�p�>O?��br///!v:�����C0w�BeJ!�]��N+����*�f͚���2$m��t���=^34>:�?���ܩ��������5�Ȳ�O�hn'�A�;�xZ::�?8cC�ʇ�,��htכ޵-�)��P���U@��`$`1u�A�e��	M�`TwSH���̙3�ar���0�O{{;>Z�>vmێ��/ǌY3��s[&r�f]�fa�fe�խ��0�;4�[ܗ=ý�qfcәz.ݦG7789&��~��.��f*O�ĶM�QW[B�K~~��V���.�,2e��ӻ�m��d	��vm�*X��0$�T�V�b�s�D����B�f��蝼4#��/��gF�A{kK�F$�j��j�P��	&w��'��f�Xq �eٝ`,;v?�n�رc�`�{ｗ&w�-���W�b̄q��p>����B�3�MD;�lS��	�.S�Nŏ~�#�9�3C��5?�ǥ5�k�>���±��:��%ʺ>��]��V����Gqi_��@. 
��;hp'=��:0y�8��>��nP���UZ�*'n�7��L��/�݅��S�7i�AU�Q�<�&�L�D���Ǹ���Q]]B�CcC#־�
�oނ�/�#F����p홅���7�{a��s\޼V��[��L������?��8u��aℼ�<<����k�
=�`2�{�nC�%s�>�!���O_P~N��`��BU߁���;B!�d'"��K�-Ŀ���B���]m�01T�܌�P7�>;>[��2�
�S%K������̞	u�t�Ǎ����TQQB��й�>�Iӧbּ9�/( !�{t��cώ]ؿkO�7EHw������3fL�0��a����%c��~���C(V�wy0����ʼ!K�-���<!co����^.���MMq�J���A�$wm�{N ��x��>��*m*�����tu{�pf�N�����?�r��0���׃��r��	����)ӧa���0p����c�3�ݑa�5��Dڞ�<��ƙ�������;iin��m�q����q�0�?���4�[�7۝&0��e��v%���ԞL�����ە���!����ۮ[�la�ޣ�`�!����߸B��-;�_XEqa>!�d/{���:e<�Շ�����f�7�'����fh��R܍Y1�ciɄ��߆�I�&)ݟE���#G@Hw�X��8\qg͛�IӦ*��B�#>?E�p疭hkm!N7/��:1�C{wM喙>'��	�R�V�>w�:���s9�'`_9���{hp'=��N`S�P��iR>4#�
9	�2�{d^/P���`�&���U����h1�ir�c�x�b%�A�hr'N)ۻ���c���X�|���{ީמ�ٙa���{G����Z6�{`7k˰nq��1Lv�	ݫ�����ػc�"��sB�"η��s�!�鎹=~�]\�R���L�jZ�i�n�T��&���"!�8A��ʧ�-tt}�|�'��7��}���_�	�~�Y�w����_��&�!������N\?�?Z�u�B5+Y���n�} ��]�����h���ac�Ygʔ)J��=�܃�Ǐ�����ֆ->F����1w�M��z"!�d�{�ء#ؾy�π������z
'N�V�/��������N��$5�d�Xj�0���I��]���X���
�8Hz����(�1u��Ք'��V�X%����8���9�J�v0�� �"w���I��t��V^�IB֒%K���+W����8A����Y��b΂y(--�-���t�|�d�S����N�
Lm�w#��X�����W����m��Q��}س}�bZ%�rss�b�
�r�-i���%@�"q�=�*uCb{A��`0�b0��U�*jr�J�����in'�b���\<�����O��W?�ɽ�Q�ؒr��#���_��t"n�����N�4�BH�'��ځ8��L$A0Z+�e���؀��YMs7� -P�S�!jk��`,��.��Q�JT�զ�g��]K�u�M����E�g�܉S�q�طs7fΙ�1ƁBH��'���ͨ��!n0b�<����M�=��翹=;C_?�����5Ci�g]8�y0VB�g5���i}����1�Iz����8^���#�T{*!�!���vP�̠m9�#��9�85���b�A���"�6�]��={�Ťt����ҥK��U�V����8E�mo��	��맜|�_��Iױ��,kbVv`nwj"��Z�]Im��/k�쌵g"w�n:֖a��X�7b���:S��Cm'�k�v���6�ban��������7ڻ{�^'0����*��bP+RE�������B������oƷ�<^�hH���܊o]�3�K:�W-��������]��Kp�˒�y��x��� !����Dc'��GIC��(7�Kñr��Xڟ�5C���`,�SM0V$K��J�{�:�v~�̙x��q�����
�8������w���D�n��Nc�'[Pu����0���'?��3,��2��矹]�q�E��$]�Շ��vyb0��n���b��>w��t
�W1L���I��#E�lh1:�ڢTb�A�@��7Ot7�1���@6U�ʌ�q�B�v�س�@FK^��.� ?��z�j&��'g�� [�.�.Y�9�梠Pot7{�[7;5+����Dn��k[4��7܇-����ü#s����-ý�qf��	��mX���]c��r��EsSqq���_��=3��[hr2/O`�$.$����`��)D��D�Ǳ�iڃL` ��}���W܌���Oi3A�tt�K|�g�c�3�FQ�y	A�����bǁ�8|���cz�㮛�'#��>�<:B� ��=�{8����FK��x��f���.ꆱ4�@@7�ĊeɃ�T�;ľ�Bc0V�t@�	�f����E&��gϞ��E�{uu5qa�lmnAmMf/����B�����ؼ��� !n2r�H��>k֬�4����n�.Q녩ñ��v�`,IH���Ϛp�����J��$���Nz$g�;�?8�:+�mL��y�@��"�H�;���@�ʀ�(�R�úm�m`�û�e˖)�=�M��UDz��＇�?܀y�b�����ݳ�v��iJm�gwf�wÄ.]�����n��L6�Jj�a��QzeX��=��;�8z�0��؍3�� �mĹ�+��/|�Ss�ߦt�捩��H*��v{	r�J���T�����.��&����vB!�����/��}�y���n�����U��o��Ƿ^�t܀�"<��-���ߢ�ݛs���"����I���N!�͋�}���"��lV/���1�����������Y���x�~���?�ɔz��ǔj������<� *+�2K����c�c�ј5B魈.����у�A�ۨ��~�ۓ�W�P�&�hl7Io7Ȓ�u�X��a�@,Ӯ�Qs{QI�t0I3�x�ǲ�T&L���Cq� Z%3�'$o;(0
V�w�f02,����{��ݎ��t[�{��ʰr�J��y�E����6l��>Q���-@aA<���,l\�Ԭlc�w&�L4�;�8�ܮ����.��9߳�v�64����P=r��v�Qn���M^^|�A�x㍮�ۍ�mJwk^���x
�F��el��.�$0���*������c9��B�C��u�͸������3x��MX>w�9ﬤ��N���~��_�ۗx�}�B��������BH[0���C1-|P��5��ljv�	Ħ9ڟj�F�{��]�cA�����fBݯ;��t��Ν���E0ֱc�@����N�ʹ����w���N<c��ъ�묳�J��݈�uA+�zc���.��Sw~6�
F:=�u�P4 +dRC4��,�ak��.�I�����h^��������Z#B�[�	V9:�*� V%��b�1�]��F�X*�X7.��{o2�kq[�:�s�ӟ�T��z�xA����f,<{fϟ�$�'`��n��끉<�؀a\��lӥ�s+���zps���7녹�+�<1���<�@Y9�l߅��f����/���W��n��W�(��{=���ęU�������Tg��P0h*Pi�j*�(,*�ߏ�	��^Zۃ�#(��EIQ���N�4�� _I�����?�u}��T'��~H�����7��>~����n�h[ڰꗯ(�8n R�����I���N!D��:�)�ǣ�����sN�4�d�H��1�]npW�\�`��~���y&w;�t7k�"��g�Q�܏9B�Fkt?k�L�;!��&��VU���	�x����s��i�|1�gB���v5��v}�c�C��Za(	��Χ�ʻ>Ob�g�4���0��}�KK�TY��*P��D�J+\A3/o;���݅9��.�H�q@k�Ӧ�G~O���3S�J��%{nѢE�`%�B�z�xE[k+>xo=>ް���ż�PRZ�Jj�U#�w&r���S�}u����wj���rhηe���ƄNs{z�>��+�w�0���/),,�#�<�����U����N��V���I�Z��?Sۍ	:s��H��;$U�����6�T��n���w��/�G& Һ���)ǉ�{�o�w�M�q�d-��)����z\~�4�:y�9��{nT�_�g�N�̧���������@QA�r��?�W.��vҜ��;v؀�chn'�b���N�2y�j+����Qc��!��}h���=G[/��]SY0V$K���&w-^��O��c	����L�%ޠ�G���sgc��� ���Bu�i�پS�����x�ĉ���'ONKMЈ�fu���0,Ӯ�����e'�]]�a5)�J-1U�gY��!���2v�'�A�;��T5�pr�Xj+3Mq7
TV�*y��ؼؗI*Cm�����t���y�#ar?u����v|�a���>c�Y��x!�W�������s{�|k�1ۗ����������n�Dnzs�l}�XK���7������!�|�~�߽�� �k����f�\y�=�ܞ��TI��p�Zv��Z�d)�;h"����N!$5w��_�Ζ
�n�-�oj�W��/<�K�Γ���܅n���v�d>�+N���7�+nH9v��H4�B1��%�h@�r���fh�^7�[�j��z�1Kot�&w7넩�%B���Q1������8v���2l(��>KIv'��L���
{v��	�S�*��&LH���o���y�f�7��S�e�X�k������
:���ϯ�㩿�����
6��SƢ���i"C���wS�;�r�$�AO<�A]7b��2\��=7w�ܘ`u��Q�%��o���c�X�d1��8Іa�y&�a�u��pj7kٰ.]����2gϠl�^�W�|F����s�W\��B������ԈT���!s�J+LY0�ǒ�%)����
B!���;ۻ�K������߽���<��OI����V܀����m ���]��c��Ǫ/]�����N!$)u-!0
Ãe)k�v��j���]��Y�*)��h0VB���jlW�[�N�/���4�O�8QIr�X���!^r��
��|G	Ě:k�Mԛ�!�/�w��cǱ{�Ԝ�!�@t��cǎMKM����0A��Y���!Z��v���h�0�P;4�ծύ��L|�w�kx�"׍폖3�1I�n0���`�vИ�)�iE*�pe��5�DЦ��7��H&�C�܌3���z��I�(߷_y�?�/���l����~�O��f��3֩�ܙaݖ�܃�\1�K��oB��=}�V��w�Q�b��$�_�~x���q�d���ܘ�S�O��0H�Z�E���ݮ�]��`La����ۧ"��3�B��_X�֎ ���������N�����4���ן֡��߿i�o���wᶟ�@s;!���l>�uS&�����f�c����������5Cm�PE1�#^/�w��MF�����3�Nh����0a�y��\��v�!^SW[���>���1e�tL�:��� ��t#jGR��gAH��9s���>f���xF�c>�}0���.Mo�P7L��Tj�A��v]r�!�=g�$l-��������	���������Pe�� �?��Z01�!�t�9�w5�!2&"�DZ*si7��axw��.�܅`�o�>�.�:�<DB��ys0c�,�(����v{���p���Im�n��e�:���n�po:�_�:��CM\�EKAB�������SO���v,JqSd��Ю�W�)��].Ti��*�H��TJr�=s�Q�R��b��P��B!�m~���PR�o��-L�:e�_on�|~�oo(S?L�"���vB!Vy�<�'BsC��f��J��n��ꂑ4wm�P<dI��pT�b1,.��7�H:���:"9T��V�^�m�x�$I���c��]�2s&M����BB�״���B���ݏ��V�N,X����1b����tڽ��S��I��G���#?%��!������ϥ���r�<Hf@�;�U�h�x���T�,�4[�}���P��� ��RD,$���S""��j����=��[�L�8?����裏b��ݰ���^�_�Ȑ����}��/����/Ӈ�݋��n�vqb����رe��<


�4Jm�mhmnQa�/����@юL�������K�HuHb�¤kwg�_��Ȗ�߻��MҒ͎������^�{���ֶk�B����ZT��oe��mZ��L���=?h�������[�345�Q.
��ٵn}]]�{�F�����������~~ר�t~���گJ�wQ7>|�r�5{�l���q�"ju_�R���ZIo�	VR�J1�����O`��O�hn'��"��_�"�q�y�����{WaK�q��G�܋
��k�I�>��N!�.����+�ci����X34v�R+LU34�
��X���`d�z�|zM��zQ'�Ώ=ZIr�ᇱa��.Z[Z�㓭صe;�N�ig�D��@!nS_[���p���rBH�Y�l{�14ȳ�^wֱ�]��!��k�� \��j�0E(�xN���R~��ۃ!��X��aA~>^?Q�u=E�d4��^Ǧc�v�xt���B2$���%�OhD������dE�RS�)�P��Qѩjt(_d���v7'�ūQ�F�駟VX�֭�T�W{{;�@��kէO455�����b�����W�����br�N����c���	f�ƆT�>��&ꖛ{O%&r;�p��;wc���}���t_�Ǌ�QO����Im�.��:�|.>�z�y��k5Mm�"��M��X7X���?���M1ۢ-�ݱU'O����O�R��0�O�:ٗ}��SG�c����i�o��={#�T�Y����������[+����ɼէ�
?_��������a�ԩ%J9]�+,�6e����zc���	T����`4��O����k$�B�����9~>�P~}"t�A�J@zk~�w��𭫗x�/��	!�t������)�?�1��5ø�]�hpW��S������jz��{_�g/�2d~���'���~�-Q��
�;��p*?�R��M�i|X��K�1p�`���k�+�P,A]M-���ǀ ��/�kk��RX�]�kp� ̎�MMhok�e��&���v��3���]����[�練�������x�
D�.�����~�
��-�X˗/W�唖�zV���:�fh�����O�w~քbj��S�������ۃ�������	�ma0�hp'�����i�`45�F��I�)� �A�BJLd0�S���F#�Ơ���v�����='�-p�c�ڵ ��{rߞ��cА��9kf̞�u��P����[2پ����Ec�sý��`q����f5��e"�e��3֡�^:�}úW&x�}�<v�w�E剓 �ofΜ���Ǎ�(e�?�z������v�Im�br׊R�H�.����w�e��`x�"�k�K���F1һ7| &����f�8��߯��8g�8e~�#hmwv�!�������m��y��U�{��տz��TaΤ����t]���w��{x�B!�{l?с�J0��x�Ϥf�c������;�k��iL'HHqWuUu���Yݟ��V�q���S�E�z�)���˰BQQ�����g0�x��_KK�/��;,ī�����S����~H�&MH08
��`��A�?�������%�}|�����o�L�J8ըqc|�����1b�(��tS���;aN�����<3���J�P5�;��~�Z�� �>� �k��ʕ+�s&/k�n����)��Wk�zc�$K��9U8V�`,%KIp77�kk�f����8;*hn'��W"��=�l�����Z������[�փ��t)�5��p¶R�n�ʭ}�5N�??����U�򗿀?�9]��＋M~�ig���ٳt) �M�f�p���������>ֱ1��ذ�����5,��?�7���nѶT$���݇��f�	,\�P�ap��ᾋR�Yǩ�ݙH�OmW1ڭ	TZc�^���/%���)��U������V�T�wq�����7�oI�F�?؍5�Y�cU��D.Y8O}�JL)h�>T�����n��靈����X0u4H��w�~B!$�y�<��'CSmUb��]c;��CM�;��c�t�h��R7�uYqTc{d^����v��v���5k�(]�_x����7Dw��mĎO�`���4}*B1���������v0����?�y�X�B�Q+Sk�F�7��KL�>'Io7�!&�
�܃��ꆚ�a���c&H�A�;�Եvb�(��<�|(���bL�����Fw��] �'��6�|�i�ܭ%2$#BV&�܅P%�-q��?���񝶶6l߼Uy1�ƌ��c%w�;5����%��7����Dn��ō�2��2����p/�	��v��'��Q���U.:	��-[���]���:~	\qaJ�,ǖwjR�%$/�甶�Am�AU�
�No�̫bUp�$�b�e��Ogn|f�L\0o�]�[�<�I|��%x�[WB�Q5s�0��W�;?��l�s�wB!�������b\1��m��ρ�4�d�CH����XO4ܣ(ݟ%i�q��B���0��Q'���Hk}������~�;�'B���W�<��S�`������!�tv�8?rL���3�$�����{��r���2�&�t}o��.ϒ���>�=Y�0e0��Ƃ����=duC�(*.��G���UC�o��Nz5;N1v�xt�ԋPI�)�p�D���-�F�2��(V))��id�jt�orO&�h�$�Jy�.�G�5x�]w)���}�Y�)���B}]v�؉�fb��4d����V�E�'�'�NM�Lm7�=Sۉ�3�gp�� �U���t�ȸꪫ�j�*%��M���8��(#n�TZaJ�b� P�����FD*5�!"P�-CJ�{|Y�ʤ�`�����r�n�%���י�U�u-�6fH���L	����уAHo��x5!�B���-��#0��@��s `�t����;�6��?��v�x�+쐰)Ф(�B��=K

m�(P6!�UF_(e�Zx�{�@�jl'�^v�x˒��邏�Nw��>Yϧ=t����$ǖN����~��.���.�r����z�\�Rc���,�ǨkkVHu�{FF�=�\��}����7"$��t���#??���M��((*!$��ڵE��K{k�t]B�]���wu�	'H�J�T���H�z���js���5������ĶөNm7��,�d���a|3X5�y��EĞ��NF=�Z�qt��q�zC��l�W�BZ���G�R��*훟^��xc�\����G�h��=�w�#���>UUU��[�p8@�]�7_}--��J�ݎ;`�v� '7W�o�Dn�ֹ��#Rzhc�o46V��ǆdX�8��qY} z�&ڰNc�9"ma��.���2m�ؚc�=�w�����fn���%�Sjc�B��S�������*c�,X�*Y�r���z������6�#������� �.�BC�NB!�$��nr����m�n���Ak��-��;?�F)�J�{���9��+6f�D�詧�*%��~��� ��U�W�R�k&Jan���ːckV�B{�2��-��͕��~��1�Z�:��j���v�H�۵�X�����r9�����⚤��	��4��B�;I	���Ay������-�He0���*�H%�*���5�GSp��������xΜ97n���Zlٲ�؍�M����ه������v�v��ﯲ%�Es{�l�&�P�F�0��s������P��sń�:��ƈ����eXٶ\*�����;"���:�,��`�[Zm!+ZsY�<��T�R{Au�'�����ss�6yA^ă����CNB!��	�BI4o��0�y�;ש뀊��1���������u�:�ۛ����,cy�%O��x�8�s<�cPYY�����5Cb;�T�o��
�k��8��@������X�b%ּ��bG���p�Wbƌ1�Zs��Hj�ʚ�|�.�U�X�Zb8�}�X:�C���ҭN�P����k��R�.{C�;I	z�����b���`e*PV�m`*���J���Ms����F�cl���]�]M����փ�_~96l�W;zBd�貖Vi)(,@�6۠a�f�W�������O�z�&���uǆdX�8.���s��	=&�T�gk7V,[.-b] ރr����w��K/�!��ւV��UȲz>�ߢ��L��k/(�	�In)�3��R�v���BO�H`�HE!$��ݴ'r�(KB!$q��<��/�@_o�B�АC���v~�� /ݣY�k�R������E��?ۥ��qӧO�m��&�׭cj.�B��b)(,���F�75 7/��䣷��m�280����ۉm����u�]�)S�Ĵ>hu\<j�њ�_/������ImW������|Fv���nnn�j�y#�/�e��aC�-`%��-.T�5����/@� X
�J)X��ƕ�MeP
Wfo��4w(�*��M�b]�	��EOd����cB�������e�]��K��;��݃%_-��¢"4o���n;���-]F���i��9>&x��qKm7k�1Li��v�0�=|�����#4oڰ�$eee�ꪫ���Zq�����]ml4��R��U��v��@��\N�}����J��A�sB!�G�G�X��Ԗ�B!$Q:��bk�f�y��B4����c��=�=�����I�}j�A���)�rh�/�@�Sit���]�Us�ո]w�,�j�--- Į�tw㻯���K�Eiyj��P[_��lB�ːÁ5�V��u6���J��	�+;�#���?a�ĉa����E����KknW��C�P,�ڡ?+0�%�`��X.��v��azF:>��!�0�;|%)Ň+�0{�D86��ܮ�` ZiR�I���u�X�V�T��<���4���(�����p�B��Β%K@H2нu+���KiWV��m&�y�IRjS�Ck�𘥶�-�38U��4���E)aj_�f��!��d�n�V���x���^j�����`)}A��`�^Л�>r�?��X�r*��}%�x��B�mX��wB!�$�[\���GY_��g�1#��%hQY3�z�6�][s�Q��)�B��f�X������<O?zsk�4i��\q�����A����"dG,�|��U���Ԁ��Zdd��C���ڕ��޶��C�t�@,�*//�g�/�u�X���vm�0�P,�`,�v������N�E̵&s"�v3�$��%)ǫ-i8��}[:B���o[���\y���c��B�ʠ��'�*�փj��ԂM���UTTছn���_����$��:���O>Cye&66�q�fz���10��*�=n��n��ذnql��|��z�ƎV���NFF��T7�k1�����-m��"}a�zr�����S���z�vi�SJ�{VN�\W��B!�.���!�B��b�f5�c��=�.h1(K��[3���:���ʘi�w����1�����B�[�|��u��7��k���B��;,�Ų$�KL��Am�DT���|���!4~Q7\Ѷ\
�FSB���3g���/GAA���V�%��.�c`n�	�r[�k���c��vhhn7Jpr�=��[��E��I��y����<X����J��nx�O����4�X�Oe�o�I"��X��V�9z���+紛x�1�X
V��ŒX%�>��3 $ِīu�勏?���'5���	E%Ŋq�G��Je6N�=��qFc�����c��n��ݛh�z����X�zM�d�0m�4)����4,q�l�h0����򺜾�m+,�A?�]���i/('0i1h R	��BW?E*B!�b�Z�	!�b^ku��*�u���C���5��!������2�u)����%5�x�+**�7܀;��=�I&���޶LZ233QY=�k�Q]W��Z���#o��׮ê�X�r�����d���y睇��,[��=&�㭝�_Ԛ��B���cik��`,o(��klw��U�v��aA�x<�B�I.xuKR���n|�W��ۥp]A*�p��U��,V	dQ)M��}:��JNv����j�{�D�h��q�O�`_NN�ϟ�	&`��;!Ɋ2ٽ���M�k���q�����c��nuRc�}�&���Fj��?{LL�LmNOw։�����ظ1ed�1g�\p����K2�O�*��#��/LI[P�����e
��8e�ܮm-�Kp7I`P�/hD*�s[�к�׺�B��'߷�p�ٙ���#�k6mIr�2p繇c�m�a'����7����@�G]e�GG'}�l��!���<��b��ǴF(п߬f�4��������r0t�?�!�z�@]���=�Z^(��D�����/DYY��>����Dh�"�G,��?��k�뤄wa~'���0���9�Ծb�/X��dE\��{�8��c�^��j{f�en���]��6��ە�XnˡXz���ڡ���:uk��.����C�+,�K#�{I6hp')˲�NT�L���V]1*����m�4����܁�7�1
C�R����^�M��2����l���O<uuu��k���B������E��s��P�0�#���jT�}�V��0�GhX�:�;����o�T	7����[<߮��X�j��l�`�$]�k�y���SNAzzzL�'�s�K���\������j��G��On�����U"��e��n�d�����	!�ؓ�Vlĉ���^r��1�p���^ŏ+6���ń'.�5�Mi�y��0��'��+A�AfF:���8�gۃ�Y�ُ8�ƿ�bF>B�����K_"V#���v~V��KrW�jס������v{��k�ꚡ�h��U'�w�Phg��~:���q��ף��_>"ɋ�庇�ݮ���	���mvN!�����DJ;;=�ф�^s饗b�̙Q���K�Q=�c��+���._��bOm7KnW�إ��r����v����>Q;��sNI6hp')ͧ��8��C�jJ�zPF_��jS^�
aK��.��
V����Oq��*2���.�����*U�NBT4+y{���X�`���J������B_~��i����rm�D���kF[7����n5���o�	>$úű����n�\����p8ذf6�[�5+Wa� ��Fd�ꗿ���K�~� PE{\,����v�X5�M\P%2�ۇu�)��]���t��+���:K��2<�*>Q�p�B�	�^� �4����C�~�4���l.�۹v%+3g��6��3Es;!$)X�Չ��ZT-�s����4c����.���P3Ԇcy����n�S�w�ۃciI�:a(��QO<�����Ϣf�b�
���q����"(*)���jL��W&B��֮-�/�lڰ��6jkkq��bʔ)q�Z��N�v-�ڡ:�s?�uCM(V���q0�6K�jk��±��� �k�م�$'4�����a�T��΍~Qʤ��@u_��� h[z��i��e��PR�;�b�[ό�ڡ��nr�Q��<y2.\����
_�5m�٭[����>����QZV�ꉵ���AyU�d�Wb��n4������>Xk��,�M�a}�����ذ�׮�:7u���LHUU.��2L�:5*�پx���=&������v� ���D*���/Py�+e��^��P�kn�?'/o�.y<L�!�b��o���n��ogs�?�ً�4�B��o�:1�i"�|u7+FwM0X�л#���B@��?'��]�Ь�w��W3\�d	M�X~���())AgG�dx/���2�z����v��[�FJm'd���{H�6�|v�ZKs�q�P���P,m�мn�2�҆b�B����N�"B ��5��6��I��+U��$�E+�0�"��}���`B����h=x*}���Ms��X%����C3�kG�ūP��<����jjj�$��n�	���:�dTӱi��|����kJiy��Q3�cǍ�1Fj"w�1�p��a=s{��{���0��jl2���#	R"�}kg�n�
BR��w�]�D;�x
Tј#��h�M��ւ�@�1�����{o���T�P5f�i|�[��A'!�B�I�ȅ��<�ڌd�o.�+7nAuy1!$YX$��&U��cm�Z�aѰf���ѕ�U�۳;����L�J�Q'�em1�8����>�pz���n�[o�BF#BOl�o���Za��T��B��RVY���dG�΋���"k���~O�hgƌ�?>
�^4�g�:b��|.��]��9�P,m0�����t�nn����j�B��$^Bl���W=��9k%����*x��r"��\���5�q�}�u��X�ǟ���=R�)�BT(iV�H����J<�� $�G>���O?Gn^���0���UU(X|46��`հ��<4ý�qF��&ڰ>ڌ�=���q�zlX�}���}��� $U�5k.�袸Tf�!J�s����MaP-r�A��ւ��԰"}����R
Q��T��6�7�}#��B�>7�y���H�oq�[�bnx�m�t�)�\�B��yyYfO(B_owj�r�P�ߚ�D��Y�v�_p���9��Dc\��D��0�766⡇u�:!J�����SZ��7+;�+QQU��	�_�ZIN��X֬Cff&zuDBF3���8��q�YgI��v�Z����q�z��X?4�2�
��w~��c���f5�`����b�cYL\.�$4�⥽˅�	Q5���]Z���vT�����e��*��8�4�!XY9o��ą��~�;)��[nA__I%���}����,�WV����U(-/Hm��z�1�plH�u�c#5��=��� �1�c�Ftl؈�k֡����2�5��3ΐ�F֎��9kn����ܮMafn7N`��/�]N_p��a��E{A�6��V��	!�}��7N>x���>�a%�uv#�8�\����؋�~X�_�T�]"��d�1�����W�������.0���=�jñ���r�g!^�[����#���پX�q�Itk�Bk�7o���q뭷bpp������U�WH����PJu/KU�.DlJOw�T?ܸ�!
/!�@nn��u���^�*�C}��h���S�������"Ky_��XN���kvW�ӫ�۳�2�r1��$?4��`�!�Ѐ�ͭH3Ɠ�` V�&'2��Fw��.��`8�g�����'��ڂ�M�b]�q����c"�C�>��={�l�����C[�H��t`����"�Uƣ���W^(X5|Gj"7����#2�GjΏ�	=&x;!>�uut�c�&tlڄM�7b�����Ÿ��q�A|��.������v�X��Z�{k]�
L`P����)�0\�����k��R�S%��dg̘��S���C!	f�]�p�)�:�1��'$�9!z\��[җ "}��َq�!{�B���n��3��e�&w����f���3���LMHr=�J�gar��e�/�j���lΜ9����j�k׮!��0�eyK��-�A�V��ld�XcKǁ�D��Z+u}&$թ����W^��w�=�B�}ў#Q�v�h��҆b����͂�ԡX�ڡ�.h��4����{�EF4�����9qDs:V��z	*b�S��%b��KRʖ��o�R"�ț���b ���c���.���eeߔ)Sp��wK-?��CB<�+�-���b��.�,az[Z��#5���jV7�8���!�{��a=���@Wg'6m��Q���7�	ѥ��W]uv�qǄ
Tf��������J�*����@�m1����HYp9-e�*��v������ ������=��w��ڎ�&`��d�wG�Bj+Jp��DzC�k؍��~��vb�s���O~�x���ੋ�^��t>;p���Ď�� �$/?lt���%=��:`�:a`��5C�����<4A��?����h��徽����w���Z,^���2���Lx���Eiy���-+��!�Dh�;:�)B�F��M�08���(�k��p�e�I&��Z�:.Z�vm��(K�*�����`,U=�gl^;42��eKa3~Z9BF��$D��G5U��s��T��R�J�������+�7Y(E*]�J�S)�x�e�z4��X	V��UUU��o�=��򗿀Ȗ�-�������,��t��Ri;N������î�bal��{�a�1��s�HU�ҹ]�G����� !$83f̐��E{d��can����ZjĩP�����~mr{0S��1���Moţ7V�9l��{B!�_Z��;	�/}��:�����/:S�ƃ�6�Y#�G�� 7��^�����؅�]�!�=�p���Nt��>Y�ġM��l�\'ԯ%��k���>��B����]{�x���2N�z�vκ�:�y睸�;��/��At�Uv�/��E��]$���,��} �9�]��E���M��N��c��y睇��<�55�v�k{ј#u�P���n���2�V%�����b9��|�Js;]��N�B�yey6�.BOw�D�Ȣ�^��g�˻\���ъU�M��f3�{��	��OolNN�9����㦛nB__!�8X�r������zM�e��U<��8����=ѩ�FccaBOVc��=�-]]����eC�0kBB#=='�t�͛�����Tf�%^��ܮ0�+D+���<�!P�2Kn7j/(��>arW,���eO��øC!$:4M(�3W����|�[�?�T����1���&r�ɿ���	A�}�t5n��� �BF;���qԤ	��X�>���fx��ݟ[�9����><����5�"\�{2���!�FͰ��@JF�f�m$��� Ӄ	�"�f�vm����e�}���R]���XZ�R�1��L����������)���#:��J�%���.��9s���h��b�Ϯu�`�ve��j(�Y0�6�ݿ�
bb7^�˪��R~��>hp'Ā'�A�8�S8 ���P�KS�������,UG���
c�,P���9!�����E��hr��>�v�a����5�\���vB�#^�6�� -J���%A�d�X��YJJP4�Y��vӖ��~wk�vC[�ű�2�'��]�����{�G��:r۳e+�n���(PTT��.���կ�A�*P���]~U0�kZ���0lA�
������ �2c"ڻ� �2�ر�/�p
�\��o��9�r2�ĥs��@��6�C�:�w����x�6IلBH�y�5�3q,��v�
--�k�i�z�<�}A�?k���Z��/�������j&�h���_��ט8q"���:�]��s���i�Fi������,E%|vv6��D���oDOw7�:;%#��)2���𨨨��W^�}��Ǵ��ݶK0sD�����ܮJm�1��c�c���=�C�3��v��XP2/��LF'��&Ą�=.��[�F,W��C� �X�6���Ղ�b.e"����6-M6��s�E+y�d�����'oO�:w�}�dr���/A����^iY�J�ʼ��P�
E�C

QP\(����&x�8Sۭ�C�{�v�Hi
==�[af�����7�������&\u�U�i��l%P��øP��򺮹ݻmM��7��t�,P)�����r��	!d43��/�x*���)���鹪���Km)���~J
rq��g��2����t�BI���7�a���dٴ@���^��$w�~�����q�F.����R�����ќ��|��gt>y{��ƽ��+��,YBHh]U$v�EIfV��I���zaq1

@�|%��[��Xb]d�I���~�	�»t��W���.�^(cen�GQ������B���:�X.ej�y�0�۳�v�����|Nq3���Nhp'$?lt���%=�*Jm`N����|��/Zi�ӛ_Nd��vЛ� ��!~�E-Zɷ�`r6� ��������]w݅�z�=�X\L����[��X��_�
�'h!7/y#�"�!g��]n��������L��}}�"��==ҿ����[f̘��/��������a������]O�ro-^{As�rqh��J밨�!�$#"�z�M�y�
�Uc����w����Z��$��o��a_Z�q�>�Qz�#��Y?�e��A�=��7x���BI5�����
�3�=�X�j��f��_3LS��60r��8&�V"b	�����h���U3��)�w�y'���?�7� !$r�iO��.���-d�����/�-��f��ė���vw�{d������&��E-�9s�����/�M%��>;��ܮ�'Z��ܝ��v�N��J�зx��c�����Jt�3��^hp'���t�Цzu.W�K�~#|��P�o��`�fl���7�+��������Oo�H%>�s�����oFg'Ӫ���P6��[��S�}
û0���`�V��fdf�9�Dvn�s�G��s���TJmY088���~i]�O��}���^���vB�A���֩����N;YYY�5���/��v�5���]��`��n����&��c�{�b"V���s��[��-!�{�v���sמ���c-#���{űx{qn}�}|��*Da����_�}v�έ}�����G߃�NƤ��].}h!��Te�f'J��c�`+���*k��BE�PB�ˋ�-Yc�e������J������'R��=�mr�Ƹx�(����p�u�a�w��@�>��Atl˦�}�Y�RmP,��y��37/ϳ^�/ൺ11F�Ɖ�܉[����W
����ꮄ���7�v���裏�y�d��vh�q��9xoC0�{;Ak�=+��5À`,�SSC�	Ͳ�%�^�Q�U[�@�h�wB,�j�s���ױF��e*�Vz�)��g+!N�$2$���q�h�Yfs��+��3g����_=����]B����,X�OCMZ�H{��͑��"R<K�d*��ʔZ ���v�ȭxM��&�1H�H�AE��.}�Y�*#��Q���!鹉u�����W�ş}A�:!I��s�E��?�y��P�&�x���B�B�@e�^Pafwi��J�IW��i/�_T���sC�r!���b}��/x�⣱�v�����k���w�F��؊����}'����A�Fާ�F>�de�?��{��F>�T�b���J����.�6v���.���翣��B!$��z�J���`\�Z/�����a���W@�PO���&�a���4���]�#i!����-Z9o4��OolFF�Ν���f��r�JB⇨�uun�=�����˗j��6(��R�07٢F��#m���ъР�җ� ,����R��>)(�uEB�ŤI�p饗bʔ)��&���1��8��]Q?�N8���~0�q�g=�z�P,����,����~F��!1���8���]�+-Z�'V�o4�}kҢ7�v[W�&�`s�aV�D��~��q�}�a��x�@I�8#�p�8cFa���"BF�3��#�+�ۥU!�9�oҪ͉��[!�mq��c�f8��RA���a�}��%�\������Nњ'�sDz�`�vY�����[k�����ւ���ZAʡ�^PY�Z_�A'_�	!d4�~s���	\u�/qƬ=�JflS[.-�d�5���6����p�AR����;���Vl!�B���\�=i"�V�X�3��y����ϊ�fݟ�Z��5�[q��8F���4��]�����n�/�j������}�������3��}B��t{{z�%77�g�#=#C��yB������Δñ���R ���c�Z�t��M��Y^<N��%���+�-��"K�';Ep�'KQ����)��}}} �$��bƌR0Vyy��ꁱؗps�X��
��v��v��v��}�5[����%�7�:��T�X�bz�D��b�剐��˝�WV���b��l����Y���X%�T~�*����.��&�{4�	�[XX��.��'O�-������ �!�yj�x}���!��!��D��9�#	���3Ϊ�= ���*P��u�yr�YCff>���~�T�2�y���7����p�y��� vd�����m����@I uX�ُ �B���[ܘ�4}�k��Bx����a�qP����0�~��uQ#T���55C�^(��&w�]�F���ت�*�z�x���q���K�!$y�%�b�A�_����7_}mx�X�V��B�����78�䓥����26��A�sDfnG@�PU7T�CKn���S�=uC]�u:?�M��K�DBR�		�'�ֆ�?nHj�$�JJ�JO�ҊW��Ei���ʠw3��d�O���.Hf���|�̣7V,�g�Fcc#�������B!$���R���P�LV��l����:�j��X���خ'L9t�)���?�j�jK��<!�؛~���A���#���u�o~��.�6w����B!d�#L�/�e����г�S�O*�i��Z�j��z�z|�=�Lir�Ɗ����_h���
e��"����O�v�m�믿�֭!��s��,B�����_,u~���ݶS]1����ncs�\7��jð̌�RJ����21��u}XF�?�KJ�b+�$��o<!a��_�T`��U��R�R
VZ�J�R���&bbmr�:.Z�������X�G�)�"���;��{�-B����G���L⹋o����f$�Km��=m���{��}�'��ً��,('�T�������߼�;���Ĺ���0_o�N��]\7̟?_��\"�졌����9��#1�%/��*��]��*��v=�J���sn�mď��@!dt�j�q����1�p�Ȓ>&1א2Α����~w=�!��B!$�^YU�Y������ӌ�?k���ݟ�8wh,و0���
�Fݟ������q�d���x���?�	�/���Bh�@�;��n�Ν����5��G�!$�T�����g��$�D�މ������V�s�=q�e�a����b_2����XúF�p�>��u�y�Ex}U>��mIjA�;!a�b��ٵh�2�DO�� ^��E*�`�qh��.&�h���>A�c��eeeR���/���o����P�ݎ7�:nn.#b�lǘ��.>�����@B�/~/�sO��]����l6u$(A����|NN��X�H�ss�5�/-,�������A��&+�]�6{�8�쳥ߕh	R�k�}�6��/ȷ����ݥ����Q�-u*��2XҀ/���N!��k؍[������?������C������M�ZB!���㝍c1}���<��ݟ�5C�Ρ\I�ޤ)��v��Z;4���a�7��k� Zckjj�`�<��cx��'uCIm�M��5���D�_6��g���;M��"e��e�y"�ŹU�N��]��\��¯����x�s�?�x�v�i�Aj�0��2֎�A+���06�{������j��QZ��0,E�g�w;;;�m�^G����$
�	���68�[݈��6�E����)S�*M9��1}�J�� �b���"�w���<�#�����o�w�}B!����*���X�Ad�n�6����4������t�,�]�;t*������[)PBH*��+1��p���9�!'+>�m��>���x��/0�JL B!��d��o_eUbJ�*_��\/��Ú�����Q��J����^3�+�`�͛�����rV�^�;V��!���Y*Q�O�sO��Δ�?{�7)봉 �=�k~"��E8S��'��NxG������,��uuu��������P�&�>he����$�]�خ���h��\N]��Q�P^���1i�z`<6�&.X��DB�;!���!��P���eҶO�J�Or74���	������`&w�خ]��`lA4��k����;����~�BIM�u�hK|����v�
Tf�b9.�v3c�O�2I`0La�Kn&��%�t�oI\�B!�g���mϼ��}��LE��q1=ߏ����-A�@b
}�B!���.
*jQ���ݟ5چ�n(��69��O^�����m^�W�0��+����ӦMCss3n��V���{���BI=���̙3q����"f��P�M�:��9�)������:>�t}�����!���X�ވe����.4��Y����1�Ѯ��dCS���4���U�@%t
WJ�� �g�B�D�H,�vAA�ϟ�]v�w�y'z{{A!���A$!�|��8��ӣ�V0�c�/�v+���6��jH#L��e�J�ܮIa([�Z�A!�:���?!�BI.D�������k����oB�'�!�w���c���5C9�R�x����.HthV4�=�h;a�)���g��]w�B!��&���8��3q�	'HI�^;��h�ۣ��Y��vq(C��u��M��J��IjC�;!Q��7�4O@_�i[����1��ݕU`���خ$��_q�L�;
Vf��h_$c��%�<�l����z|�� �B��gҤI��K�/�E"@i�)^y���=����͠˰��X��vEC~Q1^Y���!�B!���瓕C��� w�2i;�[/T�e�A�P���ݻ���]`^3t{M�z�����ܵ��ء��X+�fdd`�ܹ�~��4����BI�5���^�w�1ej��#��ve�0h0VaX���55D�XJ��2��	����(��t�T��΍>�J�ʠ$�h�_3V���W�h=�ݎ�`ξPK(�h�Z=Vޮ�����#����.L!�2����g�ƹ瞋�c��M�
��d�onW�/�	T	^�J�ܞ���7׏ŀS�EVBH��ï��WaM�V؁�vn�!{oB!�B���_mØ=i"��}z�Y��s�A�PQ*���]M���ĺ���F�S�L��wߍ�n����*!�2���G}4�9��Z3{,����nX;t���ܕ���H/��E-�"����(�r��m98��=]��}�P%��=����j;`��q��Qb���+тU4�	�Ġ�����Yg��=��7�|3�.]
B!��*++q���c�̙���h��#�ˮ��	T���0-s���hjWTF��R�ҊTY#ׅl.CW?E*B"e��K"��U��O���>���6!�̙>�=����\� �B!��^Z
�\�~����^(�{���}�xMVZ���[�&w��X3�fPVqq1�����X�`:;;A!���GEE�T;<蠃bZ;Lֺb�s�5C��a4����v���ٚ�ݡ��.��-�����wB���0�r{�q��{�_����	+��W,Q�\�B�`�� �b���B�'�y�n��nx������駟��!���L�>]�&N�U�v;Y*�}�2�k����M�VZ��4"UzF�����NB"gI������㯧�(��>']�7|��
$����=m&�8P�zp�}��B!�2zx�5s�ƣ�s��ܮ0����X(T`T3L�������]��5C�c�r�a�a��ɸ�����G��B!$y�6m�ϟ������
C96�u�X�ۥE���v����uC��^���\PZ��Z��OH2C�;!1`�	�km1fV���G�/�+T)�X����*�ocf�G�S������c�:��c�mk�*,,���G��^��[�r�JB!$���˓:�s�1��Ȱ� ���3��}�JqJ�O+LE��ndl�jlצ/�jd���q�`Ֆ!B���O�+���K
r�ܵ'��;^�+�Ǖ>&:�`�v��c�������7�kA!�B=S�Km����R�vuxJ&5Cy[�n�ً4hǇ���j���c�ӊ���|�7����a��X�������^����B!�$/999�7o�Ν;*j�v�#�����I�0Ts������
Z7T���v��_R�۲��9��wBb��A7��4�Ǻ�P�LK�dT7�"�,�!-��[�*^�����V�w�����m���.���kLf �B���w�]t���#�Bݎձv��ܮL_���]ܺBk)��t��SjK�C�&��	��L�Y��x`��{0���U��8�������`8��vB!�BF7���++�pX�}[��w�ݍ�v�Pt��j���]6��ռf(�21����a,��233� ��~�M7��o�!�B���v�MJm�v�mm[;L��b��v���$��d�}��ڡCSK,(��F>/8��#D�Đ��a|�^���y�,�7Y��w;�E�V���pe�� ��#������X+ǆ;��]VV�k����n��6ttt�B!�E��;�8)}A�0�E���X;�S����|��~k�H���FwS�J�4�b�M����j��	�%�L�"Q����BmE	������q����/���w�3Cs;!�B!��������م����0�#-GM����]��#�� �k���j���~{<��x���裏J�!�B쏨��8��3�^;�C�0�������bn׆c�kn���i�s���ݡ4�k�?���5Et��Ę����6�;�Y!�aIh��>㻩@�<"z�L�i�Ie0�L�
g_�Ɔ3W�m�|���i��p��7��?!�B��;�/�S�L���=�m;Tf�B�<�06�{����V��C���v�oh�`f�֦��,N��4��,H�����/�K
��{^��]�X�矾�8L�)3Cs;!�B!�E������\����4�wS]%`��j���&w1Ә &w�z��#��ŲF���8�!�G�4���B!ľ�/����ԩS��Vʱv٧W/�ܮ�!Z7�;+���`,Q;����[�Ǣ�As;!F��NHh�4���ZԻ���a/V�H�0��&�����oe"�L�`�}���2�A�]SS�;�o����N��B!6!++KJm?�3���7*�P�&B��M_���e�{l��C�"�6�AޖƔ4��e4�O��]����c���SP_5KWm��g�*����ڇ9W>�!�B!$u��v�+��T�Hj�!!j�����Տh�1ɺ��13�ۥfm�z�k����v��<���<��s��E!�� R��Ν����7(((`�0����~��e���ˊ��}H�خ���&�k�۳���QW9�\ �C�;!q�N�V7����s��:-- W!�bUzz��T$�`ev>�}��g�H�3220k�,L�<Y2���� �BH��y������첋�Z��H沫xejn"R�-A*�K�خ4�MmW
U^�*��o�R�"$��Ի#�n̟;�p��;�IK���ڇ�hn'IBq~n��,�+ʕ���߉z�B!��TCt�:c�f���Y�ñ�V�UIT־$s�%����)w~�l��n�brW>�x��Ý�h����\r	���~��X�t)!��x����?�{ｷ�m�z$s٩vhnn��:?���±�en7Km׮�I�%�㱮�	B�94�G�\=��k1�w�Ȗ��n0�g��j�{@���T��+�9ceV���e��Xm�����nÿ��/)�}Æ �BH������ܨ
J�n���x�W���ւZ����n&R��۝f� �J���P�7�d���	I$���=����/��}�O��v~�#��(/��Lm� mO�҈Ң<\p�+ �����z��uk���z9���bD�f'�+jј�L�$�:���:nD���]�UuC�P����a���ѬZ�?Z��k���4�|���$}�B!�G���t�I8����l;Y��f���v��a@�P'+Z�v���]el�C�4�Cq�?f�i��Ųͼ�#�
4�g>]������1�K�V��so�T�(	V�ڧ|N�������x�t�A�2e
,X ����@!���"�E���?;찃nA�.T4粋@e����nfl7��(�7�;u�z�vS��'T9�UV��[x�F���ɝ�v�l��f���2�����~sHj1fL�&��uM�3]x��)eI˚�=�¼l��Ǣbl!Č�7!}|��$-A �$a�
���$מ|5Ñ���
�Rv~V��S�5�h�#�&:�;}�t)���~ !�B�ǎ;�(�EQ`W�z$�ڥ���on�3��r����C&�v�C����%.�[�&�in'�*4�� >]���'6���u�M�k���n�{��d���9�y"�7s+���WUU�n�A���N��B!1"??��vN8�)�!��T���(P	��:�-�۵b��0���
�ܮ�^p�6��/.���;!L�'.?逸���v����$���љ�B+��U�c�%�b��@l�0�?}�q82A��Yx��ˤjB���vc�P�l����C���m�������Ё5C��D'�T�Z1�Gc[��z�!<���200 B!������c��g�a�����XϺ�|�cjn�t{V�����B���v��}(Hr����jk���1��n�梟b
�$�ڝ���&�nmS�K�ұ��D��L5����cx�5�<VE�p�鍵��$��b9���%����ƫ���:�B!���~����Css���h�b5֚@%�7���h�ܮ5���*M��+4s�R�����6��/.B��X��G�m<M�4��ddBY�*K@R����j{�����_/?G\�8z Į�+��?�?�^��X���q;oq~���8�m!$�Y7�1�0ah���bR+�خ�y����T�B�Ь�>�=�v^^~���Jz�m�݆o���B�.�=W��ϟ?;�3k�qاgnW�hn7����B�"2��u|����]X�� }��4��@�mwbFCе,`_D�n(4����z��4��x�O�%3�zY�J3^b�Oz�a��zl4�e��|����kp�Aa��駟@!���)--řg��#�<R��_"ŨH�cul<�P[��Q����>��us�J����ʪ�<��ؚx��in'��4g�$KZ�������~1�p̔��x��_c�Oah争�RR��g�>'��>��򘟯j\���ɍU ��p�z���(�o�/���ڵHV���]><X��^��\3�[Z{��v�	��?�q)ͽ���B����"��HnO�����d1��5��p,X�ۍ��ۅ�]�v�1�7b1�턄�$����p`c#�ٛ�n"R���Y����S,	VдT$3�Ee"C�+�cO�(��`���>�:u*�y�<������!�B�#�ifϞ-��+++��(�Ĭ���MZ�[[�d��А3ts�7�!�l<�o����d@��ǌIì�m�s���y?����$�nC�{��'��!{o���L�1��܀��������HH���i|Q^6�~���.�Z�X1u���c0����1'!D�竇�gu���I�[g͌�t�Nc��f�u���F(F&��5�P�srr$}sƌR����B	��*�S��ߡ�����C;�
C��ݳ�nh���Z0�lj���1��܊y7�7`���6  ��IDATJ��		�	�o�9q`c�yY��Mn���/���(���p�*X)�aUL��(e��v��Ǔ���SO=ӦMÝwމ�>��B	ΤI�$q��?���E&�����*n%N�
?}A��hrWR.���%s{i^l�
�RB�}X�܇�B	dJ�x��dmG7���ǘ?w��9�'�}�f��Ի $^���p�uO�ֳ���BK�df�K�g�#.y�u�������������X���޴�?�6!Dar߻�c�D��a:֊�*��Rw�����5C��i��%�fI�/�5�h_�)677�;��;�#�W�ZB!�X���g�q;�0_�h�
��v��rl4���E�kP7ԫj��c��C2��[o�pHeno�'4�4�b�js�WM�pt�nr���{Py�B�
K��)yd�B� �*.ES�J���HD-����&,X� �����ΰa�	!�=���p�	'��OFnnn�bS���`|�T�
7}!���#VI��+�@e��n`n/(����p��N!d ޶wj�I]D��c����b�q8f6m��#�}B��[_-����õ���3�X>��;7ཻ���}��]���A�:18�OR��;����d!#ã�]�(?Y#ۓ�����8?'�ǿ�eN�����!���j'~>�[[U�[�*�����_��������҇W3��q=Z5?���Hk�b������>������E!�c���q�QGa޼y())a�0
cC�*���Fv��ݻn�������B����wy]��Z؈OV��NH���N��X�:�Y�pl
4��IKzFt�[!PI�[�8k:�P^$�Ņ*�]$�h�B'n_"�|�|����Mʊ	>��V���>��C��^{�{��k��&]�B!�����q�9�H_���9�%@E2W,�+S�
��J�����skfpw5��cn��J�КIs;!��QC]�X�e��.'n��wp���t�u�,����� $^l����z	o/n�mgj�5+#}�����$�����<��	!���݉iuM��V�ܭ���[���ļV��SZ���x��Q���=ܹ�n;�r�h�q��a��������o�?��[_&�BR��N;I��=���w�vL$�ўst����c9M�������_҈���?!рwBl�k-Ø%%�/�8c1B+Z��+!TɷR�;4��(�<I�O���k�m��/�W^^����Gq.\�����BH*SSS��O?=얂V��i;Vǆ;�����v=�ʸ�ఁ�]ahw�'0	UJA*0��/���vB!A�p�tdg�_��-/I���/w�4r}��h�r�sk�噎K9���~#�ɀc���$ux����ﶵx����c}%����e����k1!$�_�Č�F���w�5!M}0�y٭^q�ӽM���\�>Ǻf+#{4k�����5��SC�u�]�$���z
�<�z{{A!������v�Ν����QW+�n'�̮��3����R�͍����4aX.}s��~�W3T������D�WTIA^ku��m^�C+R�tS|���`�� '2x��y�!b[\�$��K*��VE-�c�L��{��-�c�=FъBHʑ�����>Z2��*bT4戗y=���!Pi�ĭQ[���a�J_�
����t�핒��9B!IDiQ�8�@��d�t�Ʈ^\��[���왇�"&��(s�o~���KBCnv&��㑰W<�O<��g �CۚNr�#���Cp܁Sa7��l���<ZVw�B����.L�oDږ6�1�X�z�[9�ʷ�-����� i��U3�EM�i�B#=�Sp��/�^}�UB!�Jzz::� �u�Y���N��a����)f�C�����v�`��n�N�+h(����Q҄win'$���N�M�g�0f6�����4�P+�?=���`��Ifٖ�ޡJb��>+���1�����f��/�9�h5{�l�ﾒ���g��.�!����~�퇳�>�m���mw�)���"PYI_0n-8���-]��А~{� s�V���/�Z��r��&�b'2������b�mk�:�r\θ�Y��؅)M�q܁�5�ۍ�N< �}�#Vo��:����~�g9n��,��d&�!I���9�}�͑�.BH$��܅i�M�71���z>m��������w�C2�ۨfI]/Qi�Ѫ)Z����W\q<�@<���X�d	!��TA�N�<Y��瞾��c̶�9�N۱:��<�ui`8��vhP7�3�w}4��&vC��Y(�^ ��V��-n�4�uhp'����m66 �����d-�|ӗo�+�j�J9��p�Lc𥹏,�ANfHK��1e"�Z�R>�h�R���!y��1eee�?>9�,X� _~�e�/HB!�Iss3�͛�3f��9db!FEc;
RᎵ$PE��hpv���AD*3s�Y{���	x�%��vBIB�L���]p�϶���4���- ����}�sI���de��?����z<��XҲ�=�E�z)�7����/���U�_���j�P�#L�:#�7n�,��B��ʺ�\3T��#15�h�c]#�G�����>�}����s��G��͛A!��fJKK�n&�s233cR���^;T��=�r�PYC��ܽ�C�]���X�Z�+�vh�e��Y��]؄�2JH,�����V���؈�nu*���^m��R�2�<�-����9���4�4i[�#0�A����(M�z�&�h��c!Z	v�a�w�}X�h��^�]��B�h 77W�N<�Di}4�Q�n��Xk���/��4��i/�W:/��������eG<GQ~�s-�ƂRϟKJ�t�&�����f��NGq~N��->�<��q�����~BH��d���n���e����!�A�
���V��W<�B�N�\�j��ܢf<��>5C���QS4#:@w�q�9s��������B!����̚5���oQYYV�ʘdގ�X�$�-_�PZ�=!����F&wW`�˿m�ܮ��,��Z؀�V��NH�����$��v�dr��n�nsI�ֻW7���V�U���P%3xE+��HwW]̈T �/���}E�dH^G�J�G����x�	<��3���!�������?��v����&N�s�]�H��*P	�#������ghw�TA*=�ʻ�SV����BI���q᱿��غ�o~��؅��M�A�|��J���5��C�|�����9t/�t�n(/ɏ��C.������ŏ��KB�%��vb���/��
xA2�u��B�;@�	�3������4w��X#���h�>�7F� }��K�/^̀B!��)S�ଳ��ԩS��x���1G��
���@� s�b1Jm�^7�1����������m�U�#����NHL����$A�ܧ�5!ߛ� V)D#��s�VhVn�v�/R��*�1I!RAn;�Hpcx�G���i��M,E�pE�P�H��>�p��S\\�s�=�gϖ�^y��"�BIv�m7)uA�
���l�]ŭh
TJ��5��/L	�H)X�)�P�Jb��`(R9�SZ�in'���g��.�Ӹ���AIAnHǮٴg��<z �.\��h�.��Ղxx�#�ɘ�HQ���w��BF��rb��zT,Ð�O�kfD�o|uBU����@s�R��#5�H�|��&´NQo�N;�x ���*z�!�^��BH2��Ѐ3�8t���h����u��.�B��*�jr�P�~hT7ԫw}���v|V��j�rJ��~(n�n�f5`�j��	�54��D��}j�P���i=(��b�Y��R�
8�/V�}ij}������E+9�Ay>Y�2�����F[�B(�U]]���Jv�ax�G�t�h����X�8NN�Z+�D۫D!R�E��D�ȟ��s��>�?�g���.H��^�[<�D��'���D���}����.ĩN8�P�����1v5��{l$U4��"���]���/([��ܲ:��Bs;!ɀxI:��=���
t��し?�Ʈ^ؙ}v��#��$��>�޿��w� �E$;��ۅ d4�����=��+A0r8����#A�!�W�\��.�1��L�/$��@k���U�T$����C�Z[3��ӭ�i�~�0���h��beZ�U�v[�9c�<��x��'���B!$(,,����O<���q3��sL*��A±t��w���p,�Sܧ���'Z���4���n�0�f5b�Z��	�4��d|�r��6����w�_o��֭	Vj�J��{.$�b�����a0mME�4��D�`�|���B���m��3��1����.���R:�ʕ+�bJ���M�D ��x��盨�gee%�܂D�����D�_�����^��s��߼x�~��|s<1��x<���RI��3g���X�SV�$Z�J�\���*�G�֤��/(�*�"���@edr�(��[@In�7'��o���w�}Y��̎%9���_a��ɐ_R�0�����r)H�Ѻ��7n�[��ɍU ����u�7�kA!�����C�j@�s����EY7���U��݊���f���*g�X3�GGҫ��i�Q3�R�-AXVj�� xꩧ����L�-���+jW�$�痃�䰚x��?{�3?�D���'����Z<w��E<���{A�~����u;���ӭ�wF�T��?�C9'�t���,����G�/s$c�P��Hh�����6�{n����Pp�{��ݻ.X�Ո��NHܠ���$D��w߄	C�U�ҍbݳjlt�]D�/VYi=��If�"8Q� ;D+�,\)��^��+J�A�Jt��1Vƈ��������^���7oF$����d"H��X�|ip�/�evM��^~�I�}"����a*~�@	����>��g/��"=H�,//��8eeL�ŧXoG��`���=4�J-N	ûn��N{AS��������ڒ��:;7�W���yٸ��_a��-�������p�/&���L����)�u��}�#����2|x�� �B!��uC��G��ro��[U+T�b���
��|G�w����Y�P�'��=�v1:>5C�eY}<��a���Ə��.��f����ߏ�?�8j�����v]K��e����)�$U�"�Yև��g�= �ά�w�&K#�F9L� !� Eƀ ��c��:,go���y��ߵ�������%$`�D"#,��Q�a$MN=�߼��vWUߪ�U]�]=s��ݷ�	i��3���|����y�ݞ�����y�3���gϐ���>������_,������Ax|:sƲw�tΘG�b1�#4y�#��nޡ�34�cY���;>�y�v�v~ΟG[im@�����; 
ou20u.5%v$+y�A�"�X�Tҝ�m��9)R�����u�,�m��73�w)Zeb�xNX���)̦� (AJg	�-[F�\r	��������^   cٺp�m�QSS�˕8�3'j�V.�e��!P�50��w��v�H�s�&4ӳ���C"  ���K\��'��|Lrc�u�vSTش��:{���     ��~� ��ϡ��v	�C`	�'�&Gf��ͻ?'���=y����A����y]x�a�`����Us.\(v�~���?��?hÆ   ��w�!��}��������w�;�xoi����^}C�b��w�����v>JJK��,z� �� ��9|  m����I�����ɭP� ������1yS!�'+�Pb�z0-TY�i�j�AtO#�*"�؊0w�����k����ٮq�4i}��n����>tO��   @��}�٢u�N��D~�E]�
��_�*mp�T�w}�*njl�cj�h_07/�ĩ�p�lo7T|���fzak�v�   0����I�vPT��o����_�B     �0hm��������V脡��%���td'���I��ŗg���I{�|}����u6��WO0�׺��5����Yg�E��v=�������v��E   @.ijj��~����}H�d��5��^�]��:����ڵ�����w|v�+v|��>�+��׻���vx� ��(p6�Q���tZ�>�7ni$+rnb0�d$�96��P%5�D�}�A	�ԸݭM�i�J^'W"T.�������|={�l��W�B�^{���x�	q�   	�9�S�8�x��y����Zwl,�߃Z�j]V�r��4�+�TT�D�T5��!P  �-��������"�    Phl;����t�����c��(n'�&��ٲ'��a%y� <C�.�#���ǌZaP�aО`<�0甕����_OW\q=���b�{�   &t��7Ӳe˨��"0_0�9Q�ú��;�� ��o���<CS1������v|������}
��w@�@��Q���!�M���ۨ��;%X%��av��!Zɛ�&��@��"��L
W��Ny���=����+�����R���wz����sM�st�͟?�����n��F��/~A�>��B�   �s���-��B�^z��g��8�gM�_;�˵@e�䶂CC���N������-%ʹ~v�  �{^۰���Koo#     Px���g�&�ES�Po��.A6���)�n��M����̕����9:�Q�UUU	�pɒ%��ϰ���   � ?~<�p����|�&L��w��n�{�����af!�|��o��cs{�;4z��r�ʚZzz�D:܋�O �	� �t���d����1V)�Jf7�&�*�,����0r��̐le0�K�DU�7!B�*2l=(E+qXW��������.�慠)]��N��~���v�Z��L���
   ~�3g��_s�5TZZ�wqJgN�Z�s��vkc;#�(�@��w�*0�jD�ri_�in磤��6΢�n  ������{;�o F�     �{��؞	t���j?dnq���v^��1lϐ�BR�M�!?����F�#�u�=�:�aÏ}�ct�W����/���   ������.]*v|�2e�oP5�+��Ϛ(z������z����_�{�v��q�o8��n	���]��k�O�G��Rw�  � ��#�CB��|V1u9l�SJ�J>U50XĪ���!-z��B���Zd3C�փ2�n�I�*�<�>�G)X?�lD"���l_�~|~��w��{ٍ�|�������{�9��OJ6l���   @&�u�������@5nܸ��t��:��c���N���!���d�}H��])R�)���Jz�s*���ւ   ���Z�yE���!��7ѥ�M     ���HЃ;�i���>|`���4�[��v�aJ)@��f^�������x�f��J����/H�/�{��v���ɓ鮻�%&����C��	   ��7����3g�1?���XT��^��*�
���C��v�b,�ops{��zzh[5�ǐy 
 ��(CV�j��R�j۟��V�
2���Sc�g��'�V����I�����dн(��`k�OZ�J�v���֚0��q����O/��"��g?�u��!�   ��1{�l�馛��k�����@�(�X!X������}����a7���ڕ������z�P=�F�  @nx�͍t�9Ǚƾ}�s�o��u��t��TY^�{o�j�@# ��8oQ3͙RGQb�C�f�V �0���RA�4O�����&w2��Dꂬ�3�w�Щ�]��m(V5�g�ce���Rϗ��u����0�����вe�D��w�����    '�/������[o���F1���w�Cw��z�hl���5�����lo��<�V���PT[ � �0
J��M�tM��n�m
��T%�Pe|�jeQ�L�r��$�M����:螺�H��i�A���U���pu�Ma�v�x���y���:��9�C�/���~�󟋠;   �_#�ΝK7�|�خ��l�Y��5�
Pn������@e#N�TZ��#�P,��j^�k_0	S���	u������?D   @���V�c��c���������HQ孍������+7PmU9m�w�n�?��vw0�9�q*M�PM;��-{Qԩ_E���{�W6l�� H>����'ŷcye�s�p �X|�sΦ2�z�,�;�CY�e���X�q7�0l'��ar�������E�]��q�b7�c9{�E�|�a>��r�!z��ͺ��&���{EPq���j�*4�  Ȁ��%K��-��B---b,߾`PsF�wh�����s�oh��5�C'��T��볭wh�۳�p{�,Z�ZL�� D���]�ZJ�7�۶'GD*�p�jb�he0�V	�h%稄��he�g44(�����71�д�w(���Vˏ]�ȁ�����f������;�<Z�f�򗿤�k�  ��	�o��F�=m.��\�S~�D��^P<3���sq�8�"LǍ�v{��lO70��TN��,P�Ll���WR�  �c�b�ﮠ{Z+��쥨���ʹ����մ�`;�	�n��t���.����{�8���7���u��S�`-��>@_��TWS!ƞ|�}��?�W�Г��b���3	  �:�Y������H�m��~��K�Р�94�{����ӵ�G�;4x�F���Xv���K�Я��տ+������P�j�������u�]G��կ��#   ��B.��b���F1��`�ε�~��wh�[�錾��;��u�۝��<ϩ��*Z��|��&Z�Z Qw F9��]��Ltds�&�(S�R�V��ɌS�h�67����i�J�I����U
s#CR�J�ܓcىPQ��%Z鼷�:�1>�>�l�����/ӏ�c��nC  �ZX��馛�ꫯ[�#خ�J�=�kxy�tNjw�┎@e�[��*_[*Ī��3iek)�  �7�KО�N*$�z�F?��L_���Th������T���������ڻ�(J�������7�]���诮]L���c�;���6   �Yݚ�����l�}CRܭ�!ix�:�?z�1�^�lpWy�EER�J�9cY_g�	F�S�:ǯ���8o�<�������鷿�-�X���  0����GߛP�=@��F�Wh}���˱����ή�z�X����/�-�R��|�&z�;VUp`����9���{���@f+CJp"��A�2��^Z����ײ����V�sqV�J�L���32��GΊ�وJ~B���^�/�k�9'�1>�:�,:��3E����^z�   �>�s��hٲeB�*---�`{Ps��:}&^�
��"N��)՘]��N�J��kn-�jl7�/�7��/ �    �b��zR��Ҭ�	4i|U���6NQ�7M�D`lû �  j��2Dg�n�����34�ۍ�!Q�6d|n
�+<Ñ+����*�X���<��3$ˎ�F���'�+O��5��	r��؜9s�_�"]������GA�  � ����[n_�(��~׍f��)Ԟ<���y����\|Cǀ�����%�����fzc�  �� �^���6SmA��Dj���<%@����S[�O+�w��aE\sD��&�p��z�~��ԫ"u3C�!� '?"QP�R�B�1t��O�=����裏&o   4�9���N�k����;�<�<*�v�X���A\#8��x�'���s7qJG�rk^H���*׭!w�n��fz�5F      ���go8�>q�  ��Wv��MtL�.�����к�gH��a"Q�k�g#�/,J��l��EZ��]���#�u�=h0bcc#}��_��n��~��ϰ���   �.jkki�ҥ�kƌbl4��:s��Z_;y��\��7�;?���*��Z�e���ȣ]���7䣤����E��BN	����; c���ґ�YtZ�~���5܍7qJ�:�$yc�z0}SSb�ҍd�~FJ�ۇojR�U����|�%�+y�ea��γ}m}��~�����ur=v�	'����Z�z5-_��zzz  @a������t�u��駟�2�������?A^+_��\�v
�[��T�J����ۍ"U`�B�b�U4��m�     0�Yz�B��_@   �y�@���f�i5���������#�x�5�=C�|�ݟ3�C�Gv}&C؝�B�%ړ�s��)f�����
cl֬Y�/|�>�я��;��$   �͔)S��o�����&MJ��`��u��;T�3�C�o�j�R���-�X�;>;�+*+�厩���! � � �1v����xZ;uwq��Ū��e��ܭaw�ΐ�TXE�l�g���� ��a��r�|�555�=��C7�|3=��Ct�����Ç	  @�)//�+������Z:��c�X6����B�G]�J�s�W����~�(NY����S����]C��mmW�Uee��nl6���      �v�m�J�v�U�qf��.���?���~�'���  @�Iz�S��iG���=p�34�cI_(��=��S�}���g����g��!:
�aT=�l�e;���@w�y��~�a��ر�   ���"�~�UWQUUUV�`�cA�mޡS�=y^�7t�݊���3��*�P{�gEȽ�v<=�"�E��Bw � G���Ȯ	t��R�:r�F�J���xe�S*�N)��T٭��f�V�I���i�A��nYEFK���������#X�R�]5�?�����b�
q�۷�   D�	&Q�n�:L.��|��s!Fe{k�]>f
T��q�0e��D)�9c�]%R%�)s��1�n'P�D*Ŗ�����*z�H��D�     ��NmU9���7PUE���/���y��   $a���i��q�uhr��7$����3���3�2����C�Zʱ�~�zh�&v�a.C����jkkEȝw}��'���w�y�   D��`�����˨��,R�v�X>��w(����*�����C��5}Cۀ�C1��� �Ll���WR_,N ��w �(��qz`K-m�I�m;m�t���|������	?;��,\��˸��5�.���f�$R�yUD��E�ǠE�\�XaΉ�X]]�q�t뭷�3�<C<� ���   �̜9S�Y��;��`�j,jV>-��faJ-R)�)�ւ:"�N�BR�ro_�����G��:zb�x��G#"      c���+�y�$�y�~�����   31�������Ӷ��3t
�KR���g�����Aw;�aw�_h��#��W?/�к��z�`��A�_��rQJ��������^˘   ���ŋ�ݞ�;�<*r�Z\H�v��F�wh*Ĳx�N��V����w}6��ߐ�Y�BU���;�p{U�lZ�ZBC�� ��@��1�P�H|�PK#ڪ����2%L�+kK�5�lq7^S��.�S����T�LR�"�6���D+�"��5�uL%2�r���%K�Х�^*�U�V��;ߠ  ���~:-]��.��@��-Dq�Ϛ0-'a*y^j��UN�v>�l�[
�k_��ZP!R�L�NnG�C�      ܶ��t��6�<H�ߏ   5�>�ZJW�k��6�gHd���8���-��7���z�V���g�hqWy���#�a���l�??����(�ڭa;�8����$�ׯ��+W�O<A}}}   ?TUU��_N�\s�hng����sN>����5���;T��nޡN1V,������n�n�a,6H����r��� � �M	:sv��n?��'��S�!�Zc��(X���N��aڂP�ߥY��7m����KA�Ma�ڝB�ټ��5��p%[�n��~�V�^M�ʘ   ���8����)��"����]��`�Μ\�Q��n�c�t�)�XR����3�4��{j_P�T|��~-oM�^      ����4��n��u^�@�>����7@   �y�5A��i���-40���<Ì��P<��X$�d!�9�.w�6����BU���3�B*�>Z<� �������ԧ>%B���oh���   7L�:U�q�u������X!�Uc��+��V{�f1n�u���q��^��?���]�q��;��ή�za
4(dp ^��c�4����;ykcp
��JK���%
��Ķ��vO�SE�-M��H�F^#H�)**�T��xcc#}�3���o�]��W�X!B�� @0444�UW]%�S��2w������U�Xe+LY���T"�5؞l_��T��*q�Q�2�T�D��k���VT   
�����Ʃ"l��{;	  �7�JK�??-U�s�����Oһ��   =����6S3�Hz��pWd|�η��l���ܭޡq��/d�*���'�n���D"rO�n{�WO.J�v?~�)S��[o�o���z�)���M���B  ���?\č��!VTT��Us�ձ���wh���<{�n��V1��o�۳�oh�K�JiSb6��}�  �� ��ҡ�t��6����Z�"�p���Y�R53$��m?(�*�-�t�!L�VA	LaP��r%<e�����n��f�馛��_��{LX,�  �n=��E�a
S^�FQ�ҙ�����I�J��)��v���8e����8e��l�)�p��H�Uk|.�y;��   
�������A�3&�����3��/   }n[r
-l��:��76�O�:  ���}�tx�L:}����I{~�9N�k�Y��靟e���oh�Sa��P�ݓX�B3~<à<E?��Y��:Q�2��lִ9t��믋b��~!  ��q���/�=�z�b�P}B�1x�f�P����!�Zۭ���?h����U�5��p=��D��� �  {;���މtUcu����lE+"�5f��i�A;�*%TY[��J���>��I�6ZR�
S�
S����uY�\�x�8>��O��O?M+W��;v   g&L�@K�,�q�'Ƽ�Mv�Q��$`}�0e0���m��*�����!�ւv�v-����^j�B�;n  P8����ޒ
�3��i˞C�z�  �GC]��=m�t��"��  @���Ct�w2]>������Nޡ�7�ls�b��w(���Gq<.�T9��7Lb���~<�|�ؽ�w���-�q>N;�4q�ٳ��x�	Z�j�B  ���3�Ȼ=�s�v�uQ����LQu�����C�b,�p{zh�2,7�06|���L�L��UM��C  � Ƞ?�����ʖ94pp��V���`e�KLAw���20f�*-V%��Fa+��z�D+�s�\�6�w���Κ5���/��n��z饗D�}͚5�&  @�c�9Fl!�����Z1�Ka���(�S:s������Eu�=S�r�V�)Ԯ�gn-��������^[WO���~��  j*�9S2Ư9�8�  @��	�����C=  �?]qz`s]�2�znOjM���k1i�0����[܍c�~!#�B5~<�0<E�9^��(����O�N��v�������W^y~!  8PZZJg�u���.���21�����Q��|y�V��8�W�e��y;�0�p{U�,Z�ZJC	��; @၀; @I"QD�[�>��B�G�؋O��͏b,� �s�`e�~�M�������)�ȩ�A"����:S!���&�bQ>�'��ݮ��l�{��ضm=�����Sww7 �X�ۮyA��~��b,�n<�"V��)?k�U�0e��[
f�U6��q��������F06"R��)�Hen�BԠ]�}D�z@Tq   
���U����$   ��������J   �g(QD�Z�.in�����mX]q������r#���\�%���B��;���.?^��:�zN��t�]cܸqt�E�c����/|�G���   �ĉE)MMMbl,���c�
�g{m��a�g�P�w��s�o��}�ۥ��RbR��'�^ &� yjs�N��Ds����xK���<4�,u��x�$�`E���lg�؉V2�.Ī�J-T�E���E�ms�2'�u~�������s�ҧ?�i���?N�>�,=��S��/���  0��υ��~饗
a���.5n7_w|4�X�d����B�,C���P�U����Z۝�\[��T�*R���,tQ=*   ���	������4i|��   w��XC   �����贙-4�k�3��z9�^a���K��n��_h���8l��{~.�5+|.�к1�9Qs���������|���Nz�'D1�믿.tO  k��R.���~�������?/׈�X���(x��1c1V����ש��v�B,�%���Ụ��	 0:A� �ʺ=1:2q}�z���P*��pã����JK3�d����`'Z��܇�;v/2������z�7�:�S�!���B��������E���;v���{z��h˖-�  �Δ)S�K.��8��!4y����KQ+�k8	S��N[
�(�P�s��lav�m���#���)o�77�   (d�j*m�-�;�֬�J   �cp�{�8�>  ��vRӤ���r/����>����>�C���'hW�%}C�?(��I0��d%���3$�5��������;������A�׽\�����.]*���Vv���~G{��!  ����3fВ%K��.?�#���g;�+�P5^a���F�ޡͮ�:�X:�X;>��~�r�gKН�9��o:m:�p; �� Zl;����lvuڟb��˛���2׹���d�����*PYǄXemf��������@U�U�!�0�|�ڽ�QAW:�gϦ;n��vZ�~������A  P���Wn[��+�.�ն�xԃ�(	XN�HR���{5'aJ�C�vBU��v��{EU��5�v�G�  @�3������Ʃ�    �ȳ�P�ګ���tPg����d������N~�[����Tv7�c�1�1r؝�,Y
Y���vS�m�ٮ�2Gw�Ϻl�7��:�����'>�	Z�f��
��y���#  -p���Σ�.���>�l�'2��f�>�~b.�����C9�����<�ۭ;@�c����S{k�p/�C F;� ���ӊ��te�l��,8��W� ��Y�<�I
T雰�p%�(5�N�b�0ejrigP7��U��]���u6k���y�\�97�q~<��q�]wѓO>)ī��zK�4 @���c,��/�X�-ps����t-��|�X����z�S�=}^ue��n��`��ĩt�=f��ۥX�p���J�l����!   FU�e��o�N      �z����j����znW������]����m��r,�]�=�/�mr7{�d)ʒב�e/4���{{}P����'G����z�~�a���,�� @�a��k��ɩq���/��;�C�B,Sk��7t�[��:����3i��R��k4 c� ����V��9���{������F�op4*���&*砻Q�RWv�r,�����vc3C�HeE%Z!b=G���՘����������Z�v������O�S�  �7����/��-Z$Ƃ
�5�`�j,J��k�Y��R"���$Ly����H��Ӑf�=%N)ĪXl�J��ҊM�qC�  0z()��1�㛧      ��P��V�]��L��[\u);���?4z��6�d�=��j�z�ZM�#�w+<5m�ks�cQ��|�^�r�>��'���_/�6�b,�<� i��شi�D�����Ɲք5�O���B��\#�:x��J���]�����w�
����l��=ao]3=ފR, �� |��5M�K'U�����͏!��'�nlp7
W���t�]�Π��Aw��3�U�v��@%���Gy��U�ʇ ��P��`�G���~��1��9s&�|�ʹl�2z�����_֖-[ ^ �F}}=�s�9"�~�g��B�Ϛl�%/׈�X��)�9VAʩyAi~��M�����TZ��ǘ!��=�n���5|�}Z[�<z�u����   �H���na�gM�ڪr���'      
�g�т�f:�tw�+C�r	�Km*���BØ�U����|B����0�r#hJ�S{����a���<���˧7�e��k�^�x��c��=��Co��&=��s���SGG�B @d��a�=ĳ�>[|-e��5��`|Pa����Q���X�R,��c���J?�l\��g��[	 0�@� ��-�c��g2]1��:H��(��q����Z%%z!w;�J�7~F�ʮ�A#O5�J��9�\�k���ݵ��裏���.��~�iq:t�t�{��Ӹ=f.�luuu�Ķq��Q��?s��(���F���|�ٳx¿�|mߙ��;������������O�o�*_a�׃/İ{P��䣝H�y���v��v�@5����@e��.���*Z�;�6�@  `t��7`{�����>��{�]     ��x�@��UM����Sw���F%�C�;?'�ڗ[�]b�	�x�~���&�>���\�e�Kyi�%��.���������;�T�=�����g��uz>��nz��W�g����z������ �.���"����̻�3Q��S�Z���;��z�r<��w(��Cc��T�e��<��3<C�)��'�s&ҁnx� �Ep dEw��\EW�̢����7G�J��~�C63��gW�b�*��t7�U���
T4r6�6w�5^��W>ǂ��͸�5���x���O�^~�ez���u��aG��^�����G��?����
l���@���5&_���������H}S�/��{�s,,����Z�?���Yg�E^xa�$����)*�|�q
���;4/$��n�v�p���=����IS�U�5���   @�t�8o��OO��H��j     �z�j[-]�\C�������n1V���*Ŋ��ܝB��]�����5׵��B�ϊ�ڝ�#$E��|�����P{�A� ���]�iMUU�(�������z͚5�7d�T�竜)�A�~�3�?�|�3���U����Οk�j1Vex|�N8A4�_|�Ţ��ɧ8�<�\��������X�;>�l<CyTO�In.��8�R �*� �fh�&���bZ<��&�lARS+C�x���7X�6w'���8���t�D���e���Tm�f�ʊ�+��8�m=ʂT>��l�u������#_�җh�ڵB�⦆ݻw  x���8��y%ۦ�s���0��X.,�%�e�T^[۝�)�p{����оP9y��T<|_�q   ��:�r��)�w������	     �B#'Z�ZD�47S���~�g��j<�*�A�r,�������^�v���3����:?c~�������:��p�>�!q�ݻ��{�9Q����;����)���D����a���;��r*��LA��ۛ��;��?{��>����$dS{CC���a�<�B��TF��?��;{�<G`��ҥX�ޡ�g����5���0�A� k����sia�^���$������p|���$b��4�����I��4��a'X���w�-�XP��(����
N�B��@�t�E(�-�]w�Eo���hk���@;w�$  ����^����nk��&hQ�������cVa�(X�ϻ4/$���*�慴Penmw�L��������k[���9� !  dä�U5��W�8��:�W�AX���Y�J      "��<D�4����"L��z��9nis����_�|m��|n*�2�m��G9�o�=L0j��h��O�N˖-������W_aw���3 �0�P��'�L�w��O�:U���#��&����B�{�}���&c�`��R���+<C�+����f�IooŎ�  � ����)�BKf�Pס�����A������,Z�O�f�3�-�w'�*����@2�>��n
���X�*3��t��1��~��;��~�ɟ�惷%\�n���ք� ����?O,^�8���P��5a�[A[Q��E(�,C�r:T[;;�S:�vlE�240TU��+�� * @�|��K����V>�v�?�=������8���dO[���8���v�*����t�gD���     �"���5���ɇ���H�+4iZ���ӥX��{�d�Wt����N^a��,��������_��l�u����9�^y��8|������A�= ]xw��;�Ǻ�:1�0��(�Uc�����=T���P�4�b���w����G��I������� �w @�t��i��
������l��,��U�=����.�IQ*y#�����Nb�Q�2�U�Fw�6�4a�V:׉�Xs��?.Z�H��smٲE�����khk `�_W�9���Ρ��N:)��'���ӹB��Y��u���A�.���J�R�S���N��T�v?���=C��<��:��b�  �����64\VZB?��5�PWC?Z�
勪�2��/^�nw����ᯩ��'�{w/u�7yB5��篥��%ű�	     (L�uѪ��tes���4k]
�0ᢁ��ܭ-�	�Prw
��С͝F��$��}�{�s�c�����xPk��'M�DW]u�8:;;EН��_y�:x�r- `l�;=s����N����Z1���������Y�K����\���s�c�����z��:�v�p��7Lۇ���Xv>��nϩs�AW?��D4��  Hp ���7�i�&:�t7��o�4�����%螾Y��G��C�NbU�1�>����^T�׋�h�� �5��sMMM���멽�]���x��h�޽� ETUU	1�SN���ٳS���ӝ��S�
K�ʅ�%q�\�t��	T���t�=)B9�Ucn߳Ml��C  A��@;]������V�X[�q������/��S�D�8���o��~�w���cf��yfm+}��W����::oQ]{�q���H_��<����#      
�X�hUk1-��L�z�S����_h�o)K�F��3wv
���B��Z���Q���6w�o�v�r�����_�ܰƃ^c=?~�x������Z�[o�Eo��(�z���0�������;<��Sš�ӳ����ڽ�G)خ˕�h�/�2<D]�0p��l�Z����Q<|_v���^iE)  � ���FM��#m�&v�f'�*�6W���������GnO���*�`e���n���hejN�Ƃ��x>��b^x�8>���Ѻu����_ֻ�+�� 
)H�y�"�Ώ�snk��/�*j"V���U���ۍ�Jv���bU��M������������;�Z� � ������k��;s�N�����]E����N�H�����2��v��o��os�1����|�N�?���Or���ϡ����H      2k��h��9t��6���P��R�~n��sFx+tO$��ݟ�~�])�|�� c}-�B�6w/^�D��F�-~aP^��<�Z�(��O}�S�m�6Z�v-���˴f���(�������>��o��3Π���>��:�+�p4�ݳ��S��m�g�`{Bx��p��wK���`���V�UYSK�v������ jp �N[O��o��+Z�i�m[��ʦ�����xOV#��F,}Cg���Tb��R��8�-f����읂��T��_�)(�*�k�\���������M-b���'?I������녀�s�N�z @~�mO:�$:�䓅0�`��@)��$X����`���5Ԯ�|T�ܩqA
SI�*�nn��SB���o-�
��s5�]U�яp;  \tB�W����>���u����4&���h�j�9O�m��!�>����O|�z�[�SYi��<�~��k��/�7m�{�      (dvw���:������2���XV��i�紦��W����X	C9����F��X�%B��0}�j���zr�`�B�^<�(��Aڭ���y~lllǵ�^K���"��ꫯ�cϞ=�
(��3��,wz�R,޽�x�i�۵�<��UO��D�0{����+���+4�=�T���z�LZ����� �A� ��"z���3����v0�M�6��6���4�`�lv����N!��V'��]�2�V�`D+�X����B��r-D��g�vڴit�e�����Ɔ?����/P{{; r��F9��cE���N���]�q���s٬3��x�D�0�)��$R)����TV�ʮy!S�J�S1�s�F�*����� PRI}#-oM��  p�����%��G���Y�5�#߼��������|��v4���Rey�����6�6�������]�8����~�՛�/��:C��      ¦?��K���f*��F���T���چ�-~aiJKK��l�:����Z��C�(}� ݥ���F)���ot��;������z��Z�^r�%��y���b7h>x7莎���o���Zb���X�w�)������F=خ˥w�
���ܼC�p��w��	:��v�_��B����! �� 9�]��{�lZ\�F]���6C��I�rmf�d;��Xelg�[�����G�ж �㪱 �\	Oa	Wٌ�Fu��Z����ؘnl�y뭷��7��wny��G��0�1Gu���?�xѴ0a��0)��A�R~��R��27jaw��$�D*�}�O��^�����TR���n-�$T95��ظ�2�V�H�[	  r��[�C�G�i�Ǿ}����ц��}��$�Χ�����n̏V�Bg;�.;��y�gM��߽����rq�      @����!j��H�*�QoOOJ��BU1�S�=c��%��~�gy���·�$+	?&�K���Q��	����͸���u��y~�?�8���z�����;"��~!7��+ w��0K����X�>��w�P�jf��J���;T�ٝ�C�b���;4������>bEe��J�A 聀;  ����v�ч�k�����U���VN�����[R�R�3X�4ދ�ܭ�u� Lb'V�q
�) u��ׇ5���ds��Z��������O�tg!K�{zz ��w�_[,X@'�x"-\��-ZDS�L1�ѹNX�s%Xy�VX�V�D�`���WW���0
U:���im��V�*B9�/8�c�T3����SC�{n �����I���}�r��o����� �_����]�� =�������q��-�7~�     0�t(F��hɬ�lۧU��S��\#}��a�����0����������?�ҬD�����w�=Ho�mn��:�ֹlϏ7Nj����[������+�П��g����{B� m9��E;;�b�z�TWW�:�?�v>��aB�Q�[ǒ��o����om7z��z�N;>�Q[?��QA](| x w @^JЪ���-4sh�h��ݭ���X��i3�3E+�6wsC�J��υ`���he�E+�^��^ǂ�r�>�qݏ'�s^��9o��m��{�8���>v�����oБ#G �	��ܮ��v�N9�jhhH�"Ю3'���ӹ(S^�FU�"�[
�*�p�}k{�,L�B��ւvq�V�y����&Z�iH܋ @��	���ہ����w��|��W�;ν���i۾���O�E      �:��|S]��L��[3�Es�
嘲��R����7�osOͱ��y�c��w	?U�?&d@^��q\5� {���B������4i]v�e�`<H6lHy�z����_: @
��͛��a�0<�(��a��a]#*c:ޡ|t��!v;���ώ��P{Vޡ�3��"�_��&Z�ʾ!�C �7p �7v�h[�L�`Jui������Ūx�/v���������U���t�J�݋��p����习��̩��?9��?8­�7n�w�}W�X;v쀈��'����������4G�Z�:U�*
!�(�S��,N97/�m+����.NŅ�}����A��
VUц�i�n+��{�� �0�R���77�Ǿ�[��A����?XM?���2�7��rj��F���� ��~   ����-C�2��U���n۠�]���X´t<���p��۷��s'�P�ڶ�����K���9�����1��~��;��:�����B��X�4ݹ �=C.� ��?hg�����C<�3����\'�9�����c<�>���;��B��s��=�y�	G�P�3b�,~�7�P����#��;|�o*�ߊ�v �?p ��C�|k-i��ءm��vyC6�XVVf+V%_������ܓ�U�A�*6�uC�P��h�$S���$Z���B��>��1��s^�5���\�D9r�޽{E�}ӦMb�µk׊�w���h����	nV�����:��ϟ/�k�q�������~<�"�~�]�j+R��m���F�Jݼ`mn7�T:�
�]k��
N�N��^N��  Q$
!w�ہ�����o�@_\v��qe%�󿽉.��Oh��C@.��'/��xǁ(p畧��s    ��M�b�����h�@=vfcY�2�`��?LXK�F|Ä�3T�b�}Cݐ;?:��<|��i$=D�G��̧����|��s����9��Yg�%���W���rA�cmݺ>!3�3f�@;{��%.Z�����Lst�����?��'�͘��wȸ�����q��[۝��=x��b,CȽf�tzt[�"� �� �H�H�c�q:~j3�+�E�}��m�f�k[�ʦ����`���n��vB�HXnr����c2+�/�t ^���8�����^G~�>}�t����c�"�Y,d�����5�+��*477�;�*��p�B����(���DA��&a��ܨ�Svw7�ʋ@�l��1�P�Y�r��乢�"��B���|�  D�|��n�|�7���&�ҳ:��ÿ��e����)��# ��o��p<��f������:z(_p���n������m��8   
��X�Vn,�s����m4�~��k�p*�2y��R����&=���Z}ô?ȸ����������%c�G!�����5t��e���ds͠��ͱ���q7h^��X��G�m�z��E�B���s!�1�C'�|2͝;Wڛ��R���<��e;'�P���\����Gu���g�ޡ����;��ͭ��v�����<D�w8�G�S'��8 @6 � ������i�dv/u�kl��)�*���]���(XI!J�s�tD+��&Ib��|�ڽL~E'/�����:�y�9~�q8���������l�B�7o�;v��u�����!f��!E(�X��@;?�P{]]]�\�k5o�V���̍�8e��bT�Y�2ۍ��@�C�k�K�Bu�xz����mC� P8�#�p;��G|��WS��z:�i��\����7��_�_�Y�����H��k���;^y���3���Aˆ���c� ޽�w_MW�c� �y��z�    P���=F�&̡3�SW��b���_��&d)�˧�܍���oh�
U��/t��9y��1ae"�3A�~^����E��нNkt��g��|6s����,�:�����`���;���*�BY���� D��������(�S����z��s���X5�0W>�j<�P>�O�v�v7��/��=��l��ޡN{�kk{�Dz�`�9� � "Gg������M�Tܱ����f��rÖ�ق��<1"Z鵹;ݽ�ܭm�#��X%1��j�V���:�s^�g3'�y��բ�	��m�6����w�߾}�8@Pȿ�3g���|p��[ZZ���B9�˵���*w���
��G��a��0%���mE*�Pe��┍0elc��<��\D�8 ��C�ܗ�#4i|�ɓol�ۿ�p;�FOߠ���'��N��q�A�sNh�o}�
��& �e(���|�A��.�>w�DZ����-_���mړ������~�77�Y��Α��w"x   �v�Ѫ��ty�x8�ͶKu8�-d�]���cx�����KPU�e�j��l8�X�i/1��{>`X���|�lר�yY���9v�sهY�h�8$��c�ΝbWhnzokk�� �5'NeX��3�+r��w)0�7�;/�/��Q�úF�>cvޡ������;�ʰ��v����C�_��;7y.�ܔ���p @p � �,On��I���� �tv�������F��N�2�2�#���9�n݂�)��[����d��3E*+A�VA�97�q����9?烜���e.�d;���0�mooA�]�v��w��k~�o|� ��f͚�
��s>i��ɦ��|��j^�
V�
�{/�`���^�����N�]'�Ώ�!s[�J�r���i+A�0ŏ|��V�H��  2����?�ӎ��{Ć?g�����ϩ�w��;Bw~����[����>�O��v��~� ���{C]5=�n��{9=��5�iڤZ���?L���A�   ���D��o9N��B�b;D���b,���Z�&ݓ~���ݝB�����ih-];�%&�j3��{e;��sA��fN6�x�]ٌ-aM��A.ǒ!�7m�D}}}@�������T���#��C~��GM�h���	�Y���_3��# ��lwkm7���7�v�ͥ�Z�ћ�  n � �4��h{�$��i��ṑ�N��7��F���Ħ�At7
TR���
W��+����t�=
A���1�e��9����|�s��e;�_�Oǟ|���0���!�����~!l�s~<p� ��c�{2a��3g͞=[ls��]��?01i�$-�@�}������y<��v�/q�I�򶥠�0�(PY�t��s[�ʰ�`m�4zrW%�C� 0:xo�q U�_���u߳����u]L�7綾��J d�NȽ���~�w�����Q��'�
�c9f�n�9y���ہ�	���_���̫�ӏ}�   ���m��IM�ζ���T�a�3LX=ô�!v��{�7��C��;@�#�j#���lƃ^�v��Z��A�Q��2���б�!�����#�����^ܳ5ܼ>o�<��i�ܹ�G��bMM�i�W1b�sƊ�`�jL��T�Ct;����3?�",{�Щ���)j۵���S�]Ut�7F  � "��P�l-��ͣ����'�u��
U���V�DR����A�d;����V��*^Y,w�trnX�A�	z���{���y��~�s�ٺ}!���:tHY|߷o�ٳG��y��#�^x����z!2qco������)S���ܶ�'��u]PAu/����Y���uM�E,�cA�S<]G����m+(��:�l������������n   �%��E:�e:]q��y����O]A|���� v ٣r/-)����4�~<}��?�1,>����on��U�sn*�Ǖ�U���(���  ��C=qZ���>��B�[i�����y�����d)�!����Y�R�b�&w�r�0{�D�;@����1*�`T��0��x�~����ӵTs�ί�����:JF8��^ {���޽;�C4��yx���o�7�?� ������`%�0����<�0���?�u>������!:b%��Ot��Y]�e�f�㳝whjl7z����Vx� �pA� P0��;H�6�MC�spW�H5�f�����-M�j���Πr�G��SU~��޷!�v,�a��Fu��Z?�u���<��~�ۭ)++��S�����z���t��Ajkk��9��Y���w�t��wd�iڴi��ֹ���;��Չ����?W��g��a͏J�=��A��Z�]>�����)��(J�ۇ�x�V�A	T�p{M�$z��x�s�    ��Ɍ�h��zq4N�D��^#<���Φ�4c����������ڄ������G�;'Аyqq]z�QTVZb;�w-��^��  ���S�c4kB#�9�u��,�Rx�v>��3Lq�!=�d)����n~��3T�����=ƨݳ�n6�OX�>o7Gw^�>�j>{M�����:���> {���ݻW��G.�b���=A~��w8��>"��`��"�y������y�0����+��Ϛ\��^�flO>�Ɯ�B'�P'��KU�%w}6z�N�v���� r	� ���/F���:kv5적�e�}�g�{��!�����1)J%���`�ngP�18�ݕBU©��y�5��m��k�^�ϵ������l��5�n����<����Ǐ���f�:�����]Z|�@<������9"��2$��d�L�Ϛ[�u��,6qX]���o�ǡu��5�x�l?����R�ҙ3������`��u��	Tn"U�@������H��J����8e#T�aG���bӐ0�    <k+iѼ��q*5�����@G�j���2�׼纳�S��0X����W�D`l���Կ<0|�8d��ΜsB�nnG�   ��l��ʎ	����۶�6�;5��=C���g�tO��N~�Sݭ�@�[2�a����{�l�u>��΅q^wN6����o��Ǫ����w��A��d����â��[4�Ỻ��	�߭��V��9�.K���ȏf�9����:�|a�/�@���\����G��h'���96>�f�]5��;��<�f��Ss;��E�i�fx� �܁�; � yi� M��AM��C��*KC�j�A��3� 9�B�jB{��-�n��B��qB&�Aw�k����ky=�e���~���ӽ���:��]�~ܸqB a��	���? ��w�X�������uww�G����k�:��|c����9��0:�` �F|��cT�F~]YY)>��dh]պn�~A~�a�Z��B�}�V�
�g
PjQJ>�Sv�J�rn^H
S*��CFN┛X�!NY������j�M��CB�}    @���b��=Wӵ���Ǖ�Љ-�)Nh�No��5�[p��g���x�r�n���n   ��}J"A��&��f:�b?�vw�c<C�b,'��tO�~�ݟ����/t���'�w������Y��u��չ��g3G5/��v��ָ�eo������'�eX���k.������9��x/�h��g͞����G���ȏ�{��<�����񱅱&�"��hy�N�vU������7Tc�J���T!w��m[ە��A����?�N�M�	�!  � � (X��i��J����J;��@���T��M��*^��dh-ns���:�U�@�
���)e;���݃���x�k���|6s���4�n������u�ð�,�� ��F��xX������/������M����O/�S��y�K�����y�?^kC:��s����5, �Z~�ya�7^���Q���WH�U���(۽�.X*'q�*R����[:	S��*q��|h(F�&ϥ՛�?Ʊ   |[�ݿ�2�p{�����;.�~�D��-�rG�    *�;�-��芦��{`��˩���3t�GJ0JD)���w6��N>�*�Ϊ��P��ݑbш՘�����l��s/k�:��|�s���^��~׸�ӽ�g:Y���8 /��dA?�k~Ώ|�\~d����c흃���a�{�Mx޺^���s��s\Iϐ��9B��X�Cz�\�%K�x�]���	
��
�Gr^ء�B��St
���vav��خ
�����_���Yz���X���1��<�Vo.���  @�A� P�<�%F�&̥3�PW�!�wK3�]��Ѹ��%i��*Z���V�*�vϾ�!-RY�a݃���������a�Q��:�i���u:�u���VX���d#@�AX�\�o.��|�)��t.�aS�q�`�v�✟��P�N�1���ܮl�c\y�(�K�6"�   ���	մ���PY�8��N�H[�"0��w��v`d�������T���c?  ��Ѫ�Et��y4�v%���EXr�D_���_(���tC�� �vhh���C!V����~�{ϵ_����=�����\'�yNs�Yc���5t��H���~�?���,̒�w���G>�H���",�\"˲�9�3ң���#9Yv�A~>x�_��~�k��a�ٽ�j�C��a{�z�v�o�s���D/�X1�o����������(m�u�� �� �Q���!Z�QC7M����6���h�r�n;h/Z�W���Z�6�w#|���N�=�k��o.��9�v}���z=��~�;����~��|�sE��l�YH�U���ۜ��=�v��W��M�2�q�l���L�J'�.�C��z�Lzb�8�@�   �B�ނ��q�0��W��v`徧�   `�=��Z>�.��O�v9�����_8����<Y����ٮ�]wh~��;�ɡ+M�Aw/ss�hw���z�A�����<�s��;�q[�{/��sm;d��s#z��Q���X�^��B��z}~���?̗��9�n|�!���zkn���Y��n��M��zb{9u � �/� F�D�~s�fMh�3'�Sב6s3�%��7oeeeC�i�*!�hemrWW��(P��|lCn�]g��k��o��}�nN�Ts���Y��^�^��{E�\�[A�W�Av���t��C�ʧ���j����.�Sn���v�慌-]�����l.�m�Z�    >�w��{�>v������c�\��n   �W:�㴢��Θ5���v���Tm�C�P�z^<Ä��=�3T7�K�Q��8�Hw>(mOct�/rnX�A�	{��|6s��S��3�m��:������~�R�+a}��\7J>b<��j�:��`��[L���j��3[�ݛ�UM�w�;>������ho�\z�!  " � u�l����j:�q�uo���&��Q�hu/f�J�ɽ���n|���]�!����	'���0ƣp���l�d3�i��|�5٬ӹ���e�^����r)\fם�*Z��l�j�nw�2B�6�v��v�(e	�Ũ�~�nk1����
   䚿���hׁv:�e:�n�N?��k �!��������i��ρ#]�W�� �B�    �yeg�*˦Ӓ�C�{p{�Gh|���.)����EX����T��̇�3����aw�9��\d����	Y+MN��=7��ר�yY���9���;�n��:��^���A�g�ȇ��{��N>������=_H�a��&}>��1؞��p清٭ޡ:Ю*Ʋ�=�ۍ��n;>?������ �� �Q��[c4�f6�;��:���*cC|D���Mv�R�J(E���;?�5��s�{��=)^�2�G;��>�n��\�=��a���F���@D�=���7�^"?�G�E��ȅ��{��F>E+V��úFX�v��}۝�!��l�n�i_�[VV��{S�Ϣya� D��2��������c��/��o�F�O���+� �Nl����?|�     �L�`�V��I�[��x/���f��������_(�C�h�'ˮ�7Xl��EYf��vW=�|C"��{&�Aw>g�����ָ��习�g3'�yNs�滭qZ��V�:~��{:a�>��f�>�h�s��c��\����j�����{k{�?��5�C���iO���7  Z��  ��5D˻�����г�L��!��屙�D4�g
V��uI|$��ʐzW�38
V���vB�݃��xPkt��g��|�s���^��nk�Y��ϵ�y��N�F�������&XEM��f��`��5�n=�_���ڮlO=7���ۇ��� U�ϥG�� Z� yd��)��_���*ʨP�?w.��O�Ow�!�w��        D�������tYc���n,�Rce��ʂ,�����]����ZK���aAw�\����x���r��Z��A�Q�j���uNk�\��5�z���+?4���{�0��ss1�a���6�*��mm��S�e-Ʋ��9�ھ���� �	� �1��7TϢ��Pg�>��A���k����^j���A�*IXR��kfP�3�V�\܅'U&�=���e�'~�=�k�\'�k��r���{�N6��:��f��z/���ڣ�0E�|	Wa�VA�Kt�fm��|ە��,����TZ���g���,���}�[��h���  ��ʳ�-�p���E-���>I�|�!z�        ���H���8���K�ͽ����!����Y�Xb�g���k�	3=ôo(�B�2,�mН�a�L��ۍ�������g�%�Y��:N��v���u:ku���Zپ�X"�?�l�1(1����^+W�b �v�q���^)V\x�q�p��_��Z<C���մmp��!r �肀; `�p�;N�7U�y��4�{���������f'�J�?�+u�]������&X����aw
/�n7D ^�:�^��9/k��׽F6��u���:��^����^�eX>*"ZP���x]����X�r���į��v�P�Qx��T[	*ũ�{��vǐ��qA!P�{����zs�bq�� Ѡ���F���w3��ï�������!       }��ѻ�tyc�zns�
u��Lb���$]�e�:�3L���v��_�]�u� ���h��K�z�n�}�l<� ��:�
�=
�\��پG�Av/��C���^���3�>�ڽ��z�X�?O��q��v�R,�r����x̰�3�C @�A� 0����!�X9�.�5H=v��*v763ȃ�(�6��X%�b�kc��]�=�Ҡ����0{F��p�K�=��nܫ��GPMU���a�SA	S^ĉ0Ũ��γ%��G6�-4�j�	V��t�l�	��*;a�*Nŕ�v��v[q�F���0���D�Z��   Z������Ӥ�U4�/U���:c�\��7K��       ���K�6��Σ���Qow��+4���w�]��c�6�!�۔c�����g�{�]!���;e�s� ���:����e{^wN6����o�Fw��z/���=@�N����/�@���B���v�]�7��ΥXv�v��K:�a�?T��Z|Ī�Z���@��; � �$�{�rc	�4}5�ޞ��f�J��n|���`If轘�܋�����@e|W�e��[�=��������ݸW�����`������09��QD����$,!�,0&���:\��e�1��p}1~��t16� ,�BB�&�
	�6�<;;3;������]�U�=�=��<�U����ݙ�>���mC{�Tq����S��+�4� �$�!�%�̨k,�h���v�Z���^��.3���/(��v��JmW	T�k���v|f_��qS�"���f�'��/F7�ԝ����o|�m��c�A!�B!�3��<~����;֠8u K��Z�,���^����X���:_FY/�%e���F�F�;GU\)�B]/n�1�qI�������5�o�Nܵ��f��e~3��c�������v0����f�X���d�g��G�0�4��8{&��{�\��CBHgA�;!dE���~����vL"w�``���T�ҋUA�{:dr�Y�p:�:��,�=���5�W�"�AP��*\�i�=�fN����㌉3N5V6^7G5�d��:Q�L��Dҟs���E��`պ��ϯʟ����{N�خ�D&��P��-x�)_Q���n N9�������8s��j��BړO�� ��S��������΍��q�'F������_�'�� !�B!�t�"p��"6�]�������i�(	�2�f2�]�3�w�齱��I��$�����V���϶��c��/�c:W7�f��k���F��c&��V����n2�]j���f�	e�4���Ac�>��ZS��}>%�]�%�X��G&��;gFpxw�҉��NY����mc�q��4f�Ψ�ڑъU^�{Ɠ��ن0��`"V��M��u��sx�!�'\�m�=�tN�}���#��X��y��6kخ��sڝV�ZI<'���Zi|��*�9I	SBc�����]%L٤.�M�E��]"N9cu�v��� ��p��"|ew���A!��'�~ ��ǿz?>��W��'oю����~�Ÿ��u���*��\&�Bl�����ç�y�����k^�}=~����U95��>t��D!]��s��!<c�*�^:���Ey0VM�Z�e&�t5+S�vk���B](�������jT�BY{+눦�M��yQ�u�G]�v=�X�x��\��&�D]ӆ�6�7�f|Nq׌��(ɱI�[�����L�6�a�z�O�����vQ]�|U�����QR۳==X߁��:�v��	!��R���B�Ƴ.ê���U����D���g�s3�T��p�VoA(>ĦvS�;R�4wS���7�pՌ���ү[?�:��َU���3�k�F���>g����%�Z�$Z��tc�!h��`9q�s�3�#,T��)qJfrڋ�R��$/8�v���~`)�!���053�_�����%xٳ.3���{:��e���Oczn�B�3<Ћ[�������+�?åx�{n�<�'ֺOܺ���g��lZ�
����@!�3��`�}�p��<.�:�Ɗft��ce�C���&��L�T7��B�|5�XFwu V���ͪ��J2�j��q�����ج���V�>�z^�k���۩��R�n��z��nin��u�X�ݞU�C[c{AQ?Z�	w���	�	!�����،7/	E+��@� �5����U�av�&��7��z�mA�2�����o��bV�;�NQ�+*-���*[�i9RLװY/���@+���ψ:��(�q�(XE]���v�0�0�{�f���-�>A��Id�6�����}xl�����yBi>K������ޣg�~�ќg_�_y�����I�>r�B���?�Gs�CO6��{�Kq���:뽏c����J
=!�����b	�}<�K���%}'17;�B�����Za�������3鴴f(JxW�
EFw��V�Z���֕�������؊Za��	[��['�I<�i��g�f��m�'Q4�jS��/���}���ZTG,�$al��ݭB��EiZ��~hR7��XC�8�[����3!�����B��/TD�+7����1��]h��%�"����^7�ׅ�tM�R�V^c�hB����]dr�}BCu�@kJ���B�l�8k���g�jl��9�sMְ]+��q�򱵻8���׮��J����^��w�2��)��=���$�|[

��u$qJ��༎XۉO�w��e� ��N�����[����f�o����5���'p��y#���������$C�?2\�͘�_�_�[xp�QҎ\�k#����+J������G��p�__{�x�SwT�3�_�[�ɡS ��P/��]�ŵO����P?N,͢�x����<��!���<z2����q�I�`i�X��.�cej;?�ꆞݟӁDw�Za��.��ꄲ�Za�SW�5�Wi���^��(곙�?꘸�����k���I=�ShU-2�s��_N3��85����Z?��mRs;�glW݅��ޠ,�k]Qu�u�R��:ar+�����3!�����B<p,��ӫq�4J����(�Fw��r��	T�d�h%JbPA�JezwE�PbC���	W&�����(P%adoq�V0�)Z-F��Yݡ��rW�)ZQ��k�	S�6��]fn�S�Rja�����-�S����<Vo���8��vBYN>�����s���#�}���#��_�w�ӝ��/��q^�����^�K�m���;�ǻ?t�Y$"���;7�s�y=�{*�/.������
��ןǱ33�v.޼���_�+/�To���]x�-�$g�������w�?u�Va���<�S�gnw���V^/���>��B�\�E���El^��M���ٓ�zB�X���탱j;=W±j��tc��t:S�:uÒ�(6��0�;���vqHVR��f��ev��3&�8��(�esL皬e���Y�$����^��6c;����CQ��=G1������R�v(���2�ڄb�r9�N�÷N��n&�B��	!D�+Z�l�s7�p���Ƌ������
ƂU�^��^��i��u��n&Zɶ#T��+S@�
&4�W^�s��[)^�ε�Or�l��zQ�U�1���o�NԵ���f���Z�ώ��r�VI	[� Xٴ���ʟ!a�&q!hn׉RraJ����D���v���T�v�Y5�������P��%��*���=x�;?�y�k�qrT;>�I�O��\r�:�����|��veۺq����I�~��w�'�~�����g���.ϼ|;���^�_z��v��W\���66<�_�ux���H�3�׃���ո��m�����������ٲv�?�7��6B�|O�q�� ��t1��8�/�IC�t�X^c��v�A!]������j�06�7�%e����4�CP+����^�.��$k��#��X�x��\�5l֋�~7��zc��[QG\�b�1�T?tk��ks���6�#z�5��4�Cݎ�E���m���8ݷw�uj�Ԛ	!��b��|�}<�K��ē�`���P�*8i��v�A���v�Ӂ4w��=�ۊ�6����.<"Wbӻ;O'8-gC�s��o�N�q����9����M։�f���T���-�p�ѪU�vݘVVI�	�Q�k� 垅�v�E)���.Om��.Ȅ)�8���ٞ,�l�m�
�ϖ���n<��D%%���z-��u��'Yy�����ƅ&��#�tJї!�DO6#l���w���1z����7����W�˷����Ư���R��N�E�=�����w~�B�������$nڱũXZ
�b	v���EuB�>�螮��ݟӵ���^<µC��=���I�0��@Tt�hM�^�lC{�Zb��Q�Q�wl�9�y�kخu�($Y�l�e�S+��Q�$eV7���N�6�]������v���X��a����vO����܊/���B��	!ĒGN��hjϽhٹ�X\\�T2���hUOe���}�L���c�V1���/�������/��fn���k�g;V5^5G7�d���k&��v��WR�k� e;>I��J�T?c�"���njn���4��S�����;���;�z�:Ѓ��o� ��n�1���|����YO�a4��/����z��=�ĩss �BV����s���Re�V��<\�]�����Ç��n��y�D�8	B!�A��������u�9}�������2��Q0�~UIt���+��42io������U�CY���ae-T+����ܠS�qj����1����	uu�(�E�<��6kE]7�hJ�Ѭ�90�'Y4�I5BU_�����ިz��5C��uĠ�=�`,��a��S��}dr�ur�v3���r���B"P*�pϾ�6���K�?}H��P7�[�V��Zz{��^3��ū���o V��V��(��c|�E,��=(^uj�m�16�Dc���g3_�F���z^7ӌ�A�5�m�o�e2�S+���L�
�	�="�J��nl7���2S�ij�t;A�0���02��yfw���!���[����_��o|���k��\�k#���7�����!��R����#�|��?����~�>�G��h����w|0����7]�?닐I���;��|��q���#���!�t�g
�m�Wm܅��0;��f�Z��ce�i�3��au�g]�Pot7��j���ݩ�ðD&wO���6�����Ю����7g��X����t�mױ]ׄv�Z��fR�n���v|��u��P?tk���`��gh�T���!6s�ga�Г�^Lj�g��}pdGrk�=Nb;k������s�|��vN��U��03uFlt���]Ѫ��P۽}��N�Bp+B_�{����Xw�_�	Xq������+���C��W��:&�$Ǜ�3�o���zI<�i����s�md��*C�ɘv��)���ڤ����8��R�X��*a�4yAgn����ف�𕽎с���iʿk���_��#��_}>���v��uc��{_�W���x��iB!�NoO��x�;�c��������ct
�����/�o��2�h~�_�y5���7�>p!�t����j<�����Vw�ݣ��{��i��d�p�P���EuBU��^3T�
h3Ǽ^���v�c��j|7�k�N�5�~v�ӌ�3Κ�TGl�����=�z��0Kan��
��v������r�3��w{��:�k1y>��<��!��Dhp'���s6��SCx��1L,��¢��.2�{�L���@��$�;/�3&_�J���"C�N�Bɟ�Jw�
Yu��T���iN�{����3&�8�X�xݜ8�Lֈ�^�g�t���R�J��n:n%V��=���@�����f�S!c���]+T�Rڝ1����ԉm��~ W`�!�t:��>�9z���:6ܯ�qr_��o�k��_�Оc �B�����[^���%�o���o���½������;/��'�7��j����{�B��B�T�zrp��qs��C�l����X�za:�������&F�p@�,KV?@#�]P/t��Z��T/����K���u�f�u��(u�8u�n�ju-4��E]c���PC�:7������m�b�j���y;>7�v(Ih��<Wo�=�{q�N_!d�B�;!�$D�����ѓY����P:w��� 2����#Ni��Gu���6���kpw�+q��_��
`�v���J�R�VH�&5x�j|���,P�R�JZ��*�A��K������%Z�����v��=�2����>w����+J�
Tbc{8q�&�����Z�	�8ևS{��N!��7ڋ�����xu%�U��� >�'�����G���� �B���l�����MO�X:��Ǐ���/�S����s�߾�Ȥ������N��/���@!�{9s�������ɝ�j�<�O��E&wQ8�*KT/,�ϕ��t�����[4��YP/��~X�!.s�0�z���g[�z��:a3j���;�+I�[mog��Z�Y��u�V���?	û��n��^4��°LM��@�(�v���X��G���,+���I<<;��vB�� �����0�B	w�.a�+����ų��"U&S9g<��x�3�{��G���+)�{��v抅�F���]eh�ۅ�D�B�>���;w9��Q�u�G]G�Vܱ&s���͏�V��mh�a��ĳ$?��ku�hWpҍi�`e���Kk�S6N�r�('��D���*H�)�HezxS�[	��\.�щI<p~�w;�v��	!��w�,^t�?���r<����}�Ļ^������g@!�t�����x9n��	�1������),,u���N��գ��.ߎ�/݆o?r �B���g
�cWoZ������ka��>���f������F�{�V743��v�.Z�e��RJR/���F�$��~լ�8���c2O5�f���xF'ӊ�c�hE-�Sk�]Q?�=}����=j��ol��G����5�����ކ��w�s�gBq���B�Ĺ�">�;���;p��,f�G��Ne����e�����3��(d���sc+Bw�´O�*
�)�x�No��D�RP��Լ�R�W��̵헍1W�R��:G5�t��ZQ׍B;�ϣ���!�ڝ(Z-�`����~��T"s{]�
�SPS��TC��T%�0��.��m`0�=�8�D"U��ў��s�#L��N!�ι���O>������M/�F;~��0>����uo�B!�»�p3���'J�S���S8~v���~�۸l�z��Y�)ǽ�Ƨ��N!+�����`z7^���#����vۚ��ѽ�F!�c�����eY~�{��,�}�xh]mPD�^��Wͪ&mx�;�d�j��\�5l׊�R%ɯU�k��jh׍i����X`��α�F�
�>c�[O�R;���~�w2&/¿�-"_����M!̀wBi2����Wo��2'1w�|������t����zPbt�$4�[����긆ѽ0��ī��p�%O�{I��,�������(╮�*۔�V�2��ۮc���NHkX.�-����n;����ɘV	V"�{4�W�i��SAs{�^'D�M������h�T�ąb��n+N��$i�nOo/��[��}��S!d%�/��y�?ށ���{���d���;6N`��!���!��l���9o����}��-���x�;1>2 3��B!+�|�koý�p��"rg��Fa��1�v�c��F�U���Z�LwOůF�V��k��M0�m���(�Q��'�u�n��|ӵ�X��iv�1���6�یo'�{�L�?������ZX?Ԙۣ�c�R����n�2c{QQCtk��`,Y�й/��X�	w����"!�����BZ�}Gr�~j�ܶ�G�����j[f���*��=]��F�t�yX���Waӻ(�A$T��#�w\I��P���jv�6���Q�����5]'�I>��h�����6�����_�����e�vq�^���Ku�)���7��D)o_P�%/�D*�[���u(���8��~�B��|�'F��W>K;vx��wB!+�o�`/��G�mL�-�o>{/����@!��]*⋻�#��0{������R��Za�0+����]�tZ�%��hlv��/F��^��Kv�@{ۖ��n�gL�q��Q�����ͷY'���,�Y�]j���en��b��[Y?�ĊR7�����}��'ê�-�۵��ڡ3ndb�sv�/Կ��B���N!-�TJ����]���
�U�!��]�*�
W��z��ճ7��*<�fw�V�A��3���UB��ZD+�`����yY��~]��[�J׿�U3����1���k���I=��i���ĳ���ܢUR�V;�ڽ�2��J��\��E����]����N�!>U���2c�I
���^_�]�z3�u�'vS�"�Re~1g4��� �BV����~�#w~oճ0ĤvB!����^\�v'�<p��S(z�5à���p4�t��^pj�Հ,��銮��
�y�T�p,�к@,i��фe�Bxj���)I��m��Or��8��(�ustsM盬g][��l���|���m�v3���4�~轎U?���jMj�~S�8KV;t昄byw{V�
��à�]XC�axt��V�+{���B�C�;!�,sK�J:�X�V<ws�gU^�z������D�L�$_Oi(��kUE��V���oBC
�t�`��+b��U�6�@)�����&�T�cf�X��~�x�Jן�@�t�B3tsT�L暮e���Zi$�5ie���$+�q�Ni��*W>*<���.�l����H6��*I�ab���.��y�L��}S�ط��!������.U�)�����R��?!��Ng��"�}�_v!�������(��m�K�1a���s=��S3decc5v��xj�ձ��u�X&�wY�[#,���B�{_�U�FX��k���4��g�4��̍2?�:6k��F/�c:W7�t�(��褠��y&��V��U�_��iW?\�ꉡ1�uCy�P����j����Xn1�ecn7�r���!Ln�W:�����ބ�hp'��e��B�۝��n��O�g�b�#RE��9����h��oE�Mh(8�����P��"VY���L�$43�'mv�2�t�8���c2O5�f���xF7�
1+�gD]c9L�-�`e*J�*A*hh���P:a*(R�D)�����S۽T����ctb��M�ѽN:/�)B!�z�w�
�m_/��*���2>��A!���`v~	�B�	�Й�<c�zL.���B=Kdv���[� �]U��Za����Ou�c�±��Bw��Ю������Ix/٦����n�/c:��u�f�Mkw6�I�WjPV3>�kv[(�ɘV�ڽ׉�k��u��9�ebp��ښ�m������4�_�W�+�vH!Q���Bڀc3|v&�ͫv��0w�2�=�1��ݽ�����y�"LW��p�	�ݽ�U�DwU{5L��aP�j$�7�W�%6�&5z0����c3N4�f]��U�L暬a�V�g$��?F�;I~��L_���J1�dL�M� �d�.yAdjW����5�&N�S��V�R�������V��}��=B!�KO6���W�K�I�8�Z������}B!�{��+!�;
�7��ѽ'��ݖB��,..�j���,whC�{#�V3�
����ݠ3��kvO�����p�p��i�P�elx70��k������7g��X�x��<���kخ��ڝV�%�1�f�r�e�QL��Zb�@�(�X*C��nX�����s{�f�����n�U��Ln��SX�Q�]C!$
4�BHqx:_>��5�W�������*����4��E,�V�+Sߎ0lv�OtW	XJs���
V��╍��;V$^U�,�@e*:%�����k��g�f�n��f<ힾ`;�U�v�1I��E����.PA/N��(}ꂙ0��m#�M\T6�	����^qjpx����N���B�d����m/�O_�K:��vB!�{�U��B�=�B	w�-a�w#��������=�0��k�L��Za�Z�s�a��.�Z����ٽ��:}ڀ,Ϙ�x�+�7�;$evO�?��q��I�Wͳ��[#�zI<k���ץյ�f��P,ﵸ~Ni�^�������bi���X��[p��fN��C!��	!��}�P>�����������>�L�G.V�CbU��6����t(��/Z�����u�v�X���̠.�/X�E�� ։U+ĩVSq����⬳�fv�q�����W��\��R�I&�TP�2M\���(#a�.H�)�(�^�Sn�+:��^c{� �$������_^�K�chn'�B��|�wB!�[*������V<gS�g�w����J��*�]�Up�f�J��thY��,ѽh]/��9z��F(���>f�f��S�Mj�ɼ��۬��3��V��#+ʼn��^��~hS;����Xn��&KW/�1���׳r�y��v;Fw�$������Bژ����Fq��Il�I��L#�0�{��A�J.V5��΋wg�\��
P�T���%Kso�W:s��_���	V��aa��A�j�Ѹ���������7Y'κ6����Y4�s[�j9L�E�*J���qE���)[�{0�]lj
S��V����8��J0�䅠0U(���ߏ�ѭ�}����	!��y�n�/�|����vB!�����!���L���)lَ��-b���J U�&�0��±d5Co{�����T�Y�P��Ov�6��4Yh���kVI��^��_˶'���qꋪ�Q׋󌨴����?�V�m�tf(V�OߵI��=�j�qꇪڡ��4���É�ạ���&˙;�z�=ч�;����B��wB� �}(W�sWoZ����1;=-��I�"�J���	Wn:C8��MhHi��Tw[�J�ր�f� ����$*�)iq���6�DY7�g��!t%��8k,w���R��Ȧv�E)�X�JYP%.xSt�viZ���^�T*qJ(X�b�����o ��-���"���!����ů��:i?��B�ʀ	�B���L���b��.<m�fN����u@�]��j�DwQ�Pov�����B_}���)y�!�.��m��b�_߷	�J2�*�8�X�xٜ8�L�ۮg��I=H3?��Ċ2�SB��5�h�C��)&]?��E�<�M�f5Dub{�;>;s�'7�N��n�	!����N!�}G�c�z�jlϜ���s�4�um;B�m��>�nr��W��y�������TwSs{���L��aqJ���k��J����Q�����7Y'�I=�[i���U3��c�ѥ,4�����Ȧv4)��Qڂ���T$�= J��)m�T�j��p���iJ �bƛ_t-���gJ�in�l~꒭+z��r��?B!f,,�A!�4�}g����v���Dw�.вCU3,k�<��y���^ب����UcP�'���uB�k�:�{wl�.X[�cE�6��+��g�n~����mB;�e-w]3����n;���?=��{+S{m����t����^�%��k����}5Ī�ݴf%�bl_��?;�}{��{4�BH����B:���}��0�]}S�9w�BOU�*��v|��4w��cvW�=�n:C]��$4�5)��?��4��F�
�W�������L���֬�i/�*��׼�t2�ɚI=��h����s�-}�fl���{[S{Q�T�R���L�!J'L�M�6�TE�����il'��W��T�ɛ�/���y�s.�+���y�������σ/�=��O��� ~|��z�O@r��BH�9|�P>�ؼj�>��4�g�XYA0��fX�/hk��`,�ٽQ/�	E�B띠�/T�N��ژ݃aX���k�����Ǌ3�t��ZQִa�M孠[�l�%Y4�|(����#��S?���Mj�E;>G	�
cy�����ؾ�1��?3BH����B:���� Fp�q��¬ct�d�[J��u�����Mh���S�i�v��*lz�W֢UL�����,�ݡ�w�ؤǫ���׭e���Y�$�u��^3��6��&0$���^�)�����J�����lA��]������.L��s�@�F����E�4�B���=�/��X��I70>2����yx��n!.�_��닰k�d���w��%>5Bځ�S���cgf0��Դ��d3 �BZ���|��ݯ�\ąSG�N��B��]op�c��I0�,�]�t�/z�Phv�^���(�����V��p�8�t�mױY3�����&����U�3t-�ދ�[ej��AX��D�nϚ��vE0�kl�ޙA���B��	!��g��T�(��*�]w]��3C{�Y�L��^��Fw��]gt�%ZE0��Xa�_�
��t4S�R�Mj��<���kجw�n�BVψ��r�Vq��{��]�� � ��(%J[�Q��R=e!dl�R:a�(��+F)�)�	!����W��?��e��=����[p�3Ǧ5�p��eR�K��3��e��n�j������7��rL�&��7������~�F��A|�?��󝸰�k�s�{Y�#��Z�F�6�ڎk'��Fwg��[�=fwS�{�Z��N���mw�v�]��R3��vh���:8�U��V�	��M暮u�$��h�ע��XQ�td(Vm�I�7&����n����kl����#�B�L��v{.T�;�z#���P]#��.�5�_�i�{�p��)�=�D��#T��EB���^7�=�fFw��]gtOJ��	Wrӻ^�RWĒ��+��g��Q׋�~�a�oW�,ɏ���U�dbT��&��)�Y$L!,P�B��R���onۃm&��+JI���8�����kq����B"s͓��÷�
�=�V��I7�fl�wR������7r�{��I��ן����عq�=�G��h�3��4!�����t�jtێ�O,`���ݟ� -��]ft��ܫ5�zm�`Z/T�dk�&�l���fA}��s4xO�*C{��k���%�c2O5�f�5�zN�Ҫ�rbE���X�{��]gf��Uw�N����i��e�=ۆb9׾�����88�	�9ُ�4�BH[@�;!�t!���>�I��q��fOEڛ����>m(Z5�_R���.Ou/
�դ���e��^;�J�t���U�oU��w[K4.���9q�η]/��QiW3�	�����n��M� 7e�'FI����v��]�� Ml�l%hcp�R���U�8�I�y(W��i�!��˶�ǿ��5�����N��S�x��)BH'����'�!���>W(=X3��m(�p�0��4wQ8VV��n�tu�碸^�	�Y�-?�M�nOY'�uBQ}��0��k��Ú_+�p,��&kDY/�sH�_�Vb��Y�P��g�P,�k�I�eFwۺ��~�6��Ų�r��'7�;�{pl��Ec;!��4�BH��ӹ�ы�c;+[.�9Ry���U������L �Amp�EFw�x%��fv{�*������9��%�9���cM�ę��e�(k7�٭`9Ŷ$��*#��$��{��=x��`.F�V�w#S���]kj�Ra�z�12�?��
t��w�)
քB��k�$>�?�����4��n��o�:�s ���	�BڅSs|q70ҷ7lR3G���X�Jñ,w�6��
���ڢ��]it��5C�w�6C���Vخ�X��6kجw�n����$�oE-��k��dvQ�����6�G���ljl�
����d��l=�[��i�;�۹�3!��4�B�
��А���필�⹪p��nC(Hq���%��kG!�nW�9[6��īD��oM��gub��oKoxwƸ�q�)���sT�L�۬eͤ��-4��mu���<��*�)x��'�IX��ݳV���%��L*�ąVۃ�T�ޙ;�z���NZ;�X�B�m�8>�'��ի���4��n��؃��u?!��ѓ���BH{1�X�����ܰ%�U��1��n0�%�����Xz��xG�X&�`[��_3t��n��
�}���5���g2�d۵��oK+L��V�l�@��s���.Kiw�6f��M}Poj��뇲 ����8�C���?Џ��|� 0��vBighp'�����0Է�ڒBj�(B��.�l�A�*$RL﮹=,`�ܛkvwϦ���3*��-���]8J!dU׷���ʠ�o��͚I?�]i�����Zad7����6�%Oi	Qq�)[c�wKA�%�B�$Ol	T6┱0%Mj�
S�ԁɍ��>��@!�$������^W9�p~O����E|ꞇ@������i�&�b��H!��#Ky��}dRk�S[2X�S�;?�L&[Im/xM�
���t:��!��U0���.�#���}ú2˨Vب��;3K5�t��Zq׎B��ϣ���#���6��Ƌk�Qj��P�����y�P�'6����v��(6��LﶡXEo2��v�0��142�ٵ��@��HS;!�t4�B�
dn��;v�Л]��l͠g��/�V�+�P��sD���-hxw�&�6����H<��*�>~�{H�*�S�e�jbCt���?xWH��0�����5]'�I<o%ь�I��/�'Q[�v�lml�_t
�ۘ�U�vS��q��:S{lc�H�*�����̃BI���A��ǯ�$�����B!^F�@!��3����{:�8�ܰ�����(d{�fv��=_3�g"ݥfw�`,U�0z@��͘P��5�W)j��tw�{g�c���ͷY'���zv+Y�z�rbE�ۑ�Xh�
��q�Q�������2��$�+���`��WM�8&q�\��f(!�t4�B�
�Ih�ko���mO۸���c��I��[����Q����I:C���¦wo:�_�R�uVbIn_������W���V��qL�9&�Tsmְ]3��t:���xN�5�kf���ڃg[�*�������5���{]�
T­���R�c���(�zW��X8Y��A!����	�0<�9�/��;_w#��e���1����vB!�����Svl !��)<p,�0��n�O����'�L��@�����`,}8����R��lk����q��=�����a��c���7Y'κI?�[h��w�V�bk��1I�����Q���ݞm���FvuP�M�0N0V�X���:<va̡���	!�ӡ��BH�MH
���>b��.\9���3G��吕l;4��W�6_2�"��'ZU��)�\�����(����`�m
ux���F��P]����bD\Aj%
PqI�k���(fvQ�J���k�ܳNhR������]-N����%�(��n+L9���$��qW%q��vB�^tݓ�O��
t���V��	!�+:�?���^S��zA!�t��!`��N\3�G~�(�&wY�6+X7��c�$uÔ~hS��C�b�Ѩf(��g��=�i]�O�±L��曮eݤ��δ�6���X&s��Նv�b��.�/F�ǩ°T�X���1�;=[�5D��{��F���>���s �ҹ��N!�Ǿ����h�6<cK
��cXXXP�ӆ�h%Mo�T)���#V�,u������ ﶇΆ����+dU�*q*���%Jp���-`y�)[A����4[�j�p%����P�v�%IV�L41��ۓ2������K>!��KZ(9�Yj�h���@0�;�6&6����س����@!�DO6�w��ft����3��B��u�n��.���ĺ�a��/� B!��9|�P>R�݂�7�'qan��ӳ. +b0V�:F0��f���k�q�����u��|g�ذ�]M�.hj�O"K5�t�n�(�%���H;b�η�#�k��6+C{m�V�b9��&5�j-�����I�j�1�����&|�H��P�B�thp'�"��b	w�.!�Z���҃���9w6dtO7S��4��vW��W�_̒	W�k���!�p�4��g��G�

Yr�Jnz�!(�J��#J%)�,�Y�]�$?;V&@U�۪��4BTm��=Ч�T�]֧�䂔{�
P��D�*�*]b�N�*Z�T}����&�{$���NZ;�)B�D^�`�1tnr;��B���'�)�����!_(���G�x���#��t���%B!���Rw�2�5�r�zl�;���'�v��6fw�v�n/ˬfh��N(4�W/��@����\�W8Vu��Ȋ�n�u��bU���ۣ�U�X��ø�X��p�Q7�٣��,7����l�
��cx�N�'��9*_�!�t4�BQR(�p�A�D8������C�1{�DE�		V5�Ig��m7h-\	D�T$�{X�
�''\i��:�{@�r�t�"ӻ_����-U�C*Ԟ�0���b2O�f~^�I""��Dl
�Uۍ�����>�H%��������.3��)�/(L	)ߘ�Z^*�@%�T&�|>�щI�(M�s(w�JEB�\.Z?�n�5��Js;!���=�6N��%7\*�[���ʹL��x޵OԎ���kB!�E��>��#y܇Al�؅+'1�HE��x��@,�]�ͮ��R�z���ݮf���~]���u5�(�X���	v5�v	�2}F҈>�N�?._ V�O��`}Ѥ���хb�ꋒ�$C�d�2C�I0�p�g���_[l�m���*��;�f~pn?9�ݞ	!�����B�1��!`��N<}CٹX�_���t��]gxo�W�����6��d��^,`9D1�[ޫ7���M��P��$Tɍ��5S����L��щi�%|EKè�i�'2���M���kk
~�)x61�R:a*(H	��KQ��$fv�*$Li�|�g����p���0E!��w9��������4�B!�8��o���U4�?��n0�����o����q�}�`�5!�ҩ�;�/�ڎ�6Q:���v�B�.жuC]0V��(Ʋ����8�w�}�&tv�Hk��;<}�p,����F(C��$��&k%�~3hW3{�?�$�����p{�Ϥ�(5�{��bk�"c{5C�ݻ˳��=�3���^������ݞ�ñ$��j�{}�}�ݞ�s4�3��BV4�B���\��v�#\�+7f���OW�U��$��L�:�*hzO����]���䞄�]kx�VB!�}�h'8��(43�˷5ԭ�Ώb����� ծ�R+��5������r�{���׆��(���ꐛ���T8��+N�)�6�:qJij7L_p�9I?ëVa&;�of�P�"��n��؃�����]����Ӡ��B��1���_|�����'K�u���5?}��-?�5|9�%�燾
B!�p�_��7��j�6�TJ�env����B^3��=s�5C�"Z���������%�7��&�d�f��	�
���K��D6�{�k���X�`,�:���.1�;s���D�j��ݞ�q��<���BV4�B�Lc;�~lىk�*)�d�u�J(b	�+YJ�R�&4H��A�k|O����M�a1�!	�*$by�)Q�J��Yhl[l	Z2�Vc���6�W�Q�Gp�A|j&I[*���/#�t}F�g��Z��
Q2q*	C{�^$FE5�{�R@�
'��|��ȸncn%.�)�(�����þ�a�Y�F��!�t;������!�z:O�Z��q��!�b�cr��?�>����g�I�q�hr��\����a"�|����?B!��������Uy����l6[��j���mS�Cm)O���V�Ɗ��Jw��ܻ����>�ñ<�m�p,d�>��]_wl���8G'��b`�����k�a�����{mSOl^(BuC��]\K���D�����S7��h��*C���.�!gL>_���A��F�w��9�D�bB�J��*��Bڒc3|q��l�u[2X�������f�v�p��.2��S�S�kٖ�jӻ_��9؈X�kibC�F�2�E/�������;#��ޤ�O�hl��O:T��X��]�/�E��Jl�]��'�垛'N���p{��.�����L�R��m�*�@U�D┛�>84���GҘ�˴vBYi?K�8!�����x��?�����O���o��z��/�d�C=��������!��88W()�d6K녢�a�-X3�_7�c����p0V�P���R�{� �{�3���r�Di���F�>	^�n��xm�L�䠬f�@u_�����^�7m�~\�5EUm�=C�̃��;=��%͎϶YZS�4+���1��L��E,�v�BBY���N!$Qr����1)�`��	<u|KSǰ��'3��	vF�t`{BW̒W)��]$b��+�	���n{:{�A��v-Jx]����M8͡*8�����G�7C�5��x;C�h�8󛏍9]=_��L4���^_!���{�2��LM��k[C�J�
����!C{@��T޴���]gl׉UAQJjj�;��\���q�Q����vB!�BY)8&�7��3���{9�w�������4���8z��`���9���?����BV�z���q\1�C~�H�^(�ZV'�ޛ���v�n���B_�Ц^h_+���	�7�6�����z^�Ɍ�*�L�Y�ݩaH�x�J�r�����Ƅ�����͌���tufv������C�t�Cq0V�nhalW��U�DmZ���2����3�4&6��s���!��L!��B�ƞӹ�Aov3�٘�ƞY̜9^IiH��+���+`iīHF���� �\KhxoM��Lī$�J�;�bV��v��F@ਜ਼�K�Q��1�D��2'l���,���.�W{UQ�g�ƈ�ebS�^y]�Wؽ׆fv]�I���]��`bh�R�T��v���I[���j|�hg�0��B!�BV2�|o��O�C��7_��UC����_��O�BY��;�/)�n�������?7��ct��fw�u"�X���XI�ܓ4�k�)�p,�4Kb|��냺ڠ�o��wN���l����cb0���~=q=0�@,��=0�& +JQW+���	�2������K%�UIhl�����k���v��a�����<:>����~���3�B	C�;!����T~r�A��H?֏��ի�Ν���d2Y��}���uaʻ-������n*b9$ep׉Y��ꍱ�]�X�{�7���<�T,2����S�D�Jm�H`=��1V6��05��j�6�*1�='ip�nl��BT�2�{��8�v]�H��R�4��f3���G���#Lk'�B!���1�����������\�t3_��Q�z�C �BV:�KEܵ׹�Ήո|"����X\X��b���@]]P[7ݽF���XqC���Z�c	�M±t�º�����6hRT���z�x��-�h�g$]�F�0,�q��P=Ѡ^(�K����u3C���X��v_���v�nϽ}��ۈG���N���\B�C�;!���r|���g����tmO]���c��s>����=p֙�e�+:�E���=lx��M�+�������,�����{��%}J1�+V��6�������X�3Ë��ϗ����<{q�[�)<_7^g^�iE�ڽi����4�!��]��P��瀹]jl7��+��$�di�θщI�(��;�
ȝv�nL[ �B!��<犝8��?Z�{>yQ�����۴I�́S����7B!�Ϟ���B&�Wn����Y̞=�\.�4��5�[�C�B�N�㻿�'���[���e���u�޸>hXԙ����Ў�|
�Aͩ)FC����m°��e���������D�qk��5����A#�8˭�k�>C���]�ebl�����58Q���;�|�X?$���wB!��#'��#���\�9�u�)�?{&�� ��gK��䨋X�{J%b,�x�>��w0���c��2!+�}�-�iڼ��pl��Peon����U�iV��e�AqI�f|_k3�tF��9I��q��Sz��+PM�r#�IR�L�2��Fv�UOiS�C�H��}��G�9�E)B!�B!z�$���J�|���&��x��?��� �B��B)����q�1>��l �g0;=m����n�h�0��(�=x��
�ꄭHvW���x���*�{���*k�A�g�iM�δn:����x�?.��A�`a�@��u̍���i_�v�@,�0dj�E�DO�дVh\O���C��XX��<���}�ѝ�CB!v��N!d�Y(����~������W�$L_8�s��@��3��|	2�{�6��	�2�{c�_��wHB��1�{���4��{�i�XFm�>����k|�%�vEfN��4����6���BT���>��mL�"A�onOX��U�v���'����3ۏ�����)B!�B!v8&�_�����w�Ͼb��������� �B�S�Eܵ׹Ǯ��x�x��cX\X0�jB�P�%2��j��ڢU�0Z-���NhZ��_���>�z����f�h75�{��R��x�:m�]V}V�������^(�������c��~B3��.�%}R{�ڡ��.2�g2iLl�޹~<pĭ@!�D�wB!mž�|�pD���5���W���u��(�]`z�	X"C�Ѷ�³�ɽ��nfh��٣XqD*��]3&t]m�ߋڂ�y�8o{P3�2n�	
?Q���L�CO�hh��MƘ�EcTb��.6�{�%�(U=�)�e-T�"S�̮��&���|�����0��p�S�W��vB!�B!�XX��������ϼ|;:����wp�� �B���3��B_v��1����={�R�Ig��P,U���쮫z�}ie�P`v��e��t8V�s�ڠ��%m�z�uH���g��]�I�`���	������%;����E3����b�ñԻ=G�!
��5Co�X,T��kq"?��<�������!!�����N!�mqūLj#._����,LG.�'5$`r���Hh���f���=$b�c�X|Xܒ�Y�8۴��f���Mfz�{��k��Dka*e=�:JA8Z%<Iƕ$}Z㺤-��`"@��L�D3�W?S!J6޿e�����F��%7��(YH�Ҙ��BV��qc��#%�NAQ�B!�BH�8&�_z����^����-_=~�4>u�C �BH|�%|㠣Gb��"\�1���fΞ���LC�du����Ʋ�	Znld%���Y٦�Z�a�j�"��M�b����z�st�D��i]QSS��ez��%����P,��]���~���]bv^5�����#��^�	!�$O�*��BV�����@��Vov3�٘ņ��p�x�[:m`vX*K�������^,^5�MM�^�ɤ/h���9�����鬒�#�v�O �Ȅ-�8� �K�z�|eo�`�#듭ob^�]�R����1���Yڂ+DU�eb��ܮ�:0�P%2�������R8���:��B!��9{~�f06��k���s�!�4������A!���b	�T��A���5�W�)̝���
�I�2�{û�v(�JL��Z�����p��k��5CemPV+Ԙ�C�:��F(��ψZS����(�X���<�qB�Lj�&uBU_��<Klb7���&�X6;=��&5D�`,Q�0��chx���w5�?�������"!��fA�{��ߛ�P_z����`_������\�Hta1�Ky��|a@Yٔ��JRC/������13u�&�(�+�uPĊ�����,���6��U�2�L�T}n����cԆwXlU�:Gi�{-����D&Ř�X���s\S���FOQ�=cJ�f3��O%>����T"��>lf�R��F���.3�Wۋ�k�06��S21�����TE��S�1�jz'���4�Q�"�B�
���<��g��C����}���9�w������ �B!���L�q�^�j6����\8�s3�d�Z�{��.	Ȓ��m�����^�Jk���wY8����6���-x-��֢�d����΍�U�1X�3�dV����nږLQ����ܓ�2����fv�`,���P������3Y�;ꦴ3���dʯ��z0��S��ɦ�ߓ��|�r�/������Bd����8�q׍b��1l����ym�m�`Fz�ۓ1Zk~)���05���.�������=>�ss� ���¹���Ϲ���(�\��dzsS'+oڼ��:c{��+`��eFw~�{��4�7D�ƽJ�r�&bAK$d,��JT+�u�{Y��=4�:�z�c{��Z2n����Q���T�k��LV�ڃFv�����AA�.D�M�k� ����*��=dbטۇFW!�7���bߡ<��&E)B!��\���}����u�n��3���{+��i7>x�����1��=GςB!��Oʇs���ۀ�GQ�;���B�d&wI@���nS+L+j��0,Q8V��Nh��uAXfAY��m_��&��v��}��,��RT���P��b3��k3��OnX����5E(�d��j{�P,�Z�i��6kphZ���������<!�S��V��[�c�Xճ�xxǇ�*;�:�&��?���-bf~	'��^��Ss8vv�N����J�5i4�7�գ�t�.�:�'n�EkG1T��q��V��I�'B�S�������#�ǁӘ[�BH��$5�S1��c��"\�!���pa����aKez�km�fw��]ix�	RRӻG��Z~�J�.��4����"aKvW�j���� �Ldb�����zc{�J*@�Ũ��]����mJjl�'-D1�+�T�vs��q\��N�p�kf�kFB!���ǧ*!�����B!�BH��ȕ�t�j-vMfp�x��Ә�'��-1�'�<���~�{�>TL��B�cnxW��eF��L�Q�u}��&��FUC�jf�5�vhcf�^�r����ݿvx��`��[7����:�A�0r�0B0V0�}`p��I��Ã�r�g9��Y?$��?��4��i�n��;7���k� [~�51�_9�����E�?y������O��Cgq��,H2��� ��\�s��x��x-6�-�������Z[9�L{�M�{�����x���c����犸�`�|Ջ��<mcz/`~�$r��\��������e#\)M�A㻯-�Ԡ2�;��-��Zntw��}ɧ.�ڣ��M�4�f��EmI	Vb�r%ik���E&v�}H|��I�>1�#^I��Q���hWR���:�j�bj��X
�:��"!�B!�B!��nd��B�p�Vc�u�t����fΝ���D�0��=�V3�7���&�c�j�~3��6(�O>�=ʽM�M�9�z`�9I�
u�Qj����Ѽrj�mk��6QV��.6�B��E�n�I��M�����A~`5;׃=�r����޾���B�_�;׏ᚋ���'��%[&�ͤ��c�ɦq�Ʊ��]Ti;7������>v��>Y�'Ѡ�="�ϸd#�}�f<m���?�v�y��~���O��B���1|���+�<��M���f����ރ��^�e���l蹀�󧰰� �D���he*V����߰�Ml�S����CFw�hezV]G���n;&)L�,՘VT�s�O�Yeh�Nac�8�AlbW'���Cfw�%�d��&���0����(��;[�3��K������#�B!�B!���88](��*l^5��Lѷ4���)��]V#���5���FwQ�P��r�8ؘ�eFwy�����F���]�n��J���e�Q녪>��=x���fv���Ԏ�Y=hf��	C�C} ��NhSC4Ik�������\���f����	!�=q~�:��_�Y�n���~�+cC}���͕��}���S���W<���/��C���������W_�k/^߶�v��=��+�V���\������cG��2!��Y̗�f�Lj3��&���y�,Ma��tE�Ɉ�(���R��1��S��	�"1Kjl�E�;�yU�
l/4�7�+W!�J�fs	Y�>յm�I�͘����U�Lĩ`[T3�x����8�(QJgb��GQ6���M�Q*�!2�����A�����|?�?Z��ch/�B!�B!�B!���|�p���.�(a�0��sN�{�W+�d���~��=��=X?T�E�w��]w ^�{�Ψ^(���񪳹�=ʽ�M�n��
�������+*���X�Zb��$KQGT��XI��uDU8�&���M`6�
��u�\s;!��/'�*��7]�kW��p^{9	���k/x
9xw|�𾘣�C������Q�F��o#=x�5�+��G������W<�oBȊ�P~S���|�p�ƱfhOY��dzΝ��RQiv�z�L�*�*���4�*Y���^�����yϦ}b��:(0�����6��L��^ӹ�^�'�V���mz#�(�]-Fy�.�ٽ"Z}�A�)	�{��+:9��Iu��ڇW�B�w�g��Jǝ��!�B!�B!���5���zGq����. 7��	:���n��nW+Tރ�((+�����ʕE}���n�e[lg�{Ts��OdX�]����EuD��]V��{�EE�Pdh������^�4�G�
�S{OoW�ƙ��;Z��)�kƝ�	!��D}�%��s�n�;��w��t���)�&+�{�Sq��������S3 bhpW�y�0^���xo���p��1��%W�-�
�� >��Ǹ!dEqj��{�9W���n�e��:����i,�ϋ��&"�+,Y
X�fw����R��bUX��o\��^iX@<Ѫ:_צ���ٴ��%GC3*)�K�6ս͵�,j��nh��Ae��(���b�F�j��=���
��'ë&1��C'S8q��ω���;��B!�B!�B!�dn��	:�Lj�o'���iy����R��^/����~ӻ�(2��{�x��r��nۧ��c���hr�5��k��uD}Qox����=u@O�0\W��Ek��M�jC���!c���><2���$����cy�O9_9��B:���,n�|3^q��e�0����,^��x�;��ޓ��w�໏�xr�����~�<���Za!��e��ċ�������o<���EB�Jb!�w$���)�X�K��T���y�N�Ep{Ba��J�
W&��M���]D�@JCX�
��������
R���8�uc��>8^5.ܯc���jI3��l7����'��Į>����u��&4�������dr��^*����(Jc8t��!��(b�!�B!�B!��8����NUt{��=�f����N���Y^?T�	E���
�ҙ�m녺Zbr�j��>���qofn�^�c���uA�����v���j�g�Za�����nXO���02>���*��dG��;<s�gBHg�ߛ�Kj'^y�0:؋���⪝k+Ǐ�Ň��#ܷ�H�=l�Ư�t	�u٦��� *�=���]x�5�+� |��af>BYi�J)��5���1\�6�-9���a��4���-�"V*lv��X�"�0�]��0�#�'4�{���
V���н�����o��)�_{��[��6��ɡ��c�}zs{p��ϟ�P���E'wl��afكb����1���-�p��t�Ts{P��R!J�_KX���l8�A<|*�c��t�#�B!�B!�BZ�w'�ޭx�,��/ �0;3c��nb|�mM�~�{�@�@�PT�E)�vY�구.������}��ă�*-�1��R�킱Bf��C�aX�Zb����n['�bnW�ڣ�bUR�GGP����><x���s���=!���ɦ+)�y�16ԇ�Γ�L�}ox>p�t�#���thpGuk�W�pq����!�z2x�3�����"|���/|w
E�@Y��犸�H����Ć'�IcM���Oaaa!$b�j��R�r�����njt�U���av���'j������@�L[���^�n��Za����?V&h����{��]|��j��5m!�/@����$�uƚ�m��&"�N��m'�����c�ό���,=�C���b!�B!�B!��.�-���CNM�|�ƚ��x�Dk��͜�
e!X���, +n V4��:ˬV(	��d낦aX"�{cL�O��oS��Z���X��`��?.z0���kV����cIk��:���hr���I�ۍ�6�X�=�P��N��a��B��랴o��˱qb��S���_�����c��7�� Ǧ�RY�w���چ7?�)X�¶6�ed�����W_�����%B!����ί�Lj#��&��9�g0;=U~#�lQ�7���Fw�uRF���U@�
���Mg�P�B�=`x��i�aa˗����}��{Y[m��R)�ar#{h����+�"Su���~�5���New��⓻���.����o��m��Q�^1����v�����02:�|�(����y�ܿ'G�JR�$�B!�B!�BH3��
��غ*�'���
�?{��Vy���-Y�{e/�w	a��B��R�h���Bi��Z��(�m)�z[n�C�-���=BȀ �vl�{H���#ǉlK�lI�����p�y�<r�ǒ�<_�N��6���=R���s�0Q�=��a*k�Z��Za�����q��kzI�����>������m}�������-Y5���K-���| Űz��'X?���3��(�.=�S)�����@�-�5��X[j��U���84�.p�7VΗ��}[2�LL,����Vy��-����p/�ˑkV.�����_��/>F��~������� @����M5AeS��b6�ej�Y�z"∶K{�>	:�޻&�����8N|��P��米�]�w�1�%'�R�K\�=Q�=�~��{�?�y��TnK]|��m-�<����=ں��S��O4%��
��������CކZ�=��dS_A�>�������J��}A�l��Hî�|        ;��ʦ��<N�XdTN��M���(C?a���Á�jtҚ��WO~����6~�Y�Gؽ�}
����#�<̞��`*wMdOt�h���������� �I��Y?�c=�`�}��}�r�����h
��z�!�ܹ�yd��&�C�ѭ( LF��\2I�|�L�[M��X-&�`�4�̜��'ߕ�>���d���_W-�,�8Sl~PC}O�7V�O,��?�����Z  ����XR6��.&�(��o��ިx��k��`GG�2���{'�'��5	5�
��{�<�u�����Uj�/���}�u�%>N~��(N�;�S{!ѭ�g��	O�	N{�;R
��?�`:�:�P{�ɦ��u������6U�Ď�;5�`{J����d�	���"ǭ�s�&`���#���hg2
       �C�?$���ȍQ���i͗�E&)w��i����غJ°{_A�T�x��t�v��N��=�x}��5Ã�ۺ_\�=�5������L"�D�n���7A��h������{��P(+>��|1q��ۺ� ��Z�&�Ǉ�5X;LV���46���(��ФU���E2�,W08�
\򳋎��^�&w��}	��j�#*���ɷV-�%SKCW�˭_X&ϼ�]���z�� �\8j����ʦ�uާ�e�7,NiK������L,�O\%���#���D�P'�Tڄ��;�Mb%�wݯ�4�m}8��<���a����6$���&	��ݒ�-�� nB�`{��	���N��C뉂�]������M�ɩ�����ړLJu�7~S?�����䖪6�l�I���;D�       ���-���t���nv��"��r��n����ؚC�Za�uB��c��^�U�]��m��cG���ܧP$+�~��$X/�uҽhV���}��ِ� V�A϶�����>
`�O� �ą���[G�8��놩Vp�V�s�p����k���ϑ�啈�#�|��:$~���[����+�R�Z��sg.�(&�-��)[+�P7b��w�,��&Ў�"�b�x�>:O~���ew]�  RV�a�e_P��3���K��$��)��l�����@J!�>����hKGeU*�}�':Nm����7$������{�(ڐ@*�U�>��I��G�8?\Ov�;��T'���5	��]�ɪ�ǉ�����s�N�9s�M�٭i3�5a	�G�w��        }S+��[�wcg.���2��$��a��[���A�@�����궦�O[:6�@�����?q��T���w�jH�=�h�u�h�ۺ�F��|��b*{=����-�:a��Þ��Yr�y�3�dO�I6XCT��`���X��5�d�a����"������~ ��������K��:L�|���/�H���^�󫟑�=����q�  goKX��#�=�+�W+4�XOD◈�EZ[�c���Ǉ��	��tO%���p[϶����{����J������$>,��~��{��֨��gx=���SZ'���s�)Q�`&�������or����
��O@�:��l���A���f�؝�Xe���E6�F����rO��        ����n�wu�5��\�\s@��Vikn��a�8V�����5О��a����W[l�y�Gہ����zvo�}��:LL)���`K��R*����~`1A[*k��Ǚ\7Li1��a�}|��۝.�i����&�l��HxE� �lS�s���K�4/G��Q�8u���/?�m��r(:��96�\w��tZ� �����s���{~���ܦ�A; ��#"kBʦ�Y��@J��2�k�B�Z�U|�M
�zOd%���U���ڵ��0� {���P�Γ���x�~�0�޳-Qp=�q�!���2A��-��3Ğ`"�@���`{�I���(�{�r{$bsKc�&�Չ��H]׳�D        Ȍ�MaeS�L��rZs���:;�c�����=��X���n8��{϶���Ֆh�_[��Άnߓ�`|�����H�z��5%.���8�uî�@�S9J�=�:b�������b����Εc��̲�6*�{��� �I����g���$H��sF���\��W���M5�l���㐛�_�42G�E���ɘ"���ț� h�{�wwl+u�d�� ֐�"��I{[���='�MZ�0qeL�&C�':�~0�}���>���ݓ��S���٦U����DP݂��ݖ �?��m�ǤTgev�8\�Z��.V�i3ʦڰt4v=/��'\       ������I-�U"��L�X:�j_K��B݋cůfr�0հ{_����6���:a���E�k�}���n��-��YOLV+�zb� {�uD�8�^��s�>h��D*k�����g��X O}����r�����}�P��^�\nx�5ٰc�Jɀ��R���eR��㘙���m����� ���л*'��9Jd|��@���EZ[Z�OX�q�k�*���@'�DR
��w<�}m��'k�z�dP��j��| !�T���4���V�9ի��`{l��"��Dm.iYeg�ȶ���뺞��PY        7��!eS��J�	�cE��h�֖��k����ɂ�����ZO�*�ߞ�8�����O�8�y��D��_�k�];��8پ�x0����!�!�8V�:a�`{���0�ͮVf�H؜s`���D뺾g���/f�Q��j��0o� ;<9V��EG�-��)/n�#��C.�>ut������
�k�������w�Ij�} Ȭ_$�uR��c+��f)���i�9�_{�t�}�'�����$U�aw��m=�Ed����z':O֖�m��k�j0���㡆�S��u/}OLI���&�������X�bW���M�}&���ڦ��:��       ���{q,{l�u˄\Á�Xa_����ű$y�} �CY3Lp�/�>�uC-���\3T�s�0�x�놉�h�'��k]1ɚa�0{4fw�s�Ø#u�|T�����îc�@*,f����r��rAvY���9G��O�#ϼ�]�T�}��b��%����?�����`�/j
þP$��D[B�H�����$�٘k1�s�c��b�x�E^�2��wc��򋋏�o�ϋR��. ��j��;���g���+��:L2�m�gT���X�>	�����&�?ލ�&�zNf�:1�j�]$��{|{W[��z�w�$��S�$���b��g[*�Pݎ{���%���'�"�BOj���p����X�!`�]MQٵ/�ܧ��BUv         U�/,��M�Y�e-�q�F)sE�m
�9엠�E|����k�n�a�u�������s�輿v-�c�0�x�����}�t�0ٕ��%v�#��9�1�]2:�)l��v�lkI[���5]� ��`(Ԝ�.X*s'�p���Ե�C�M�F_G�)��i���Ñhk8m����f��e2��V��e1�^�-�؛�t�-����Q�
�Y�@lf�<��'2��$x
N.���[*V�I�����^Ӳs_�����ۑp䅊����`����~��B����1N�uA�ǱpR��Xy���Qy�S~��c��������@��	�F���ؙ�V��r�%2!�$Ŏ�䘂b��%�K{kKlr�8�J=��Ez��y�&2��+�*2�r{�dRIo�?����q���T�DS*ǉ&�����Y	'��`��s�ɖ#a�MڣV��ewsT������5��_�  @���f)�Zēc��(&���:BQ�D��-${�����\�IJs-��1��j�����3��QeklI�2F[����$ϥ���ƨIlfe���1�T�hD���J��+t'�-!c��5,{��z^G �ε"��F��3��3Gl�(�����r�Ar�!�E��h�֖�ߓ�5\7�-�%�>\��q�%kK����~��d�d�4���a?k�Z�Jh�����՝��i[��g��ui�uug�� Zʱ��'%3����^��TYߺ��5�v[G�s�����W5��k��iv����eq�˶hl�kJi��":��
r�isc��~i�g�D�}��B�Ig�v�:��{��4�^nl������?Pq�_�=��QC��=��:֖�6*7�h��q��!�}��ƽ�Km�O  �C�?"�Vu��_M����%ϡNj�@9��C␀D���oo�`G��dS�Ė���`�I���$�K����Ie/7qߖ�8�y��$�H��z��������������6��<��T�ۺ&�ԉOu��bWC�v�P~=m���%*����O*� p�Pm�Rf��csd��L(��M��/4�4?����]>yw[��k
�cb�Mf�ct�C&���a;?uя_X�V���>ٰ�M*�z2I���9�������:�#�u��=,Uu�����]�2FuC}�W_;g��|U_S���4M���M���{�{}Mc  �pT>�+[W�=�9,E21�(��%��(�߄|���;|Ov%h��&���*�5��{W[�}�����o�;��O��DfВ��`O�n�3���z�t_7�/�>�`{��]�="6{�؝959�C,�4Iu��*����� �f��|�R݅�wֶ�+����:�hln��m�:w������5[��������;:<�麸�k?~��	n�~&�.9y��ay�Oe���i��c?,6���_�>�ll�����:��]�bo&�����\w���Jr�S�sOS�rH�����O/:J���il� �����Ķ����\)r�b��|GD����s4(��_:�>e�Ht�>./�W���z�w{�}?Ǳ]��dmɨ��J
�&��(�j�=�C��>���{lf�Y����v�m������7J�Zͬ9,ц��� �P�Vi?~�W���B����2�"�S\���/VV���MM���V	�S��s;L�9����<�^�8��X0����B�to����Y^��"� �٠V����in)e�Ʈ��h�+�]��\������8y��J��剽�{���������}�8���1ڬ�׷Į�  0��������<b5��:MR�4H�-"nSPLa���������h8�OR+Y�=��¤�����%�'�s�4+�/�uÞ�IlOe��W��}��)����Y�]=�Z-bw�%juJG�� V�2l�7���������D ���(7��T�N(=��������-���ʵ�g��|�9o*;u�����]��o���\<�<o\�v���|���������hX�$�*p�-,�=����-��{��>W�����Vn�b�{��L�����<{t��{�'ϵ[��m[�V�gG�տ{A:�\� U�m��v�y��~�*O���(�Y��\�������K$�!Ae����'��WzIp��T�����R�}�yl�����N��z�������;����j?p[�@��sױ�b��!&�U���$�|}���R���ְ4w��rS��/8�* 0y�r��|9z�[L&��Q��6���,-�g�i�g�7I��[F�68cQ�,����1��Z�ybi����ѿ���|�3!�e��ϗ�f���h2���m͑����(c���{Fx̲R���t�����������m͑���{=�   ��@HdgSXٺZ�P�+�Y���;D�֨�L�� |���������',��J�]�n�(����}�ǵ8��(�������
�S�'YK�3ܞ�PVך�2 �*�&�C"&���f�M��Xu��T�F$ج��nuv	��ިos�Y�P�R�կC-D�~[��5Ϳ
O���sO�śF�E���7��7��R�����
֌*pٳ�5�W��֪����7>�h�nMۀ�'�*?��H�:mY�j�}��?����֋o�fm��؍��|D�=����<���w��c\���M�'7�s�\��W� �@~�W�O�{�~��Z�ڿu�s� � n���AxsD,�Nx��	H4�p�#V�A�Iz�c��G���e{�����v���Q��rOi��B
�L&�����&��l����%(Fi��C�%��ף�Ҕ(�^  #��(r��\�ܑb#4�2���y��	s�����{���a2�y^9{I�8l��r���FY�4_N�㕇^��De�/-���^}�s�
�$�u���\����z�_{d��-��T����9�PN��'���1
  yj�}[}H�uk�*�匝yl)v�(� KT즰X�1FC	$���U�Pq��*���|[l�ߓ����?���n8���Ű��\W���v1[�b4�$b4(���a�}��T�FzT`�" 7~f�?wL�?���O�}�qe�7_���c�]y�ewAEE�ֱO�p昂oL,��$�9��?�X������Q��ap���S����ml��q���v�~お��2��|ٚ��������R�����KNp;�_a^2�T.��l՞bR  U�IDAT��o �d|eKtKׄ�Aꤗ�n��(9��8,"sT����e�I�e� !�F�$K(�����Z�H��S�����&��'�dT��������:p�ߍ��4��h4vN"){��"�Y��D&�o�l��F	��V��HkG$Zo�+�KT��}5��  @jFX��2J�cpJ����e���fy`]-^5V�(c�D&�f�xʰ�V����9|�K��g���Y�֒���JeBq���w���1:�S�S�h{��j�<O�e2�����R�Π��9��?�U�/�{=  �ԫ7w����V��-�@�Z +_�ԵA�%*9��������DC!	���!	�u���������.}ȒԊb%]74 ��d�0��^!�~�{����:6�Lb�Z�d���d��5F	�Y:�Fi�%h�F�{U׶�J�	sr� ����c���Ӳ���pD���v��*�z�k2�TT�	������=uݬ1��5�����בc3��,�+�\'u-�'�<,�W��#��f�q����������W��,�؏.?}��;��w?4il^ޣGL+�k4d6�f����Y��� `��&��O���o��}��GtZ�b7D-:�Ĩ�=�ay�r`6E�}T�qT��m2t_ 7�)n�)�-6�Y����j#Q����n�	D�����*����JiD%��զ�Պ��`������9��*  ��Q������J�vM;�#�K�r��{��! ���r�)%�"�&Nr�-珑_>U%�j:C�h�S.;����9b�+�A�ە1�s��ZX2�%_9����9r�2FK����=u�Q  ��t�J�._ �}��f6����wYE&�r7�)[�Se%,�HH�:Z4��Q#�	c�C��D"j�,�
ս��������MZ+yQ,��X�hP`�cՍfuo���iPW,1�%��R�`E�W���z�f���kT�:±J��Q F��e�r��Yy�U���}Z{ፗ�~R�����[��-����/��5��^�5�kE�T��$V�=���.�~��1r���v�U��f͏�X��Bn���O�ݼ�y��œJ�W�vf��q�|�to�l�^�>  ��I�@H�_��J�<  �0s�\���B1�mהZ	��猒�=Q%[��Ou=:z�;�T/�	���r������+뷷	�e�^��\��"?8g���齲aG�`�N��/W�{������u��'���J�   @��Ԇ�R�����/������j�� j&M-������n�Rh3�����u����{��tDcű�����I�u @������%b5g��Ac[G��-{�k߾��+�#���k/>�o�����Z\�d�S��/��2[~��2�����|s�>f�����w��{��Na7^��V�����J=zF��Sf^����?�X.���#$     `�:��9�<Az8�&��Y���G+	�����Y��3Jc���F�}0N]�+������j��o�Q&�=UE�}��X�'�[V H��(�]].?}�R6�&�  �G�Օ�$���<  �u���Ii^NF����n���.?}��n���n��w=~�Q�K�+�w�2�ث�LR~�6��6w��(מ}xF?	�����͵����ޖ�������P��7c�K&wT�K�<m���ѷ     O'��n� 5�����r��{dgm� uK��	�g��d��N+�}�
��l�[�=�p{�Y����2���=|Xh����%ܞ�؇����?��5��    ��X�t�,>�4c�����~�o�{��W�q�e��x�/~f����O)���ǽ���yW�T7�Ȱ	�_r�,�T���cE�QymK���G���U����Z�=|����>����	�c2�'�+on�+�����B     @w�'8��	2#�j�Uɾ��]��ZX*&����	�g�U�,S��N�k檍��6�.�2F3F_}�2F��S����#~���Lqؔ����1��c�    ��_⑋O�����^��{ss���\���0�_��^�����{��Q�ح�u;mf���Er�}/H$*�5,��'˪��3�X���?�����/^u��`��**��k[���gf�>ݘ�����>_�o�'�-T�    `�(p�	efA��"��Dn{�J�:�|���(W�R�,��qٍ����Ç�H8� ��n��~V�F�h&ysLr�2Foyd��q�@}����hf�Lrթ%r�c��Q     �1f�A�]�H�fcFﭏ����޲�ƫW7���O�􆻞�˱3�-�ͱ���f�+�5˦��/m��}�]�!���yY$ml�<�ޮ�o�l՟RQaPK��q��<����/�Ŕ��s;,r効r�C�     .�l��o��� 1�r�q�<�nC� �?S,E^�O��&����������]|b�x��0}�CV,̕���kg���IŒ��>f�͑��y���6	     @&�=�0�\����zus���M'-؟U�n��̧����,�U���b�#ݏw��3�M�RY�&z��Ys�	U�J���4���oϩ#����Kg|7t��'����9�58v�(Y6�\^�\)     @ߖNu��1i�_C>T���q���ަ�v(�4�s�H���y�ڇ�R��6{\�,��ͦ�K
�Տ�d_sP�ۢI����=k���[ۤ�5$      �4��%7-��F��v���z���[������}r�/�8}t~A:�f1�7�\ ߺ�E]^-X��	%�X	�t�^��{������$t�WV���������aI�'�v�\y��j�X�    @�,f��wLZ�Ր��$k�̗���t�^��e�ʐH�l2�9G���O�tgT���
��jQ��Q�g�=�W���8���a3��er�?�      ���r�X-齒_(�����^t����n����_=31o�;�hT:k��"�̜1���]�7��_v�l1ӻ���-���=�n���M�>�xɪ?D�z��E��Lc%�"�C�9z�<��     ��Y�s�zji�8n�G�|�^�[)��I.]`d�.[d������LuIYcT�8�%��j�����;j�[
=A�9�-��V'�MTq     �qԌr�?�(���Vn�ݝ�n�_�U�6�]��D���m����t>�%'ϖ�7W�(�nW!�M/�E�K�������[�w�U��Su�e�����5+N�=�����ч����.Ս�     �E�Gp��\�>��OY�'��Op���z�V�?��\��3T�w��<�>���ϓ{�Y#��ܮX�/����i�kWl     �`6�+'�J��<�ޮ'�s��_�䑊��ѿxx��j�6�<ד��)��uY�Z�w�j�%�M�Ks{ ���=�n���Wr�WV�2灿���`�w�i�Ƴ�l�/�0Sn��     �e�8']u昙y��:	���qE6�Xb����.q�k���L.�Ǫ�C?��?��V|^GU�F9�<��z=Y6�->�O!�(     �֙K&��BWZ�ō��\��g
��k��{�|��f�<������(�_��&��}����8o��.H�K �g��~ɍ_=�i��|�����?�u��Z������1���[dgm�      �8j�[�/.�Q�ˑw?m0F��d2��).���fcT���,��71�:jz�
Ba�6�,���>j      �8�f��1S��o}\��f�IG��Uۿ{�Cǜ�`ҫ�.�)���V��������f�A�_>-���n��?U|���Cr�+>����-\8�xR:�W/���g�M�.     @�F����Q+dp�x
cT�'��^���魆��9��{L���:F	�     -�Z:Ir�����}�����/�����=���W�����^�r��{�FcZ�����/}$Ս�����p���o�m�;�����h�}���
�;���t���r_��5,|    �J���3s�C R�5K��"Пi�X%�p8*#YY�Ur�i)��!�>�+��CT���ig���e��@���1
     ��Vo?{ٔ������n�:��k���L-���3k��3��t�o6uVq��S��*�Nʭ9rr���iln�ްL��[����p��:b�c6���FeP�}���co     Ⱦ�	Q�U��,�^��4e$�>�1�WV�A&���J��d�G���c5����j:d$�6�1�W���ʷ�      �)ǉ''-��c��`ϝ7^��Y�f^���(�^W9{|Aq:�?y�X���7ICk��Hup_2�L����w0��l�}�O�:k�@S?����s��?~v������	s�����$��}     �ktA�&:1t����H��)LߥT1t�k�H��)`����B���:�o��(w     0T�W�� �[�?��O�B��G֮O����U�� ߭�e����x���ߛ%�tp?{Y�~X^�p�k7}����E۶_�Z��iS�rs��[����#&���(      ���-�*ϳ�>.�=�Q}+��C2�Q}+g�2Fu��Q     ��e3FIY�3-}7��#�ZO�ŭ_[��{�S�^�h�7����%��O/~$�`X�I7�1�.�3�(-}�k��>�ٶR�6��w=v��f�Q��OY8^~��&	E�     ���C�Mϊ�|
�<zV�e��\�W7�&Y��7�(     ���'���W���W��K�6߽茫'<���3��jݷ7�*G�(���g�[��Y���(Cz�~es��~���5�����O�=��7��^v��}�lr��rya�     ��j��vh����x��nM�$�0��7;���Q�c�    ��*�ˑy�S�zkUS��iW	�n�u�N)���b6i���E�	���&��8lZ�޼���{��N��w�=�roe�7G�S�#�    @���<�T=#�<ƨ�1F�1�s�g|Dlf^G�,��Q     0D+Mc*R�yo[�y7V"�������?�����9z��}ϝP$c�ܲ��E�E�%SKc%��F�]�	2�o�f����.���hJ���R��     �y&����H�h$��g|HF�<�6�ǨQ�뛌#�9�;3�!     `�\�	��S�����n�t�_�}�o����*w*w?g����&�]ܗ���~7l���K�m�\���wA�ǡ��R�ԏ�9J�              @�f�-�b�C�~C�����r� �~���5����玝5�D��>n��p�YLr��Ҵ��aU㵂�����ۧ�ᯏ�8o�Z��>v6w              ��:vVz
R��i�֛.?�eA�U5/j��r�̚^�ot�K&����U��Y�/>�TV�M;�ko�l�YѼ/piC�M�ˮ�e�O��R��               ��`9zf���F�Q����JAV��������o/;k�QZ�}�2^Fn�}JIZ��pO�����zUc��<s��1�iٯQy�=\3g�               �K�R�qh���u�n���
�foSۗ���Gv���E���_�$�p_���{e}k����K�U����E"����q'�              0 �KOA�O�#Ȫ�/[�u��޶`R�-��\�+n�Ե�%Ӳp�X�b���ټ��?����kk������WP�e�'��Ѡ^�B               Џ��4�S���1��n羦{L*�E�>��B���BQ���M,Ҽ�H4*��?����5��-�t;,�O�|T�(               H�b6ʌ�����yW���\zrP�u��c~^�⿩�m7i���	E#/�>sl��}~�����+׼.�����큫=9V����W@�              ��F��B�Z�����.�s���������勵�w�X�?��,ܵ�Ko�izB�W�m�ؿ>Z<�d����W(����                �t��Q����5dvu����se���}�*pI��&��IY�y�Mk��mw	t����e�m�=K�              Nf�!s����}����x����H�Ӧi��c
��͕�IY�O.�ռϪ�����8�M����wF�ѫ��f}���:m�Ԗ�O�               '�˴���k�xJ�+������?�x���N.󎜀��R��}�i�X�;7_�f��^�)t۵�w|�G�o�               ��[�؛�i��pD�C�	t�������@�>'�x$ӲpO�_v_��]�YۺyL�{��}N*%�              �������������^]#Н����y�]�����Z�}t�K�>�Z��
t����we�i�}L�[               �X:�{�[��ҍW�\���7�I�>�\b6%�H�d-�^���Ls{ r�Uk7	t��C�Uv�j�gi�S               �Xin��}���o	t���W_�qi՟� R�uHe}�dJV�n�E�6m����"Э͵/�a�Z4�@HZ^t              e��nD_�V}k�ne�Y�]��>��騼]���+ЭG*��t�+��6��TǑ� �
               z(�uh�_4����u�j��(��Z�Y��٢�Y	��95�8��l�ZCk�nt��k՟�l��Y�:B              ���]vM��k�n�ֹ���F�Tv�ײ�|���?Y	��s�������ZS{�Ne�Y�]�ɱp              H��qfw_��I�k�`�?Z��qh���KV��4TpB�t�#ޫu��U��               ��qٵ&����]�RݱQ�>=9# ��[4�3,F.w�s�`�Q�>3��              ���i����m��p�]�k�T�����bҬO�H��n��	��k��D���b6
               ��������6��u��ŤY�֖��w_�p75�8��oW	t-kp���              �dNC�2
�
t��=9V��٤}���Ǔ,���!u��]�uZ����              0�Y����Qi�^{ Rv���d� uV�&�+�G�Qy��"�@ע�日03��              ������e8,݋D�a-�3G@�=�hڟ�`���ϭ�zU�@��&s��}B���              B!m�*�����dԬz�*�~,�%+�t�%;��ReG�]��F)к�P8*               �.�����l�t�n5���/0��4|"�d6��-�2�!�3�              0�� ��h���0�u�=
K&e%���4�S�6t�l2�jݧ?��X              �ґ׵��N��٭&����:2���J����C�>QC�@�,�W�>�1�               �����C5��Y�6�)G�kW���|�Q�﹪�= ����{�/�y�v�q�@לV�x����              �p��H�ۮY^�%O�k��2��l	�tT�v;m3��粕iݧ��              ���B�Z܋s�Tp�9�ըy�}DTp���׼O��:N�k��G���:b��               @o��>�P�]|3�f6\��?Ϲ�k���f��u��8ʤ�ܫ�%���`Ь���P�[�����<�ͤe�{�               ��#k��1-Wv�u*7�6I�>�6�K&e%�
Gd_�_����T��W�[g�X�<$�S�w�A�4�2��              0��#k�[�V��V�u��.J�����J��jp�ZL���,���	tǛc[�u���Tp              H�*Y�����N��wO�G��Z������ɤ�ܷ�m���5�3/��y!�K�^�QZ����I               �X:���=��
_d��4�s{M�D��Q��W7k�gi~���TTD���)׺�O�j?�               {�Z�#-C�E^��{w<|ԏ�X��@W�<��Z�������Z�=�Ie��V�o��"�@7"eO��vL4j�g(��ʋ.               �D;+pO��i��N痔w�]���u��(jޟ�ܫ�$��Ԙ���tX͆����*��#Ѝ|��\���T�aQC�               Hnke����\�r��|�g��+v{��W?�����?�O����)�ؾ,�uel��8��ܰ}�               �ow��i�Oд�)��q�z�Sqթ�/�
,߱����E��=�iY��6��<�>cL��u��˗�YWq�GN*��j��Ɲ�              ��}��N�>������r�_][�>O�>7ﮗP8"��Հ�;�e����Y�q�M����rx� �
\����`�              �SY�&u-~)p�5�w|��!��<vش1y�Z��1�HEV��|R-���Q���肜˅��.6:����V�{�              @����FN�7V�>���+S�����H�U��Gf�Q�~���F�!��_P6望�c4�W�o�7���}�\�|g��z��<�U�~��Z-               H�Ukp����q�nR?'Ȫ)e��h�g{GH6���UjXY뀻�j6���V9\+Ț	�����7�              �L��F�"F����_��슇��T���⷏^<���Ժ�w?��P8"ِ����[�ʅ��м��
WW��⊵�����7��8wb�8��m�e�v
�              ����U�=Nۢ�%�9����?yD�jAV�_xK:�}uK�dK��W5���[�ִ�B���r��F9�P�qFy�04����ō�Y�4              �p���4��f�/���"�͊
����??mt^����"Qyi���^ظG�?n���ΟXt��~�̥����A�\�cK�M(������`�               ``^�X)W��'F���-t;֏}���5mT��i(H����X��l�E�}݆�i	���X�xj�^*Ș�ŞߙMF��mjȻ��               ���/�?�����5�{���oV�[wS���!AF�p��g��_�����!��up�^�,�w���1����tZ��߻㉛tř�i��;�`��������ww�.y               ����;;�p_�u~�Ύ���iWQ5����4Too���H6�"���[��p�uڌ�s�R�Ҫb�:������aQ=��v     �
t.�8@8V !=�S� cT�ᨘ��Q�
�G�U_B��QcT���      ŋ�*���êy�GN/�B�=��Rq��i���{+�MG��zo�t��0����Z���Sf��nѼ�#��λ���ι���	�ƹ����u���v�Ɏ�f     ٣��p��L�M�|Bo�@X\v�@���s�E7S����0*N��z���a     �����;e���5����z�T��滿}t�i������ �nf�}����i��Q+�/�R|Oźu�X�<$�ܵ���e�K?����     �����l�S{�2���t���pl��::���U?���A!��B     @O�񩜹tR,_��������'��KV�+H��Ş��KZ&�6��'[+%�tpW����e�Ii�����{�]�(�'	4UQ5N���:��7��oC���q�     ��m
�7���^�4e��i
��B�/�
m�4Q�V��y�_�ڨi�uT}�/t�j�q�     @���ʫ[�d��r��VC�GM/��;�z�o?���M������������>=��eucg���٣���1�F�������w/:���ɛ���f�]��������%�    @�U�er�]�O{�U)cT&	tjoC��t{�1:w�@�*2�U�d�h�@�*y�     y䥏�pW��X��E9+��w~���������zԲ��U^�R%z�����?�cg��t<��B�N+����}��7u퇂!���ǿ|����꿱�C���v     ���N����k�̝�P��Nƨ�c����<z���9     ��;�)[��W����L(s�����o~a�y�!���~���ʟ���ғnW���%�GAj�ܷV6ʋ���13G���|��4g|ɋ�֕W,_��p���w?4i��Qw��ƴ=Ɵ^�P���      }ؼ�'Ч���Ե2ݵicT���^M0s�.�@���ò��p�&��u��5��Z     �����&�ŗ�N[���u�w?�č��|D0$Kf�Z7���IW����ʳ����]�]��o��f��*����1�EMV���J���ΙP�v�ב�1T�◧��&     @?��tH�?,N�I�/�;5����> ��V��lQ�hD�_���)(���R��EvG���P��4��{��l��.      ZZ��V���F�O*NK�V�I��S�'�o�U�ճ^�O���#��.I�c�����$�.�۫����w�	�Ƥ�1�L-����y��z�`@ήx�z�伍Sʼ�t>���� ��    �5����mrܬ��� ��Q���[���#���k�����Ey}y�1��׿��EN��+���    @:��_����%M5�%�e71��?߿���7_z�'����'+N^0�2C��A�m�Ͳ��]�'�����̮�N��/��If�{�%�$���Z�RPauW_�(�e�(AX\��R�f@B�&�!!!���3��{�eqeW�����|>��ɄDN����s���N��䷸w/n�!�{��]w׵g|��/o������޻ޒ��.r�g�    ����r�{b�V4��U6�����eq�?�|��w���9��2x͓���k�YK���������1�,7�   ��7�xx��]J=r`�nF�xƅ�����Olޖs��������-���e����X��7���MO,�/~dB��#���#������~�}�o钛�v�C�i����RR�:    �ۂ�ձzs]�`Cv*�S�J�o���+�9?�$H��Wʣ��)xͪ�s袵51vX� O�\u�H_�d]m,]_����܌6x   ZHk,��mh��5�L�t��I���Vuo�+n=�#���}��M���_�/Nd���i�w�a�z��9�������^s����/����]�w}h�!�=������U1���,   �k��#�xnk|��!A��6c?0{{�FSgl�'"�����o4�٭qƉÂ��E��������k�7�������3
   ��l)���_��-z�	;�ܥ�ˊ��v�^�������W��gԕ�J�[tu{]CS\vϜHQҁ{���h�q��ע�.,(�c��K�o�gط��c�7�t��5ŏ�=d�Н[�\���{^
    mO/����C�m�Yۢ��1x�9˫l�NĴ������ы�*c���u��m��e���!x��+�w�-m��9e���k=   в����x��#b��-z��#��+-.\��7�'�⛧��༫�������'݊Zn���{x^��Z)J:pϼ�dc<0ky|���m��t��g��WN���5���t����9����ߥ��v0�5�w�}s�W   iklj�k������l�h�;f����\���s>3*
Zt�	o���)&O��o��0�~xC���Q-���7WY��<eF��lF����Y'�4�mh{Uc���   Z^��ϯ��|��_}���JK���b�%�}��'?���.�����-�niK�m�[�/�T%�g.�oN8fp���>t��}_Z�q��_r�a�q��,�N�Ko;�	C��ثU�\�zuC�3si    �C�!�مq��=�����6EM}S�-]_��߯e������ͱ��.��gɺ�xtnY|h��A۸�����&^Y]����&�
��Ol��Z��   @�X�jk>z>刱-~�A}J�>v�n^y��~��/�N����~Ȅ�6n�?ti�m�M��۞����HU��˪�����?x��_�>�>|@�Ž������z�U�	���ר/�V�*{Y*j��S^�o�   ڏ����=�[�]�����s�*�7wӓ�c܈��yP��u���2��=xs�?�17��cx��u�X\�.��]���=,7���ַ�gT����   К�~��8`��3�����Q\p�!�]8t���}jޚC���Ś�d���;������&�k���l�����=���q�S�Ƨ�*�ػ����w������m���M�ԥS�ǘ��)}��(},�dߚ����Y�a[U    �KeMS\z�8�Sãk�V�N��k�G7o���9.�g}��QQRlF[˦���Z�������O?=*���ֲ~{}\u���ew
��=���E�f����RW=hF  ��W��?��\\��E���-~�lcy֬�[�v�eS?����0+:����sď{���/-���-�Ե��=����޻�=F�k��u-��g����=��'����sN?����ιjʷ�}�����l�uVw�X��Y   @��pMu����q��C����m�h���Xu��+�/�cM|��Q�B�WQ�ܶ&�#o��Mٌ���8��B���:�<:eMTՙѷk�������;��vB��V�LY���    �-��X���R��	���9���wh�3{]{��Uˎ�ZG^L}�巎�uP�;&�2�K+~����6~>yF4�����U��]r�����}8�����Z'��?p�}9����W~�3?ѡVf��?o�g���M9`��ݺ����Wn�=	�   �}{fAE�*���� �{*�j��o[���wf����F�o=D�ق�k��?���_T�;3wEU\���8��!aD[NenF9%7�[�wf֒ʸ����Z߂^�Hhul*3�   @ۺ���1nD�8�]Z휽J�
�>p��,6픳.���=퓷F2iRsA�.w_vĄ�_��[[�܍M�񳛟�Me5����=�q{u���/��U��/,(��a���U���z��t����w��+)�����Tڭ��+���6~zӳ�   �����GUMS|��C��Uߒ�6no�����[����3+��ා%���m{Uc\x��X��6xw��R��M����B3��e[��{]�ь�[��-�=�6���RdFw�����gwu    H�o�����=F�k��޷��C��2�O���pS���v��h�~|����?f�e�ٹg[�������e���hw�{f֒��܃����m�s�SRt�������i��«��׿��[N9�1ڑ�\O�L��3�������7��o,�   ����̲��8��!ѫ�k�c�_U��{]> �ɶd��ϫ�[�����ۣIZ��6~}׺ذ�����W+s3�&N?vH�iFw�W��įsϣ����\\��ڌ��aFw��k^{��R�   HG���ᙸ��#c`��z��n��O~����w���+�U~�?�8e^�3�]s��F�y�����ui�[#�?kE�:}q�'����)ϼ����O6�Mο��>���۫7W�:�ڻ�0o��o];�I��?�������}G���=���'�����B�]�9   ��g�����+�G��#K�w��9b�-q��[�_�cd��nX_���8pt������{h�����M��hHw�,t��������W3�^d3z߬mqӴ��hFw����s��+��G��w.޽lF�z~[�2}s�6�    ����i�}0ztk�츴[a���Ě�/�1���K�V}��o��|$������C��d��i�?�����_�������C�����ٟaĀ��s�W3�K����u���=��O���4���`��SG��y��;�{ri�{��������v�   �Md�G~��8b|�����ޥ���SK���5�l�%�j����1.�cm�[����^����6�fk}\���l+>;^yuc\t�k3��#�����|cm\�Ȧ��x�]Eοm�k3��A�8�.,]���G7��I�O   �e��ܛ���}�(,h��{qa:~���m�����^�������M:픊H�/������~:vdߏ�4�W�o����~|������M�~����9Ν<#~�����1����2�OI���<<���V�xmٽ��T�{޷?�R[�y~r��c�.>s�Q�6���H��O.�   @Ǘm$}r^y���2>��8j�>ѣ������T�?�%f,��iY�r�9oeU|d�>q́}�o�v��i�X��>�xnkL�_n�p+�ft����h�9����`�mX��.?��s3jD[^6��������7�޿O�*1�oe���Z�^�   h?f,Z�:3~p��(h�U�E�]c�]��?(�����[��zK�%s��^wˤS�Z���o��>jpi���:��?��`A�6�C��zsE|��iQY��Q������)~|������20R���>=s�ɹ/O�ȴ�K7�-ް��ʆ���=�S�Z��U��u�?�������c��>3��%q��s   �\*k�⶧�Ľ�o�����������J"����PW�3_��'�ŜUb�VV�������x`��8t����b��R3�W�cֲ��.Z�ͪh�u��7ŝ�m��gm�����#���q#<��������,��<ں�k�b�[���f�W~F��݌���܌f�M�����(   �>=���(*,�3N: R�{����}r_^yL}������[*��\^{c�u'�8iR����;O�߯w�{�7�σG�ӿ�kA�dcYu|��i�����90��ݨ�o̯�?�s��^;���SR�;�������#{�vsYu��+r���U���64>��[ɲ+�v����wү���)�ۣ���K���YR<�_��Q����M1h�kw�\��5;   �Ϋ��9zi{�ػ(�ک$�U����Fׂ�#��d�j�ax�ژ��*��9�g��,�}b^y��ۣk�siL��蘡�bH���ڵ��hb�ݚ�hM�[Q/���_�B���^�[�?���{e3:�4F�ftp��(L�3��]��f��U�9��3�m-�`��9e�����{���k}I�64{��\3�}/�����h6����    �w���<����	m8�^Ե˸���玣s?=��z�u{�����k˫�U��=__W0��8��OX�f��I����yt��.{�ҳ{�޽K�wЫd�~����Tm�^g^�d��Z�Y�Q�;QYS߻nZ��_�F�e�zv��s?͎CrǗ_��Sg��u�͵��Uu���CqQ��®��
���U'�N_����m$   �_l*����fGY��Y�6�OQ�v�%�Qڭcp���E�5�QV��+��� ;�m���M�ّ�.�ػ0z�׌��f�}�]�7eٳ�*w�U5�g��yi�R�O�\�?2ٌf���1g�17�5u���^�[��h겿��_.���>��{t/��E�;��g4{��^ݘ��   �4����O��/�URT�kD�~�/�cB�8��_�̜9QQS�\S��T���P���Xڭ����k�nE݋��~��ެ�\g^3-�ok�q{�������OǏO����MvEG���E�u�{�=2?��;    �LCSĚ�����R������z3J��]�y��e��ٝ!    ���"j���:(����zv/�;�U��c��/��];-6��DGС�L]}c�}�3�c������Ô���b�*          :��箊�۫���}J���1k��8��������U����v���5;�l����wtI��TU�򳛟���          Ӽ�[����_|��9�gк".��|4d�t�!������X��<~x�?D������T�nz&��/          :�l!��^�X���1q쐠�565���7?�0:��g�-�_������c�������5q��3;�-          xseUu�?L�:b�������.]���=���ٟfĬW7DG���̆mU��?��o{�.��UW�W=07�<�j4w�;          �6di�Q|ن���'�>�������q��g�����:E����o��o!��[g�t@���=x�o(��n���n          :�g��/���8��!{޻����W⏏�M�`u�	�_7c�8�w��7��/��0<xws�[�/������          �m��q��O��w��|l��ѽ(xw��My!����E��3�Z��o|&7,����Š�%�ۗmk���Y�          �O٢�;f,����������sD����7����-������:e����_Ys�m��9.N<tLt	��������yqg�ɦ�=P          x���?���8|��8��cx���{l���9�~[UtF�:p�T���e�Ή��[���ǰ�����g������          �D��}Ƣu��C��?`��ѽ(x�Ek�ťwώ9�7Gg���׭�T?���1aT���G���w�]Sss<�����cU��          �V}CS���¸{��ġ�㓇����X7=� zqE45G�'p���g\�d>p����~�0t�6�?�Ҫ������          v��꺸��1��%������k�v�|Y�eq��⑗V�S��7	oӬ%�ǘa}�S���#��]�#��m��^X�L_�U          ��m��q��s��̏��%N>lL�[�����Y�6t�����-,^�-οuf\u����~;űw���{DG�pͶ�kƒxtΪ|�          �%�Wo{jq�����o��q��]�	ãkZN]QS��]S�y5^]�=���o�������-�=pŇ����*)��h���|��Ћ+b���          �����«�Ǡ>%����kD��7ڣ��Ƙ�h}<��ʘ��ڨoh
ޚ��jjn���?����w�s��-Y�=� �6oM��j�[          ���۫���䏑z����>4&�4 R^�^^]�/�O��6���vz���{����,X�?2�����20��=x���֦�5[*c����Ҳ��ܢ����&          �=Y���/�{���8`���w�A���b�!���K��Y�>喘�bs�\�>������D�-�P�?n��8���j�=F��݆��Y �[�s���[+�յ�b���X��,��[��          t��������#ӣ[a�5 ����C{�N{EQa�?����|��tCY�ǅ����]A��%poA��"�����g�E]ch��گG�S���޻�(z�v�n�_ˮ*���®�����M�M��u��+<ʪjc{U]l����۫c���TV���         �3��m������e��*���JcH���׳[�)��K��WIq��-.,���.�=�uu]�k�����khʷ�Y�����WǺ���~[U��iy�VVW�+6��          `�jn���옻|sо�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          HBᆩgw	    h'.���v����HPCCC����ۃN/7�����"=��8㌱A�w�E}?��/"=r3:.��rϣ�rϣgGb���g�y�    h16�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��۵c   �A����Q-�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,,�ъ\�    IEND�B`�PK
     $s�[����C   C   /   images/ba153158-cccd-4fb1-9320-38bebad1b7f9.png�PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK
     $s�[Y�u�= �= /   images/fd2cb464-8539-444d-bb0b-3750bec3ea07.png�PNG

   IHDR  H  p   ��   gAMA  ���a   	pHYs  �  ��+  ��IDATx��i�|�q�u���_��M�HK#[�bˢI�A"C���v�	$@;$�����K>$@Fx�h�)��XD�RdE�mj!-J$EJ\ɷ��{g�r�������,��;s�S���̜ӧ���_UW�Y!�9ә�t�3��Lg:ә�t�3�2g:ә�t�3��Lg:ә�t&Og�Lg:ә�t�3��Lg:ә��
ҙ�t�3��Lg:ә�t�3��3��Lg:ә�t�3��Lg":+H�,L�HK��,�9�ș�t�3��L��3�[t�K��
R?����E�0��� H���}�>�:�	7ӟ��"4������(Z��|?%��̔}z"�Х��sR�=��K���C;�6���쁔�KC�TF���������s�7ç���k7�~^�q1t����]�cN�)��� �QZ0�g=_�o�7��|���.a�3<c]y����b�����伵1g�ڕ\�0�7��Vn�i1 ��޸+.�1��Z�^6�V)҄|��-e�k�\�z>��+�����U�U����|gϝi;�c���{�g�L��a\�(2�!��O 5G��%恌a��+ �,�+#�4n��U�]�N�&�'ګ�G)��M9d�K�<�d�_N������Z�"n������$�.)H�+�"��W־��ھ�jc�4|xm����4�������'t���:7��sI�(r�NeX�B@�z�I�	@g;��mXL�ic$�iG�T)@)�k�	�ey��0��s�Z\)�U�FB9XF�Ss������ʳ[^!����`]��i�r?8m;/H�0H�l�6$L������������{=�z����so�|�rJ`w��>7-m7\�w�����t��W�w��޼em��<��R�6[h_��|�>;�@ �(ӊo9���R!�)�g� &�ymj���{�Q-�a������':�ƽ��\�����){�9}��v��V[��7?�޼��z�e����Wָ��"�v��a���`Oh��6�k
0�(�r]!���(�1=n<k>2B�	Y��W��ךs�8n=u��]u�j ���f�e������>Ȳk�Y)�p��6$m]��禉��ɞ�o\o���GW�l���.�7�'�:?�ͦ��ٰ�%Tx�r0Ɇ��C/�qr��*� �8���	�E�	e>��}���概��$�r�]�1
���7%�Sl��U�=N�(r=KL�ϡ�QJ�0���?�+��&�#F�:�g�,���=ӄ5iX��A6|���/90 �W���y墇/i�� �Za�+
��f3,N�ң�y�s���O>��ʏ?^��3O��^�^?|���ޣ+s���5�����N��7�_;�x��^�l�	9����u�E��݅��b�i`kI�t�lvT�/������~��g���@0
�d.@���\UhE�B׏C�Ne,���s����T2���r�q�ʜH�P��o?��\����
R��}�'�/h�֮�2�U{���н�ط߻��;/�Ͽ�2�}�Ë�y�����l�r ���c?0�|���=�˱訥����r�C᜴�]`�",Ǡ�N���X����m���v��X�§^��������|�'��[��b��AAv���ag�ϥ�/�4ӆÜ�-v�Y���"�YU ���	`�]���rl`j��8V�~�D�����uu�vUg���'�5���S�.�����{�j}�2�{�y��μ���+_���O�t���+x�J�p���G�!bŌ�[
K^�����A��z�����z�/ߕ	(ɣ�$��(ykPD �Q#􌛹��}�y�G^}�5y}��xb_|mc�?���Z��2�����?ɼ�`��gގ�)����3�( �҆g��u��8���%[6�}2�Pc.�����	����=�k�Zu�>�iظq��*������/;�z�
���Ë�������{�g.���;^��}�Y�"� ,d���y�|+�;�@�4��kY�ć�F/
��$":ÿ	b�u?Q��a�����4�v}~mͽ����_x��?�;���g�񤻸|�~�9A7���?�&�#��z=�gY���kG7(>�zl��$V*@^7�0/q���	�p*� }g�u����k�R��Tu�߉{�=���*j=z��V��	 �G��kKaf��ve��_����e�ld.Nn�Dn*�3�E�44���R^�x~ȡ�=�qƭ7�c��eȺ{�oV�|d�������{��{�_y���x���o]�g�|a>3�G�7(L�7�����G@�� �E����͏����o|�/���o<�}����{oyeu��G�����j����"���*���k�x
#�2$p�ec�b(���J:^�zU W�����D���I<��)a��dab Z�k��e3��닶��&{�c�TԞn�$(|�e��r�RK�`&g� I ��֐C0%;�>v+ǃN�m��4 q�}	��ӧ뷼���{����������r� ��\���~CrzX�	%���&Xy��Ս�sl�?$�5@l({: ʺ�1h���҄�z��$������X7HuC������۬�ڑ:���E�~sO�]ëx��yۇ����Z����e׭ر	����'hѓ:��C}���m,c����]g���J�W�.���i�3'�7jѯ��S�_������7Ü� z`u���Gr��i���b7����k����_ys�ڛ �݃�͚��/�3A�^7���t�`|q����,wuF<4'�.�q�QR��'������� ���@��tJ<$#��=d輞��M=>���\߻�X߇~���W�um���O𝟰��߸��ozǽ0x���J��:�r�O�Vr�!@#�DB�1ȩZ'��y�7��Zh���2�M��#�$��у��:)�݀��<��>^a������WWW���_y�E\��\o��^tA�r;�M�0�7�y����av:�O#W(�V��b#ƛ�_���k�C�����A��ҽ�N��w�]� �A( �$8�3]���(4zg�D��~�a�}���Š:?�v���<�hw��_�<�ҫ.��� \� ���eV#����w���6�1��� �V�hER�%!g	������4Ic�h�Q��*�3:�GQ�U�����hl�y3��<��P�����ݑ�>ּJgH�C�<�$��RL����<�Օ����R9ypo //~��/��/_�/|�=��?��ů�����/���A,|fH�؄���P�NMAr��ˍ�w�~����y����}�_�����W�����=��x��U�__�ު��7t+�0Z9�����0xJ"�����f!ӫ����jM8�K���;�im+qD�E�I|Ӟ�G�u����G3h. f��Z^��o�[�t͎�騫����cϧ�����E������W?y�E�悄�f@]�l��>q=��.*@�}�˶ �������^�;$^`9ڥ
�UYM72
�����H��E�`�t�j^�3�����o���?^�ܮ� ����yc���� O��{��k*�
F{�='���gl#ǐ����:�ij���X�bۘ�S�+q!����~�������\�W�����_�z�����qԀ�\j�cj�A9֫���!Э��j;U�XW��������i�0��f(�G��\�@g�V� *��'g"���<�PØ����^��7��>��iA	a�2����{4a�A��0<��Ut�����b�Iq�jsTNG����R�c-{{%��~�Ɓ`�1�����8��/�M��Ǜ��{|��x�9��`���H�5��G��5b&������kE�oԹy0L\�#�:�X�!�STow���\A�
��K���l�lv^9���ol83 �Kg��bm�/���~�{cp�ȝ������R�Hۤ��\��e_+���'\O1_����/ƥ������.lP0����"�<ߌc�+A��Z>/�x�+����跰�+�Z,KR�T�k�����@��ύ���������~���j���kx���W}�������?��^���;/�_z��co���{+p�3�4�D�� 2^m�;޸6�������g^������?��O���|ӗ}�����7=\mp3��� X���7+�����S;���O2`�Tmב�]� -��3��,���V���i,p�iL{���y�-�fEa�(B�������d�V�"^�ť�����,�a��x2;t<$ٺ�v�{�+��zP���<����ݵ��²l{�.�>��� ��'�̥J�^�G%�,�d�cU-|	�#��i��
*�����Y�t�q�����Hnܮ�!�ӄ�j ��a������\9>�-a�g��J�-Y|v��@8�c������Y�ty��l�7�`Zs�]��O�a�4�
B$��d�u��ϧ�_��L�i�v@��%~b�{i~Є�؁ɺ�ul{҂zml��Z�3 !�����@���n�՛��ƫ���s�>ݘǛ�Ţ���������s��;��E/�d�7&�E_�Xu��e{�x��y�[�2���v�B���p�n�lssj�rƊaιM���4�0�.�M8�I�]&{646��]iX@9����65��(���i��n�r��`L}�ǆ|��2�1U�W`��ڱ���I����A�6��7Oܖ���w��כ����}�-(��$j[܄7q(��|&7 ���� ���&��s��:���Z��u��x��`�V�<�/���F(GS��b��L*J�Fj!�畩�YH�r�@�I�z�l��������Ý� ��e7��I\]|v�=��W�>��k�s}�ʿ�և���w��'����w�����U�qg36�D�� �t/~���k?��G��ӟ���_z}�߲�˟\=|��O/l�S�Ż~�w嬂d�" X�Y��t�©���V2�d�<}kaj����"}S���{��Ga5����{�Z,,�qh��6o��E����B�������ӝ�@3������xY���l�%i�:��ￔ��ҧݳ�a�����B�(/e d��3�Q,X#
��%��|L#�ud�ڃ�~�p�t.�.K���͓G��4��(J�!+��hX3�	���
��X�b���r�>4ǹ�������.8u��'p<׸�;��Y{`+ʏ _�,�į~E6E�׍/A�X�J��N��q+Zv3m&��x����xiো����U�E�ɇg���E�.!+
�XU�K�����ȭ�l�=y����.L̘��F���V݁�pջ3KO���ހ�w���tI�{;�V(ִ+�7�x���Pk�N�61mK:4�טè�HZQ���d���W �7��K��3�ѝf[
y����@k���Ms,����W}���
RI#ݿ���ekD�`$���ϋJ~5�ٱ�+Zj�m
�E�$V��[�������"ä�4�!f/fur�M�!��*N��z�v�>�������݃�����?�~�?���_��{O��_}������m�����������?�'������_������y��<w�`�t.�>��Z�B�� � <.���U���0���4W|^�w�����lŃ-��+�w���RWTq�VHmI��m��	��oA9���  ��"��ltX"�x$w��+N�,D$�p�u���V�&���4����٩�x�M�wy�ŝ��˦��d0(��]##B�aE�6�9:K�Ω�>��h/���&=�����RݒȎ\��WQ����M.#oqmH�)ʤT�mI��M�덪`T{S�5�Z���
�1�&�+�ޠoh�û�9�w5�0�����%*.���D�Ƣ��#I	m�Z�2Pu���hɻT���p=ٔБ���+:+2/z��(�D�o��z[�ye�#C��l��e�h�R��@��B�ɋ�����蓚F=�w��'_A��`�%��GKqQB�Z/��5wE��w���4v��꓏ᭅ��o�J�_���ksh��%���0�ܹ/y�FS����!i���.ɮ����p�ܴ���|V�w�4��\<�������߸������v_�o���w�����~�����v�^�ܣ����}�;�֧ͷ���w��/��O�
�n6��;8lV�!��F��ު����tS��װy�x��Ԙ��T� +K�td̯Ɲ# 1w���� �l�AHq=�sau�a% i!�A�E�5I@k��)�RI��u0k����#Ę H۵�t����۲� �,) �rKу���~"(�]%@&\�ʾ%�l��}��f	������ c�u�lǚϭu�1�7� ��-�*֋����*S!��WnTT9k�P�l�Q�,��UQ)���J �ѡ-��B�����,�s`��>�u�������l*�I�ԏ�U�7��i��s0q��]K^W=��Da�A9�^)2���#g|��lIa<�!� z�B�q5�শ�j���4q��r�� �adѥ�\��.Mإ�ݜ�&��p�-���B9a�q���,>5��iq'�:*�	�p��\m.��\K_Z�"s�[I6%{H�e")e0��[�g5��y���k�1�}'�<�0����ƽ��?�d��>�;�oﯟ|�Ϟ��Vn{��<����}��{���_{�^z�ަ����3��2}�"�c�)ti�s������x�M`� �Rf(�ܲm
�%���~k|���vӔt1ϣ�d�������>�W|�[�q�c�+[c6�%�p��v܊�7PgqS���X������R�m���,:W��?�pm����T#Ƞ ��-ѱla���0r��A'cl<[�?2���W[�]���8�i|��4���!(bp��]օ�!jQ:y��'��f¬eժ�G����}�#�W��b{AT%��Bg����MUq.��K�L��!PTCR|H��4�����
:L-�B��)�6g�V�#�*B�N�Q�NKJ�9?�xp�(���J��t��"���qzU�=�Xw��3���'��a ���#,�?r/�)����B�u��p�g�3ʸ��<�Lg>����`�T��M�^��K�}{!Я����#.��������\ͭN׾	��ȵ"���K{2ĳ�dv犍��jǸά�2� �X��{j�B�����?��|��5�CG� ]o6����}�����p��_|x���/�+(���m-�sE�B�������:�LNl�M/�t���l]QF��d��;��� M����C�eN������3y���,�R�����1��E��ӱ�XT@
u��àˋZ�Xp���C�uNj����H%83�b�f{�VT͹,z�p��P��hReph-Z�d6WG�l�YL(�I�Z��T�xx.7�3�-����q����T���:h��q~���Xw]<EeӐ Jr�$?��j�KP|��AXȭhXDۢ$	
$^�@� ���җ@e�����!�e-�Hwj�%`�:���<_��.�oFg��כ�]4v�1�L�v.V,��<O����o�5��K,L��-�E�y��x�л�����	)K0Q��7m{(�:3�4��'�c�[A�L���ତ�������f=��a�Ձ<F��ӡH�7|��C��c�Qv���j@�>���;����9sKtt
��e�������Ǿ�]?�z�-��淿qpa7���̪�0�Țk�����mx�yZP��p�dW�s鬝�>�l�lgR�����P��]�$,m��Q��~�x8�O�;�0hS�i�o��k�b���o[��?`��|Q��S���8�?�T1���t>�6�YfW[��f����uW@mw��t��:_���X&�w��}�0S�+o�v}�@>�O��mkװh�P>Q&kj���!��1��e`(�t�K�h!O�!OT�;yʐu�� t�PIo�Vǝ�#�e��rYrG�3��9]�a�Ԑ����ظNCDm�Я���	{��j�)�o��t�\�B�������|�>;�����:���n�o(9�N�9��[Q���� *�lȰ4�E��,���,ҏ��(׊q�K���3s�5��-x���Y��R��rl�Q���}/`71k�񈀥R��d�+O|�Fk�� ��.�o�V�'���Cw|��NAz��<�#��K�=��_����+3(G!��������Ɏ�����u�K�T)̙� /e�e )=#%k ��M�n��4��}��{��>l|ߞ�Z�. I�	`Կ_�"�9�	A���1�p7㶧P���\���~�qݣy� 	]4qW�ܭ�x?������7a�9��N�s�@��|�F��Ҙ�M��kb�s<�)��A�h�7�zB���|���� �?�wM��t��;e�-�+^z;ٺy7&[�-h�"��‼߹����y������zz�wY܄w�����;I~gR����[�!��t+�~���*�����٥̄hr#����μy~�̳���ݱQ���0��pl,�u�J=��j�h}������95ٕW������/�� )�Rc��0�5�-.ٲ>)���T�P���Nεv�j$a,���g�n��r���:�<�n��>i�?@�#>�hw�;O?�C �w��hp���^�tt
�k����#��\����j�>�{O��9bK����B`�g���J~��{�Ĺ�6��|ߥT��1E	<`�Ӿ�����喆�h�3P��-�
AUwض��^���%[:�i:L�$���j3Ȇ;Y����~Z0�ΊMgts�Q���>�m�8/}�"eWW�u��A��Q�s�A���Z�QVA,uEk�%0{ʱ�Q���~*�5�k�lÑ�#����<Ka����Ax�"�ֲ���V����5�0	�ģV�X.c�9�-a4���9�+qx�	E&�`@^c�|��ID��ј��N�$��t۪�&ymN��Hǌ����c ��F��u~��'�YWh��4�h��H���߭�������.�]��A�]4S`����dƘc�@�c���mQ񲣧r)�^��o�O\I��v�94���y�R:,�4Oָi���bv��Imu5FF�F���uݭ��Avv����;�"����(���W7��?}��?�=n�Lo/�}������M߉��K:?x��|�#�vA2Ic@eFc2�����c�����$�*�S~ۆd����W�e˕�VN�QU�T,�i`rd|kH���I}(˪���X���U��ؙf��f�ǣ�T�T:>z,_������F� �P���s������BYv)���,y�2)�Qe��)��20R�R*}f�ɧM�^d�Գzn쾼G+:����1��u���L�n�p)�)�R��5�M�.3X*3r���t��^os�)Y˞��3)�����p����83Zɮ+�F��a��Qّ��aMٗ(&Jil+�W�ށ���r��F�����bV�7F��v�L̾i�w�����cЪ�j�׬8���@oP�U���쭌���S��xzi��]����ҽБb]��^��N�P0،�W� .����30����;GeY�jw)\o��ۢ�1�_�V���D&��BT/T@Ƃ��:����2o��w����練:[`@4
۝n�bQ�,pl4��	򎣨bu���*�q�R�S�Z��o�8m�dlC���+�"�!�,�t�!����A�)�46ogy-�(�hqIa��M6��p3�S�'ʽ��1�R��L7�W���`ͪ��ɜ��!�+��2k,]O����=(�=*�������-G� ��N۵�p��r/�������I�(͓ �^�-T&-��$�>�ֶ�K��~�2QVk���}���g�u��p���e�)�zX��"� �!�,�WilT5���C1�hy�Lf���N._�6D��CM��N������n�A�:%��H���`C{RS&��kJ�|F���I!�5�ף|>�4*&��Z�_<���s-�\�F�>0�8�2�$��Ɔ-&�X��BIҟ�n�Wֲ0oo���g��=��[J����;�P����\h����3�p�i�ؚ�{�&��R������ �u�tC�$��4}�D����_�\>�4��D͊, ���C8G�-1�!p���9>��Mb�b�N)����;�Ft������W���n��NAr�w�rʽ�VCgmzZ�($ G�
}[[�幋r
���ƶ�K7����!��W9s&��^����I
���\UL0�8A��Kቦo|u���T-�-L?J(��l}[�+��*��V��f��]�C�n%M�f0�c#�^5f}���� 1�%l�B�7TD�j�E���S���q$Ĭnb~Vs#�E^�S�C4@,�g40��?�q�+(�ҚW���t��1�����u5h�iG�at��|w�r���貞�G���vηI�g\$�o�=͌˱�\y�OM��n<6��M+]g�iKi��$3>�F��(%�84�xjm�z�t|
��3�r�Hл�S>BC8�.�e��!�F�_�VE���띏��1s�kˏvqk�-�9�䘇	5���{� tX40K���M�[��H?���p��s�UB���G�s��)<��oU�Y/CG3AY�eZ�;0��[�@s�؄۶7A� � �ʢ(�Eb��[Y[��]�i}l)ژOc�~����������t`vE;�1�.ي�}չ���� ���vx�9�b�q٭h;�"4%[�F�2%g$�r[ �B���1x�o`��K�^tnV�����\[W�� r�Oq�;19Ϡ��W�5�a���#��H/{���̢�Zg�d	n�:Q�c,���!����BB���t!^�!��ݝ�&������5�\z�y�Q-]�7�`t�P2o-[���2b�9K77a��B�i���_�����Lm����{.�ı�f��Xü����GIy����̛5:d�!ky�6{����K����\͍L���?o�����M�P7�v��c�X�X��������k���v���G�[�%�HM����bޕ����Bbv�v��$WI�`���{G� s�������:��`�|�� \����=�T�F�6kE�v�r&�.��h��lY۟R�1q�(��`�B<��cIѭ��_X�te�0^e��a���׿mwfk#f�şJ�`�dJQ���vav������Z��H�D��Niup��}�e�Ǩ��r��?��i���T�,���d��X��s���R��X�R��� 놩0�@�|)rN�����t ������UF�B����&����:��	���O�~6���SG���iG�z�@�=l��*��y�B]ې�V
o�@g��9P�(���^�:W��N��i5��:^4dr3 �Qy=�)��a���H�T=�(����
�^>/����gEFN�v����9���H�A%w.�,�ۂYv*�mE�mZCޮ�*�N�@�؛����3�u����D����GnZ_t��^�=�t�
R�H�t�s�(���LJ庴�PE��Nyk/3�D�bq�-�p�tN$���ǎYD��u��)�G�R�Q�RT��@PPꇖ�F���C./c��JFL�@�F��<)G�@F� �yr�Jg��c�P�]B���E�Q����R�M��ac�i0��D���sX.�h�G�/?mP	TU^�ḿ_K�sԹ�����HvҲ�,�^��/+\T>F�1���w�����+af�[M<~����=;�QXRX1�x�QVר�R�(<3��_��q]J�͘&vtH�s
��k6^�m!�x�{��y���ql��,�=`�����~2f�/��.R�a�n��@��7�a�����軣S��	˚�D��̛R^��+S�i�jK}*+���9qn��¥ai3`�4��>Ƒ_��e����OњW-�����TY�ŚW;�����ނ4��rQ���D%����f`��Y���D)v��{��Ƃy��U���tvi��t`2l�J�T�TeEB�o�Cі��a�6rk�H�b5���Q�,�z$>���Mw����刣�I�������	!}a���p��銍��~HS�Z�j�15���U#�R��������-Ol�&6_E�-v�s�"�g˜2����G�@oQ��%*�r����ر*��5�;֙4�C��R���G��+ҫ<n�A�NA��wr�b1�p�����B����I@{[V�S'���T���y�.IC�4��g�b)����E*,�"K-���\U�y����2�R�	ϸC�5R;�)�0Z���_I؄a�+snB|�(�K�������%�2�)����@r)Z���]�v�AKP��]�s�=�(!+ہ"z�2����wQ��(�LTd��G��fc��?%e�4u[J=u)��9O%�_
w[�lܴJo3�K��b�s���HUڰ/�K�m�h�����Y��@���v(��и��G���1�ae�(d���k4�����I�Jc6ٴ]�}t=��\,�m>��ˣ�ٿP�e�$�Iǧ ���	D�P��hrd�0ALV�qV%�S�hܯ2%��tf,d�F�:$>J�H _,7J*«ѬW�2·\C<5�).�1�����4 9^���턗)^�X �j�lOe����3R
NLN�%��b��s�	(����3��������-�(S!���>oU�P󉍢e���܃P�WC~Z�lΣc?s��@�����T��ƀjA��3n]ʁ��R�/�#�P�RЏ��9��A%WH�dWv6؝w�66V��!�)���R�h��,��@A�OII��-H9hx����c��\9u�g�:F����0�H�ԛ/A֥Q1�t��ې̩CS촎��z����yɍOt�f+2
�<*�Sj<>�k5Y��qj��$zW[4�y����*H���ua�:�2���R��>�d��/�$N�����Dy	ێ�2�h]��>��x$�������K�x����|��T�]�d���;�s�� 1��WX&� ����L$��i�f`I	B�� ��VQ�.<#��r�>��2uI�I�(���a:,���.*Ɉ��hu3[�7l&o��g��Vh|�+�'��0��<��'�û��J�gc�b#Jm�϶���,I�)�x,`���uy�G�+W5����~艍�}�A� �mJ�!�XF�򳄫bTR��@g�R�b������߷�����;�;��A^�Ƒ�gbNv.����-�Ԧ��+����k)&���+�v�kk���Zѣ9�|�+���h��$ ����4�-�v�)	��M�K�K�c�G3�<�I�l������D����<47��ظvC#wa	O�2;^�����7HG� e�� �N��9�nK>P�\�k�BA|���y��mi4�$�J)�[k��
��\Ej�Z9wa�+�I��&�JũY[�� � �T��M�連8�ZU��ӎ��	��u�R9O�2�Ȭ�aw�\�t�"�9.�.�әB������1B졭��*�iI)"���&�PY�f����J.}@ꑰ* �L���[ӒLNM1���l����d����>�͡b$8����ʺ�]�r"�G	�<�JF�2/F:j�s�ϥ2�3g@檒,	�Ә��%>cr�~�j))��5ezS_3�3���US=[#��E��rz��s�J 1�WS5K��Y�t��n4�I>�cy,��sǧ�ݕ�藹V[�S��܃5����>k�H?FM�̀���p��.\�s ��#8y���C���/P==*�bЁƨ0eQQ\+�4�=�>��m*�9�L%��[��%��(�.5�����t�G����aJl|���1<1M����Ô/��f���;S����m��6o�p��x9kn��RA��$z�c���"i��q:K�����1ߘs���2�?7K��-�B�nQ���JU[M}��Z赶O?e,�u�����i�}1Ov�ib[��'��s���9�~Ǒ��8���~��b7$�*��t�fd^q���ze��U`{���L��GE�P`��tM�jǘZ�C�5���&�����hއe@��ژ3탠��&�'���R�O�n��G� a���aF1"�-b)I�1 j�i�rⱁ�Qp����3��B9.~A\P��|0�.4��^��mIۑ"ߗ�C1񅨑a�3s����׽�̨Ăv�Uυe�΄��$�00���LϨ��y�`*X�����}�Ƌۍ��aO-7�a�=TVal�O�y�$K�f[>6�J�/.�Iɴs׬<%=���KKw)w��b�p��0��!�����{�(��	6b��f��2�84-�i5i��]���h��o�Z����BT���	����*����u���$G(�$�Hjl�6���d X��*��2���m���9/����32x̭�T�2j���D�)
yn �qZ
P�*�䐌5�I�i8��EFڕA�O������������n��FMQ�����%����ÐT|x��M�*�dw�v�a���߸�oD�l�쎹��X�rr���ŻLS3.ډI�P�MؐA!r�fy�q���qq�Q*H<�a���5-ָ��N߁2�S�0�^w|������a��Ҿ��;{�K
A\�2m�p������֤."�V���) =���.8��p�K���	��r�x ��dkJ=��[?�eF����<�;�e9��E,W���3����3�NZ�Jp�E�+]ꖸ���Xh܌;�d�5	�L������I�O	;�%���w.�b��ϝiJ�k=V��d  ��;
9{)/h��x#˳�+Ub�Q��#7z�2ٮ���A4e)x�t�&�/���,+�i�E��}�=��Āgڍ�l[OY&�0X�b=t|�����3�&���_�E�t�m1C.�ĺ'�z>c�� ҁ1x�Ly�
��RA}�E@Ό�����3g�3�pK���>V�Q�f@�^�(6���*��z5�4͵�j�k�ޖ�VHj��#n2��[w��U�J��L1�2-�%%�]��/�-�i��R�9���P3�<�/rbf���\w�˞:�&ܚ?�D�;Fb刿�؅S\��K��Z|�9q�yk��ʰ�v��ug��L�X;��
��&>q�݃���|��Qf�&[l��[��T�-�>f��)�����h����v�l�3���I����0���>�t����?���g}g�٩	���h�7�Z�잩��o�p���AH���KB=�3�w������
K�H=+�;��E�i�Ԉ��
�mܨ�/:V�W)ٯ]�P��mb�ڡ��(W���"�=ˆ�e����3Hr�j���d� 0H���F\�Pnά_���,=L��Y�o�4�_�����g�^�v�P��@L<TRu��Q9�Z��"�7���i3=WmN0"u�T��6���$�t~_��%>��5�k�mV��±	.h��W҈'�[���6c�q�:D��D�.jc��<�;7��#Iց�r(��7��4z2x�r��n�']s��И1bv��P��e����Hr`��p���/�����ug�4�oC �h����JH}b��qlH�j���cO�f	(�y���}�X�/qi���1�]�w��#&���#�%
�ڑH^`�QM7���8ֳ��m��]��*�� ��|.7�l�{0�cW�I��ʐ�)�b�公9��*G���Q�qe��=�����G� 9ʴ�]�K�q��ʴ�3%[Zќ�AI:
��e�b��K��*E���]�3G�c�N�]6ܞQ��J/]���T��:G���D#�U�*������9y�F��P\ G.ô�Y^cE!v����Ё�eS��2����߾Fa?�r �It%��/�8����{�z'����N|N���U��x����_�̉�9ۭ�5Ғ�Ȕ��@]E%�2*c�15Ն�܃��ͻZ�
_B�h�(�,�C������*HѺҺ7F2�]�xδ�_i�s�Lv�R#?n��ʄ��g�w�,���F̀�c����x�j���v{���i��}aݲ]�0�o%/���c��g����F�{]j �S[
%-��j�-~	Ǜ=cc�2-�P�L��-�)��)����KrLvM{��%��u�K�z���L��/������������&o�`C�E9�#�'ǫ �C�r��ֶ��a0�F&e�-n�=�֏:i��S�#��;Z4����90��/��4K������-T�w�����L^=��p#��n;Ky��+[�Zs[�Y_5o�����"�̢kE"�[�c2w%7P�HKvI��z���HfUQ��"l�2"��?���b,ٺ�ET��T亣$����a�O��� �q>�
�ǁ��bA���Oi����f��=��t�-�r���=0%��p���w�R��/�
�ӎ&)���#��A�Ö� d��<�����g�g����,#Xj����-��;y$`������T%���L����ŧu?�q!� ��kFɴ��@N�3���p
jw��eS�u����U��R�FTΞk/�uO2����\,.׿�	b3^����v�$�* @+��_E�Fe0�c_�!��)-P�[g�刬0��x?O�1������j_�2���̥~3/Y�ZQ���h���9NR6����g��t�������(��;N0i;}6Ϩa)�b��"��K�2'�a�p�����uI&3��I�X*���1���|�T�奉y��&���%�}:Z��Чd�+�����Z 5���"���eC����~��w�.�ғ[�+|а"6�%h�	g��=d�9Q*�[i(�ևp��@�c)
2:W���N���N��" �ŌU�ߝ��#>�)5O�#��=?��>���jR=�H�N1����/	���4�S['�zN�X7,[Y�2����r������V�L�]~n�ZD%;�AGG��ғO�?�oqs
�2ް&�#����x�Xåѹ+1����˰���L"O�YX*;���ǔȃ��5�EG� �h,:I��'X2��/$}�f�y+�����.�@c��SlWS�X��U�,�C�bay�R�P/��`泾$}y�����#F�4"��R���ڶv�]��oN^H&4��E����mĸ�6��f�?�Hc�5�-c�}��m�MB����.S-\�yu�dוx$���v+')��u*]�vʫ!#��ӣ��m�Z�?�l蚠A5�뽻{]���6X��g�`����Q���Z$�$�`��2��M
���p\w{2�h$,�/aV�~� �x\j�3ϯ��l<����t���,��^[�p&ײRA}��t{I��ɍԞ�wM�-���h"�mC�\�Q�Χ8Oz��ʤ�*/��W��N,~sv�Fl��i)�~�ݞK�)�9���'M��Z���������_��8��l����@*�%^�Sv����qN2�?�3|F(b�Y2��-HU�m!B���C����ڧ\�X���Ȩ�ؐ0Rm#`t�\f�AE��Xn�
���$cT6��k�w����l"eU~^��]h�~�-_��亿p8��0Ad����lT����[RtO������������|�xT�m���p�-)*�b?b5���_2���H���<v�@;�i������YDc�Ai�th��b�2BA���$��3JZ�%$�/�v,��v�P��9�h<9� ���)>!x��PEG� � 0K�^��k�@�4&��Gh��)�s�����:L��u�U�儉��(y�}���W\��I��۲��י��L�G!�	�(nT���b�^f���.��}_7��?�ב�?F?
�OJ���!�bl.v�Z�e_`*)�ܴ���T�@��wK��)�p���H�<:p��e=1��@s����Ӟ�d���;����>NH��Љk%8��Mq��^:��w�����:�
�K��a4���CL�r(�i|� �0nhN�H��0�9��Pn���xP�Lq�ZF�K�R@�'+άB���ʁ`����%��2��� ��N���ǑC/���(R9di�a��q�r�@&9c�	��u1<���h� l���T�Ee�蠞.?���8�N�ҵMSRo�˥�����Aв�k�k]v����;C���3l�^Q�󅓗�3H
�d�d[[��e'L��U+Lb�.l����AVw���`TϚ������v�6d���C�e����8Sl��hrה���X����J*#w��CN�(�ߴ��R�oE/�B6~7Y{����XJ��<����(�l����7�ؤC�l�;&� ���IL��g�I0}[�����l��%�,���1\.��'��CSm0�6姰RgUp�$�P�K9�����QӦ����B:���d��˖���/UZ�4��Q
*;As�B빱���7}NZ�X2�H����M�L[�1Tz��f]�[ȝ��4���h��fYl\B��QN�w�Ei�i�a���Z�z��D���LL7�Bp���17( M
H�Zִ�UZw��v�K/W�˳�3mO��I �L;�y,�j�A��4�׋��Ӊ�\����2�u����!��F=pO�Y)zg]z��g㫮v�\Y����wd�B�\��Sq�� ���~�$M�Vg���<77�C�>.!5�p�+Y���+�j?�Ѝ����w��U�\��R��	���[�1�{����*�- 
�;{��R���ܴ�QK�̶�av���Y�F�u�f�.*u4�	����Y��A��U-�c����T<$�ֲ�35�6�k�t��"go���w��x7@[!.�BC[zN�vA�;��/3����9���a��Kν�1�V�lE��weU��9��.�2fG� 1c��ص+{�J��������"�Yn�:���H�mr�YP�P�d>�/����!N[��ߦ1e:i5����]��Ol�ofp�%T
iP�jO��;�ߒ��@�~��;�ޛ���[ Ʊ���-�3���(�0�V���h�WGL6rFf^>�;N�C��r��~W���\N`N���nj�w��-h_G��c�G<�e����tq�WߣU�� @��R�;(Ch�Ց��� TF*��u4Z>�P0�ܰ��v�r��La�)��vB¥�Oj����g5S��z�.V��H��Q��6��ӲxQy[� i��A��ہg�v��Y ���:X=�&TB���5�*Tڃ@e��btV�r*w���
����~'X�s��i�=ӁIt��S~��g`'�g9������9��]}�#�ϰR���f)s!�Et�j��I����R���� �F��8�o�q[��T��ۜ�R
ȡ��4�4{�Qۻg�7n��RA�ɬ]C���vY�(�K�� i�@�^�ߗu����V��4LE�2����tZ6�,Q�^#r��	�v	��Weaⵌ?�J�5i����Kb�b�ĩs�,�]W��ATZ�0D��A�b�S�++H������d�� F3���p�́���޽�㳬,�>��=�0����nʕ�m�q/��z˄J]�43'�D�g)J��bGX�C4ۍ	����Ux���8�Z
�0��xGJ�^s�+<0k�$��X�ʎ�T`�����H�v������!�ύ�n}W�c�Z
d�\��e�5�!�
,��W|�#Zi�t�m�LG� �Q��
`�6Z'[L0���4F���r3���$;��3%��.~BZa����Lh�n�)��W	 b��n*Jz��uD@h�C���XfD?�2�[I��g��B+�V�%�p����.+���w扛�r-�w�s��ș�{�D���31�i���P	BuC�}+�m7�v9�Ρ�B��9��*k5G�r�'��Z��`�L�W)�
�N� *�9!jWE���t�ڐB'� ��
�Y-��x�ځ�zd�Ϟ�9'�����$��
f��GQ$��$�I�`��kq�hFvR������џ6�BY���0Me���:�+_IG6OϴwZ��b�;?9�0�\����R)��w��7�1�h�s�\r�,)�R�_���$(>%�s=�� bH�鈵fDDFov"r�o*$��+�7�SS�p�BP4�S �!�,�n[�n��,���V�F�2�����`�j�i��Q�֘˜�����8� /�T(���D��TT�N��iO�Y�[�5���[��Ю��Yr�dH��c�(�V�J�F�-����ʠ��M���c�2#��Z�]���94���To��8���@~E'Gip�UJ��l��O��;=~�hu��䷋Q����%{���aw�I�-p�h�`�Zg�2P�k��B�F�M�u��:�w��:�wV�N/���M�3�Ul�[�Y�2&{�[��8��	)H�I�����_�rTۚʀ��
�Hj�AL�H��۠f�8�m?���Z%�?{����/��c5�иp�[�]<��v0{����&9����S\L��x��BZ���I�Q'Tm�|��npL���g�w'+c��@Kʵhߌ�,�M�\=Ҿ�c*�2��Q�Ѱ��o~��9tȱu�	�ݖ|��y����O��M����RY��W�0Fl�c�j��ˣ�X�(��5L�|u
dKW����w�h�R��x��Ak��:^ u
d}�{˭�� װ��h�K��E�3�IX�U�k�0i��YRڛ�&��3�Vϔ�*���$Y�kf�K>�;6��V5�� :RX����j5�����&i�d�I?�+�|���{F�!k��PNp��m�ww��g������P�)��A�9@�Z<��IWίmkm�Ӽ(���3�L7p=���{#�F6���l��^���8�7��<&�/?W �b*W�:0@z�N�����ԌOigo�`y�ۊ�2:�ls��uT������E��܂9R�@���e�W���i�<Ӵiy�+�XѢ4Y ��ǩ �~C^�e1��Eki�
pL�T^$�0�.m�6��
T^�)�(��*/hF!�L��r��0�l�e�@hi�1E!Y\�Bޤ��}�1������w5�{@��m��P#�!������؎<���+x&�Uۍ��Sz�j7�1Ӻ����Hw����c�ؗd,�T�Ko�&�bY���GQ#�� �S�L�㷕j.���00f�����[�wUN�%!W���"!��;���� ��F�ZGU�EB������f0��X{w0�x�.K��q.�U�d]I��R���Ch�k�ƳC�|7P�I�c� �����b�*/)+n�{�vgV�dE$=� 4�X�(�ߞ�k���4B�w ���	��j㖾� ���ɉ~�#8���v����Q�WRQ�d�����w-��c�ڙ���9v���s-Z��]�3���	J&�L`���?i<* o17���Qz԰,�W
v2�Fà�D�V��c}�g2���(���ZY���V�������e$�[�]{��f��(H�-Cڳ��&��$a�S'�9)E�-=���ΧԦI��{fw��P�qwW��i
@�qLl���5S�/�eCWe�v���WN|�-��JwՕN�h'j��2��K�f�*(�$�=-2"����d��[Ќ�z���cǞ��\9d�D���ZI#?4���v�;=ƌ��i
�|6��:�ȗʖϴ�d<�c�y�{�-g(Ij?C�75.�y��ػ���.�;��e�B΃��±��>z�w��w"d���T�y=q'�Q�u(TцR4��\
�{}��!n
멇H�^Fޘc>��jG9l!k�	nQ���_���ϞQs�ͶР��?�}��?�3�sV�N��ؕ�*T�Z�?v4P(�
�DU���[������#S��pWi~D��g���e�`���g���k��<^++hX����4S�NS���aF��� k'l����a���U�$/�ٝJK�k��1�"_�h��wOv�c�G� 1��[�|2��hL#7���J��4�A|7�ѭ���Ę�D;�5���֓��V�Ԋ�a���.+G�EN�ݦ�&^��i�c����p-M  ��UR@֔�վk鎱��M�p�4�)w`��ʛ����"1������=V^8�E�S6��$�Z��FQ:�׊���Qq�Le�A��FM�W��yOo�Wj�����ㄌ9���%��N���u�1�!+�x�d$^�NO���P�LgZJa�C선����&(�|��O�셰y�����v0�H���	��H��!�Ӑ �7d`�p}e���-�w��2ZA�G�w�c�6��V;��k��mik%�� �@|�Ah�5����S�KIŮIDJewˁj*G�L�F��cc�a�ޅZ�ޝ���zU�A�~�CR�lY������-���v�%'� Շ���@3�� 0(��v�����|��]��
E�tЊ�ŽV��B�t�?BӅ�c21;Ch&]�w���p�O��ҹ )�������t�cؖ-����B�p���ז��@e�l�"�,O��K��2L��~�;��4C�rqI=�~�B#���0��C�2^i�i"u�M?����-"Ѧ��	fv�;o�`���5b>�@l�AvѼ��en�WE�q17fZ��������/m�0�4M.����ѿ�w&��N�{t��yG��!E"4d�(�HX�,/��,Wȭ�Ȋ)x#{~,Z�a�d���s�m/��y�Y��gڕ8\k����r�>�x�����$}/� ���(+�І�|�����k�M�o-�3VԜ��-��Ә�w�r5L��
y�H-�{�3�"����A�ع�a�!��ZO3~�jZ��Ү��(HA�����T�1yHj�fog�rz۱��������r@�3x�����g��yO�B (J�H��!���E�'TߒW���F�
�����wO�r+h3�i�f�"��Լo�o_T�KZ���yMg<v��O	8���;׾?P܅�u(Ɩ����c��X�f'z&���i�<�ޗDk$&K�����;���n�NFA���HK�¡t�[�Zy�L�A%(5�C�,��ԈձF.�aX�|H��	r�?���ES�"��k�����H����=0���2�tvyA��k�ٮG���Fy�A��w�۠�T�
o<�t�|_I�)v�Ogw��ݒ&#TȠ�%R.[g:=��#H��<T�X�t�rd����ɾ��pVn�m� ���ŗQIK@������]�.S6o�D�����k.u�L��F��s��>�#���y�Ҳ��.#'N���.��JV�]��PLg��A	wT�'<5��Y]{A�P�I �A% dV���U�QO�\K�ry�*�Mj$B����ѿ�Ux:s[t2
R���Ha�̭���:ә� W�#o"��JV�}��2�oD�0'��H����"�b�.P�x�<{������h�v����~q� )� ��_�L�fj7�:slJ��Z����l�p!ص�"�U�ep������4	����L�V
ϰa2����oB�����{���͜t�M�2�̙N�t��Mk�1g��=:z)m+�V.*U���X�qX�~~����x]���,y�ۙn���Q _Ӹ.�D��K2b��x� �����ZK�f�8���3��h��~��c��[�3
��;��u;|Z�[[�y�n�=**e
�B#m��F|��}�1r�jp�
������}�[���Z��b�r��[�W��u�p/A�| i �����R�����ǉ�Jna��R�p�]��6���]'��ed��b��>}O*�x�3�Zpıt�I�6H��z�Â"/3Ð�])���Oi��D�8����xG4��>c�CZ�u�b7�@|�r=�#��ܐ�mxe�o�>W�������S����e�N7Q)V��G>��lQ5�q���s#Gx�)kL!����e6f;L^���7M���V�Ye�h/�lJd
�*�Ϯ���ֳ@SKx5�Ǐ 5W���h��ƹ����-
%fQ�~��L�G�B�<��"��r��3)����m^�-M)9�߹58]�K|Ɔ��@���T��-@�k�=v�x�	�0{ߚq
p=�ֶx�|�)��R�"���9�a�,,���P�e���rd�t�M��6ׁ�⟱(@ba]��~X_���	�QN5��m5���TL���UtU\I���J(�N=pDfp#�h� �Y�D��j9���6�$Ŕ�r�<���m�;n��g���N�0��j]C�E���LIl��t[��EJE�����i*H
e���� ���0J�6����h��C�Ho�gn/ږi����^G�f�'���H��'l
��w�Ф��.���͌���H3�6�l�\^8.���&V�S��l��i��Yt��徙���K��Hr�_¶��+�ؔ�&rWjv<��vk�]{�;r�gJ3��EP~�����g�9����4s}�6������(H��F��A�p����❙�"	0���[
�����>�]l0�E���q�UL\�2�O��񭱾�E���ƙ�x��q�.��c����t}R22)!��K&��Ѭ����������ׁ�>@((�{W(4�o-�Yϡ��0�U���`��s�t�Ji]��K�S
B��4�`�\�)є�nuH�}G��y1����#a��� �'�I���g&��/����Ƙ���>��U;E4��ְH��H٦�����z�p��C��1���S�g�<X��ϴ;���[��"ͱt�}�]�1�p�*�{jh~��1�XQV������<3�,R[�$Sg��� �Gb�,9IF�K�T��PQj�Ť>H��"�a���;�5��nbr�R����5_߸Q���Orklz�)����>�;ʨk�4�K�ȌLʪ�%-PT�4�ǭ�}���S'$�	������WH�y���j�����)eg���x(�,�~�~��([VZb�� s�A�<3=�؏���3�9���+E�(^��mfQ��@r�[Lk)p�1$�sV�n���K��#�N7����׹s��bP�0hHX(�eY@����k?<.H�P[;��BK 1���R ��9?���3���B�5R#+y��U�2�5�0��=@r��&F<4��/�T� �+)� ���|�{H/�}�E�\=&
2�D7�)��|��	Wzχa�Fv*��b���������@˲�y5J��({<%d,UG ���Hʄ|t�8��?j��p���e��K�Vݤ���Q���~Ʋ�-�4�৹ׅ�qA�!/|����!$��}y�$�M?㙹�++Z�]V��N'�(?���tZT(B{6�Cl�R�Sb�x�Ŀ�C����)���9����)��VěY4��	���t;�G��p��'�Hf��eu�MBqrV7H�5-`�=�_���ErdUnV�\�p�ŵ�3!�&���Z(z@��h �.��-i}K����bx1����0W�Cc��دJ��a_Vy��Es�ȜUz��p蝑�03�ǫ�]}M��C��)GE5���VY]��T�cR��-�"U�X���֏#�m_���Y����T!���| �o��?�o��&vP������O7��\�I�����t�$'4.w㔜���P>c�vs�t�$�:���{�0Y��'���!��:�g���)�m�}H���|� �N�R	+�l�"*,�&)N )lU��|7��n�]۟���d����[�r�&�
46>( ��#�� `��h�$B-��J.a��dJ�R���")��K��k�&�(S��d���W���>)S7G-���H�)��vx���,��d썯0�+ܮ"�$��w��^���G�-�(7���v��>��}�e��#�"L
b�\�3�Z	�nO�g8�֕M}�\O�tR���Q�hw��X��_���������m�w�1�0��箰 ���א�1o��f�w��҂9A��v��`��!V��{�k
���`�UՄ
p��Q����x>
gM�0��s���w7q�ة9�WWu��=�$^>����<�%g��s�E��=�Y'�����>x��mf�8qϵ�CS��ź�r�w��X��H[�\�G��|#��,ƀʎ<8f[��Uc
e��j3�ڃ�O�1>s��0 � ��yP��{R�ZdQ�tLԁ.g�sf>�N����h�$����|�MI�S�X|�X:R�:�U���L��r��aM�������ʷ|���)s�t�
��|�����>���ÿ������^}t���ۍ�����R.2�����s.qR�N~ۘ,�������2���d>�w�FG�a	��>�\D|N���_M���y	À��@ �^	�"Wͦ�B���p��Y��L>W�Ń�4�
�rXۃ���v��eO�x�<p� Wq[��VE-���Õ,-�,���o��s�K:;�Ԛ>a<G�!����OE��.���E��R�����EM�7� >�����`�)��� �9l�v{�M�x��k�)#yV.;��t�.��e���<c^�C��޶<HM�̚�塎'�8.��R$�@t�.� 6��f��Vʡ�8E�	�j!�Y��{�T(1a�ج�-W�Ulv@��@�\:��;|������+M>r=CE����l��Kјl���s�(��3�]*��8K�2�.���������w?���~��|���?�����?�U��́���/���?�ӿ�����ٟ��_�Է��*z��J�ʲ���m���GN�§Br<G-�(x� o�R!1�x�ka��?a�@C�=��S���C�B ��hW�H��`8k��G�@0�L��V��!I�~'��fH��A[3!x��� ��v~�nc���,����mHsݤyk3�V�b�� �v�<֔!���DN�� ��j�P��c>�[�²���c��*R�(� �!=!��M)�LeY��-)v�X!�$�7&DN����}䀔��� ���W�a��Ҷh3󘅼N�R&�H�4��p���{�<�X�y{��Һ>
�xB�,�,�+�`MV�b�h0���rș�	O)$�_2-tT��/N���|��<_�,c�P]�iĆ�y-��01d�ɵ&(z����G�L�N/)�,TړrT
���7>�M������~�;���[�����o������֏�Ѝ)H�������~�}�������%^Ɠ@)�#����#�S��2���a�4he �|n�!��Q	�q���l(��_�����q%-{�_�D�t��c� �Ͳp��[/%�>���xq�.S�|���h��`u�3ȼ�</��������+�]X��G��11�6�\�:�w�<9K4���$ ��u�$_6����X��,+l��V*1���(�z%�3Q(R�}נ�����j�,}&���hP�6�e�/xC�2�k�>U�BS;�ؼ"{0����4q�o3 m��� �!���*U�izsD,�<�CɼQ�ч�β���m��3�l��D��֡a��x���1�Ƶ���MHm�o����`♷�48Ȣ�6�xi�3�S����Q�pX��O�����_p��ؿ����{�Է~��}�K���2� }�����?�޿����bn�*�X�����r��,K��Ng:8�"�Cj�����RZdAO��b\�y��H�� ��n�n;�#�O ��%<4V�.���+��5�IcWC>��.��*x��"�gcB�H=�s�l6��_�b�ڬc2<�&e-��0��-xkLY��)�L#Tk�i�{YR����pd7hL��KְOȑH�m��'�� ����F��|{���9rR�����r�vScz�V|��/�)�t��~��#%w��Z�b ��ۧѢ�-V<"t:�[g9"�tڰC��NL.u�k1Y,"r ,�F^�ɪ�zg��
��"������	�)�PĽ�傛j�mL<� �T��(��qqd�c�.Ƚ�c�y�P"*��	�HA��l�=��-!�����o���߷�W���g��{���/��>�=������������?��?���Piٸ�AT��2�Cq+nW�]�J%?T`V\��+��3h_k*h(��'+.�B��p(�ou�݁��3�v@������F�\�7�	��MPR�=�,��L�sDZH�p��n�f�h��{�< ��d�XR��*�uȋN���7�HcJT�T(��y�� I�8�O<D �$�	�A1v��y0���L�0�X�#����nU�{J�(�[��+��2����xCL�a���)�6�xB?����1[T��IT"r^�&�y9�������S�%���P5 �jfgUDF�au1|����ABuI��4:$��w�E7����N	i��FӉ��b(.p�Ğ
�S"
���H� ��Z]8���b�֌�]���������[E�+bL�}Y:Ox�gZDb�;FE�'~�c������~����������Ϳ�K~Q���?����/~�O~����%sD$#��O���R��bw"� K��o��dׇ���Э�~��i�����4���@�s���J�a�n��Z| �g�Bʦ���P�_�ާT��0&�
V	}���8��,�i:�C���?�7 ��O甂@��d�8���ɕ��8�X�Fט"?M�T�c +ˍ`�1HCٮ"c�t��#����� ��fm�Yu�_r�r o���6���
a�!�N�)Z�!���M�E�b�	:LξXR	����<���64���g��g��ղ	T����l�G���ґ���0�t���6Oh����ܻ4�7?7�xb�z��neLi�q�m�AэK�Ue�J��ZUN�?��(TM6�ߖ<�i��9~���Ar�u'�l2*�Be�b�v*�	/�}pi��Et���R7�Xَ�����I���3����`y{�����ȟ���7�������_�s��ὋG��W铟{�˿������>��o4GK�խ<���~?�t?9�1�Q���Ł�ά�h���5t-������I��Q,���<�#.�g�7����t��A\�`��3*����@��ȿ�~���˞�>����Jws�p��y����J� mF�8�w����ͦ�C��RY�����F9�\=��Q�l*��v�"Ŷd�&?�F0<��*w���~���s+]�+�T��AQ�=��7(ޗ����!�_<(_�J}R�M�t��N���0]�PɅ,�u�]q�\^��;�Y��:��aGs=�E^Ȃp�c���u�V�����k4�K7�h��� EkcX�OJK0p��"v�C�]�xǭ�(w���N��k��%DI���)��U~s���z�7�Jc�t�&�+����zs�����|���������?�Mxχ��7���������ѿ���̑C�M�'੕$�����.v�Nq����k`a[&I�P�~B��m~/�����K�&�}�,(��x����,YO�>f�S�O��x��z�I�)C�Vi�����p�`^1��t�#w��C��",��������~��X�j�NE�U�Ӕ<����%Q�H<7r�*R?���.��Ɵwp�+AbP�'P�,�����l�{��v['��9h�<PĺV�AV�Y��z$�[t�S�0�k=�8��	�]�𼥉\�B���������o` L�YZ� 1j1\���Af=�C�����&��[ׇV�d5��/ɑ���Sծ֜�v�CF�2��s4�)��fC�Iօ#�+�T�%U8�Gg}�Ei �;�����G�f�9SK>ӳL�R�����~��w��������?�m�͟���<����~��_~����9����o��V�Su��F�btK��sg�An�;��D�L��ur���ߺb6����;7��:E��:���0;���46k����"��p���� �w=&����4���>�_^(ۑR ��P��?**�~esF�$,xl�;-cfu2�Ԇ�nRԩ7��^�,GlÞK�DK�O�r��8Rc�;r/����(�''k��`�jQ(���'��<f珵��0)�>�|��r�ԚK�qӘT�2�����u�S �~�@ �ۇg3�1e�}���gɦύ%���p�1���FY#u��)���Z#~'W�Pa��5�ϖ�k�MփYy���&La��h���*��3���g�커���_�;?��~������_|���7�e�3;)H��^?�������5֞e����v���XĊ�D����x#�D&�����H�H|"�H�b	��R>�$�qDl�K� ��cl@N�L�#�bl��o��>�={�=�]�U�Տ�5�����;��Z3=�=���U���������;D�Zt�B/����ZHj?�ܨ7��y4|�n�]A��|���fAR}���tSsҕ+���?]'�r4�\����E�.~S
�k���5�la}-� 3 ��Q�0���ߣ�s�R��Ygȕ����m��0څ�wICB�����{����
A"A��F����s�*�[,�`N3~9��9o�p��0�*e�J�R���)�Ƀ�C�K���c����^C�QDq�R���g�Lҁ���g8s�pa-,�q`�G��?��������_��?��_����T+�j�g?��_�O���_������N�[V��#0�Gx1�������s�r��J�ŢV:r=����7%�D�ϒQߨE(��t��\BR�0E����[|��d
�`G�C��J������$��۷��	%��:Rv�&!%�+��,��]}XWiD+;Գ&�ϿkTO�k�K̀<�&�h��`�g�![ ����V�x/RP���s��C)�P�z�'��������O��Rװq#�,Ek��`\+c9M����^���f�?-�7Ooo��am����ѹP�*D�������S]bʅ��9�"����/���_�c��w����[��W)H��F���O������IP;�:Z�:�)�p�P�Q�fs���\���Kn���-b��Kd�OI� ��dI��';����R��a�}���'��T�� C�@�UdK��-=QRMz颦h�o}�?�Y�s�8FAC������_��]��e(\wn����bUu ��DB%ǤV�j�O4*��6T�/�\�Wb}�bD���/ܧߚ�s�Y`��1�[B����K��_���Z�5n���c�D�P#šQ]2��}g�1̿����#�(bQ9嵭���k��i!�qC������_�¯��������/����[����d)�b�����������O��w;�+vL[����b�i�`%�N1�p`l��K��dZ�d��[l<����h	�ɽ�D9fw,�f�D�Q����$�8�M�Y�I儚��$��Z���
'�۽�����ncl��|��f$E$J?o�/���4�ߖ�t�_w�O��$�q�o0DvtAQ�u� ���\�Lڸ]|�4�]��ӵ|Ša�sx]u{�N�����9�Q���"�ݓvD�j����*k ,=�	�y9+x�*�8�vu�x�4�|��Ԯ®3}�nf��b�:���Ub����l(��_����=d}�)��?�o}����������������,R�~�>�7}�7}�_��rdO�7��D�,�kV���yiH��#��<��
�LqF7�L�׹̯���'M�-�ϊ�g��FR�*@��Q���� !�`�[���0o`w��דB��.�E�.DR�c�(��GH[;�6�zY�L���E��3�*��X�JyY�x�R�+�%"6�c"�D�kj)��$��#fkխvHq-{Pj�| k3V�S�柳V�g0Wy����q��ߋ+@V��f��$|[�>��b�Ɛ��YEM�?87�ٟ�����HCҵ�/�O�7Л��.<�� 7��Z�R��������O~�����������F��V�~�_�U��M��������tw�g���E�S�B�����JG�ȺعrdW�]8(��v��;�����B��>R%�&���gY49K	����hpz�����]�3�������y�,YY��{z�)!�C~Ϯ�L��!��-����In��@��E�"�T*��TA ,�S^A�\�z�r9q���}4�,r���K�~���#��F�Z�d�|4|�l�,Qg���4��/�vfa�9��ff�����b��Н�0���:�m���?��&�	���@2X�c�8A.0R�2�Q��M���(L�13^��r$&��gY=�8�l�k���T�;��?��'������������n��C��_�������-%�#uB`>I��,W�A�m���8y��,^�4	���W�^ ��^0+K�������\��8��R7��bsD�	4�Z���4>����_aC��U����iif���*8V�*Q�5[�Rn����{�u���k!�T�t��ҋr�.E
�E
�A��^��Sy�&(M����h{�F)G����)]L�� 2�}=[\P>���K;X��N�[����=H���4���a�ǃ�=���Q�~���T�k�N�DjG��NTe�F�"�M;�Y5������Ky:�-%��-�����zq�����o��?�_~���o��_�#t�KA��������ۏ���T�����M"]�C!�H4n��S�eB�p-���[0�������X�IA��������O����i3�JGqEZK��w�)Ո��1�:U ���'8�n�N�'�@*Y� �y�Nk:J�sk��<~e�Y�.=���u!�27s?�����:��p�w%�H��cR�[�V���]x�o��^f~!'��X��upp� S�g>�ѯ�]������|�����T���_���~���ov1�e�_� �EEi���Z�����|Ɋ�v7��N]���\��PR���fע��b_��<�����ֲ�P��AY���胳�^݈FV����������R�Tq%��`��s�=�u��P�U�0��h��(_����={ɼ@�#��ZE-e�V�&
�.Zӝ��5�V�L���wE,�:�JF{R)�"S>�s\ٌ�hN/]����/TUV��
�W�si�]8�w�I:�#�[�����C$>~�G����}�_�����o�~W�_��G_��~��|�{ �L~��]�82�ЭÖ�7�*�&.0t�Ko�*=%���1P��_GA�,l��F���$|�t-Ʌ!�LPN���U�v�\~��h#�Z[oA�Qn��)I�q_k Ə�A�J���R�s��,^c�7�ML�4��L[��u�Oe�����v���k�=Q�Ղ ������%`u^��$���9r�8�����) �2!�I��};�{�2zˍ,ݘ;kZ�����)�P$��'}���j��Q�Km>`}�b�#���������|՟�{~���
ҿ���o������� �[6b�ohx�e�,y����\��.:O;$+�=X	�R/iZ
I�
���U�˦7:��6l�ԍ�ja��rf���킵������dFsO��<N���RʰD�M��؅4��j̟c�aB9�4RBh�Z��6��\��tk�)�Ma<ҥfp���}�VXʿ��[��.Y׳q�*��<ϔ�ptve��s��[B�v�{bk0�(�>�N���b'�����w����?�{��� �O�����c���{�%Ț�N�|���i��rJPPn%]l� /	��ƽ�U�`S�f9�S�)�h�jі�V)e��KF�v���p���������E�/f�+���|��Q�m�A����E��k��Es%Z�𡐏�_�[IJWAe��h|K ��x�8:,�xw&p�dA��UW.w����Iq=���W/�"�(�Zz<ϋ�KfH~,�_����!|F1�86V�t.���+���Skm漉��<?�w!T�� d�����k+U��&��_�D�낒:F,�&���5V`�i&e�`ܺp.��t%뙾G�L|u��`ί�@�������[�����E�_���u��CJ�׭��%�K�3r+��>��@d�,���-\�Z<jN���e[������U/v��ٞG��)	%�	��sV>��0�����b��F/rqD���b[`;Z����cط�*�۪G�ii�b5�3�4!Ž z�Hm�B2s\"�u�x	ۍc.�s]hP��
P�w-s	���|��QX+\y���  ���!�, ����J߹
ŕ(:H��6�Ҕ��ЯdE e-����hg�����۾����T����������t��U#;�m���)D-����D�������t��`7�m�����Xw@}�ʆ�1���KԨr� �0{��{�c��kjݚ�����o�\U +յC7�ϯlR�6e5A���oR<�歀ի=�\���,�#4���G~�'�+��$�sez�xL�l��v}���o,�4�u^2J�$��6_��*\��6gd3��i�I)Oz3ۅM�PL�����W��A�;�ʄ��!I�o��ŹK1:0�����TQ&�CRO���Ե?-�*A���?)�����؛�ny�����˸�5����>].���w5�o�����Y�����z-w�������a�ԣ�邇�!��*j�x�J�!�qX��]�1���q@��������?�S��p�F*�	�,gV���X�PATp'9�xr��c�������*��cŬ=?�ή�	t��(ʈV���Z(��N�*�����Y�?,�s~��?��X�Rj������������K���`>y�*�<��Q��t�g�/#�Cwl�U��ZS�0&��^Pbҹr����K6��`>y��8���)H��'�����)�Ss����}�7�=���-���W��(d8�q�Gz�4{k�й4��[����z��\��~���S��rĂ�{	���TF���59/�!��Q�z�b9�^���˛��L���N�PN��֬ǆ�hMȄ���,����:귋�}�͕����,-o��ҕ������<��]c��~mL����V�����/kSi�
m�w�=�k����
h���ؖԇB�Q<��s�1�
X���2,a@;C(H��~�>���j�`L�37�����jlv�8-:��=��F��#0�n�-iH@1����@�=�dí��]#���a�^נ����X����C����X�.7����:4�n��UIи��ta�}�܉' :�s$%����y��I����BD��x��P�����������[(��ޡ�hY�V���4�3,Z��20ϗ[�ﵟ�5��e3�d�ڰt=h9�����v�	���P:���2��M�A�"w>��P�c-D��G���B��t���n�?�r������wk�����Ũ���k�{~z���$ǃWOl*_�����?�h.�lK�t��uZ�R�s&�U�#ΜQA���|������~�;��~b�2cK���cɈ
�/�Ch�+��P�.��&��f'�+OI^���+~�+&>/G9�M�B��n9�������Z���O��j����G��
r x� �,��u�[����w���[|�����a��ygK�*e]�0�<�vm��䍙;�l�}Mv��|v�0�k}��� }�������頾�v2���pϙ�:#H��3y�/�x��H��=����aZ�K�EmKaMBzF;X��*�������������8��\�����0��
�z�u�t/�?]������X�o
'��gĊ�y	׶WA�B�>��=7����}�_���@��?�z���!�5$�n&���Nwa-��
I�K�i}��K�{��80z�D,�^���ai�ҽ�U����6;D�c������{I�N��<c�=
F[��ǝ�R�w٥�����̯������Ѣ�,���:l����X,Sue�LZ&dU���}^&�B�St����;��
n'��wA��q*��R�h�� h�rp� Ǯ�{��1Opr��l1K��9n��9=Nׅ����t��]Е|��#b����#�^��p�&�vL����m������h%�������׹� �L Y%@������u�ޘ$�����^�����	Q{f��E�熘l]yL�v�����nx����`O�v��b>�h�����k�~��Q;��v��8d����?,)G���l��x量� %�՗Z�k���o� ��5�D���z.��p��eH�ے���Z=.z� ����"^�
^�TX�H��Sb�̅.���n��Q�c;ɻAI��]>�o������
ҟ��O�wj ��~r��r��^*M+l!����-.�����������H.MF���Ч��O��;��"�v���w�^�A��۴*/w.g��_nv��`�C)�
eG�K����-�)�՘���>?9�1s�ͣ�=��	�}�r��l�"�]�j���Ӈ���������}�;�pE^_�Y��$�|^L��8>�R�y��t�H�*N��b�=���r��\�}X,�=��E��?J��P�VUD�4�A�V��,�b��zD��5KH��{��>���̊ʳ�\���m��[��w�0�4p�j\B*y���N����Jzc_���9�Y_�[0�c�Ї��c?���I1���M���O����X8o��.�ӌ-fȅ¾�X$`w���~
�?16����<87ҍ��+�]��E��a���S���(���R����4e��H�YP�������v��G�"-6�>��>|��?�ݑ�/��#.F]~ ��߰���É琦6�k�M?�.�(0�VpW9.t[SgLw���9մ�'~��ܒx�=�Lό-�*����`��a�k��JB��P��N�J��V��RF�D�jw$Na��.,��Zφ#a5o����4%�F���ed�FK-�]L�=6Ӈ�|�iX
D�Ax��{����8{�����F��uq>ђ����I�=�ӏ@J����� �Kw���4��;ĺ�f��A��@/�3�������b4\��̪�`Ҹ�O�_�d�&@
�D�j�"_n�7�%e���2��iޥ�֚���Fz̾䏃q��Ҹ
:+���؋S���ցɄȮ E��x�-�W�ZFT��7)xG�����=����W-��_�UAԏ���(��t ˟s1~��!)R�	�R�\&�G�o�]�D�M����cH�<26��#�	9;��f�q�4����Z'�t �bV:[��[��9���*ݏ�O��#Y'�?�J�bZ��((�N$��𶆒^}�c妼oc�q;AL+s�d!���V�*]\ �Ud
�A�]XU>X��$�p9��O��/�-�Y��R�O �r���f����592��6 ����bSڼ�.Q�AٗRuy	-��u1��;�y/��=��4/ܡLw�٪��Ud�tu�X��z��}?^z
�?|���rwRhm~-����������t�ьUr �� ���-����F��J'�����鵱RP����ӂ�s�i���Z11V�\<��{6ڻ�r����ư��i0=�W�Lq#�"���GD��j(�cU_���<�������N���p/����E=�i��n@�2�}7Sp��K�TG��5��6������kU1MO*C���[��G^'}d������w�4N���4�YF�S㎴Wk�=���[�{���j�����_���q8m�Z�s4���/}���V�2t�wa�.Fa~���/�»Z:y#�M������сy��`��w@�z�*Ǫ��9n1 m
X�
�}$ܠ<�E�E��y��E;ǆޗ�]��]
����ǯ����L.Ԡ.mh����6X��=�%
�2���_Z\B8�j�A��֊Lɂ��L���; ˹��=��m�+Op��a�Rh3o�X��
L7��qd�,)D��gT��ڍ�c+yk�x��p�l�9��l~��O�RQ��+��\���I�s��{������|i��������T�L9z,l���9wӬW�\��R��Ԋz���b\G���#��}�
�����̯�܌j�H��A6m��ߊ�}H ��؋���ԣ�m��|\1�����",�c]��i��������I��Q�����C����@E�a��:�,�2��Q�z"�J'#����r��5O>-��N��O*?=��d�LXJs�c�a��װG�3�@��hX�l"���L/\(a�aF9&O;��$L��؂:�R��m�"饲������3�B���ц��Y���:گ�	"�	��e=��殺X4�,��T����՛V7O���]�����Գ<�A��5^�[��h���ķ�4�}��{*����m-��4u����#��.�ꂋ+I��7{�R6�GP�y`���{���MsӃ'7,\;s��W��@�ZT�Ϣ�.9ӄ����CQtB3Y+X�;����|2�ǽ�4�����)$:�h�
�F$� �{�Qna�شš{E��Ș��#�/<L���d1�Ƣk文Y��b� �!)I���hW�1�8�ƻ���c@%y �	�(Ckl����s�Hs�{.���v�_���w��� ���r㏂f�wD��������Ln�A�R+H�3C�Kx���N�y��Q�#g��P�׽��<<f�a���O� M��5���a�]��.�q��VHb���V�@�,�ھ�3l�B�[���0zs�X7X�&}�a��Y�`�B�+i���'ȿ�Gk����ظxO��������<�{2
ɺ�*�&w/~���z�"�Mq�vKvv@���(HM���4��%�i�E;^��*2Y:2�Q�qH+��}����%O�����*j{P}�Wd<�v��<GO{n�����5��>��֢11'N.)g��w%Z*�Zˊ��½����e&�xsZ��]�|����@�� �t�}6��Q��0iݷ��	o�z.��8D��@�q5u���D��*$m���E(ua������UFKW \E�x6a��l[.��v< ��Wx4�%�˭�G����j�_˝{��5��y��O� �CT�dnYq�'�5r�b��9Ϝ�s<��Z�J�m.,��
��U���^��ԡ�����|����o�jX�f�I���Ӡ�E��G���d{6^����Y�9v� a�U�y��Y�j�=z�����-խү΃�
�c���x���>�������_뽕=t���<G{J��'��D!!�y�Hw �9>6�^J�{[A|
iP�J��X��Wb�յJ~��짹��,�M��VM+d,t-6QJ�o�T�T�~`��ֈ�.�YVX$&ac�G�a�v���M��6iSAC�P �l)�<��Z!�af��LC.6��K.��r{B�^|X�'�@~��L���,/<%��*��kPv�yE�ށE��Ｆ��#Z���ޝ��(��e��O� 鐖� 	�$�Ȥ�u[]07��B0Z���a�"_q�Μ.�4���ʼ�k��/a�d���ܙfM�ow��k= �D�:P��y���l��##��AM8��ppY�MJ
�6}�j��I�J=Y�k"U�����UE��e��֤�]o�X�I��ҕ3]E�M�MC�Ɲ�����x�8
��.A��[���8�&G�ܜ������ߠ�X,��w�G�4JD^ėX��w|��H�<���}�<�~/���O� ��JC?�������ܹ���R���U��(ˡy��n��W���Y��]�}�U����N\}s�ȷZ�ݼ����V���^��9���	Mam#�f�\^�FX\�庿Y*�45^�a4S	��uw �0�&CC�+S�@s��m��=�$
R�/�	, !�T��ET���F�ݩ<�,B��R���R$f�Yɚ���2�f.q�5j�w7�����y��Ҍ��!p$[��)g/a�Hma������6�B\��N%��P]��T��t���Q������(�w�r?���<qw�m��ZH(�4A�����u���>UZ �Y����jf��HH߳ۏ��yF9�I$��"!-Y���@��{�/����ӕ�@��B}��	�����{��F�YQz2I8��\��C��D�l�p�
�zy�M"������L�/��j��c�U�t�G��
tE2�u�Q��5��\k��́}v��r�n|��jk����5�f���nO��oOy���z���L�|�eoh�.]8zh�~�єsZYQ/�iٸ�6_�4�Co&�@h���y2j��w�.q�����2�T�Q�R.,�����ϫ|�%W��.���Y�B�`�����Ó(H|��6�KA6����[	����q�y�n׷���Q$��T������W�hOD��0NLb��Hv%�
����Q�S��T��j��C�@�pK,�|&�}C��F}�"
���uTE�l�6y��HјJDR��(<�\T�Xl�v?wҎ(��F�6A�R�`��"+tR��5zV��o@�D򑛗�O��U��Fi��uV���1zb�)X�Ȫ�LϪK���$ˇ�A�C��-(������.SSl����\Y7|ᄗHN���-)]M_��;�/�=���4ę`cǎx����5U�TDE�8*�������=�c���?D���˭
y	�w�!��:�'ne���*�'{��t8,S
�Xx?�}S�1�]���ߟ�P2��z��
��2�u���ueV�r_3bE�g�A[@9��}�f̏L����~.�m�V��l�@2�w�%��S+HZX������x dј��3�H���Yj��i�q��H߻��������q�>���ׁǐ����0�-�V.d��TU�-ɺ�姓��y��/,��
�ۼXi�4$׾y%�;�p<��������j�����HSK��Q�N�A�!�1�ޓ�DClY�[��:�zP�ZɗKGb��˳�����������"|J�!j�m�MѶ�5��i`+�rw�B��o��n�q�|�rz`V��n��V[�S�{G�&����ؖ<�AW�1cUZ�	��U
ol���#��Xmt���{ .	:.=����G�y�p�F�t���
���Kv}Qn��&#� �Ϟ�����h>3薖0|'=`��l��k�E�=0���6k˃�kg�h�_����/0��&o[D
�L�3�T�J=U���>��x�>[{�F�c�8�J�~[��W6id�]RQ��Pn$5��P��
�{׀�}w�RA��v�3aVeL׶"�Z䷍Jpe�M?��Q������`�{Ğ)lZ旓��NiNe0몰Z��YE�HW�ԥ�,m��MŦ��=&����d���Ao�s��4��=M�XŢ� �׫�DV����\Z�%���zM\)U?���SƋ�8�OfŖ�Mo���(;]�u��x,�4�Uz�-�S~�્���_s�7h�u �٤�6Չ���>� ����%&���"P����9���ק2��4�x+����_���]`�b=[ ��Nmi�/�ҙH����)�zTmD�pz�p��=��tĆ,a{�(��b� B *�)={�&K�1S��"��d�k�t��\⓻xk9�u��,��C4���&a˱}�%��V��7��V.(l?�P}V�qA���tn3��t�m�D����v���?T���Z�m���XD`	t	��B�X��`8$r�(�8ѫ�ݗ[����ͱ����8d$%,$��<�&��
�T��<���a���I�51�}�����rmӅ�S�����f--���A4|}��v���y7��B;^��h�'�)����������A ��A���P���U+L����?M&�v[��l�D��I�r�L%��BP
�6�ף�0�cE�V�m+�V*隅�h\q�&���z�U��җA�z�j�n�/���y�tYRN�|)Jf[}�l��,-��B�6w��fzZ��}2��B�Iu�آ��W��w���G�Q뚱��#��duѰDE�w�_$uQ�9Ev�������t��s6�A��R��6q�)�%w<|��υO��*��	+��y=:��E�w������߷X�4[E�#��$�V7}��]�j(����CX�;Taz��gYu_h�� �1��~��:��Mk,��U]�=B�fUI|��"0��W����^z���K��)�6�f[�h|��k�����\}f����{���4
�<�A0i��y� %�d� ee#D9'��pr;�Q��ڭd���˂���n�a�����t�E���
���Ki�]�ER�\�@������x[О�m=�� 8�S�>� �;(E��aA=�%8��h��Y+*��4�ƚ��[���h�>��q��'^���R����/p�a3�\�_�v���W����q�7�д4�9	��*؁S��"ʞ��*��(.�_
��������\l�⼏g��#����L/H�Cμ,��W�8�
s6�"1s��J���y�����p��bN� I�_�<U���^(X�"{v0kpC�l��_WL'�8.��A������[��N�՘t^[
%�Y*5f���J�Ւ�a�o(�q�3�![��Y�)ݧ{��ny����D��XA1���I��Do�{�
�=y�0KY�EC�=�߷s�,���:v5��ZA�ջ�PP

���'��8��k������> �a��R��KW`��$<T��/������9��ݜ-ZQ�2=X�uMj�\��������<sHz��u��G�4
Rir��jB�wJ8��>�C��/��F ��Z m�Sy���f,E(���*?�+�a!�Q �"�$$Y�zg�l���.B���b\������m]�&zFkC?�30����/���RT/𨨩�!�'�G��'��֘���a�z|��'$��"�E����g��2���p�}��+�:��@PK�v�=&��H���.j�i�7��Q>�Q�,@�Gop����r�
}�0^������bG�d_���S˓W�L�%�x^ݖt���h(؞c�����1�=��8��-,�?&dk��Ҏ|��/��S(��d�4R�OY�߹`�-��/�[Y�ݢ=L>�.�����{S����cZ�}K�<���ik��ȧ�����ilW�G�~ۭ�Ɲ�Af�G\I�P�Σ �&���U2
�h{�]U����,twj��2�pAO�u+=QMj�	�?��{b�pӍ�y������u7:em��^�>��dJW�[����Mf�9j���2���+���@��Z~�a�ڌe��9��⋸��4���Ů`/h%�\�L�~��$���+�mk���`���L�7�4Y.l��;�O�uɚζub��}v)�!0~/�|-IB�ܽX�?�Œ*��*i�;��nq W$�d�5Z�DII�7�u���{����x.��<
��ۚ:<�}�7�b���M�3_GU��4ڍ�'�]U��Gm!�.0ګ���{���at��DKb�U�4��[$}��V�У�6`s��8���u㱓�����!K-��$-��U*�I��ʠ�ù�9��[��o8���h���с;��9P�3,�.���WF[�ڄ3�,�X���7�����Jm�Ħ0���ؼ��^����z��y�P�d����LOG�h,+HyVw	�C�d�(�� EM��J�
VK4�-{�Ck�m+Z��XOA�i�~�s������3��WW0A�VG�J�77R^�"�+՛��E�Ę�FO�7d��@��B�LJ���J$E�NҌ��<=��l
�0]{>�����kӘ�Ҍ�?`�d1�Oq�
/�4!�C���jV����f.���0׏��I8��G
^Z1^���0��wK���}��yl+~~Q�F����6Q��5�Ω��r���5�5�U�m<��z?���K�@:)ש}н�U�_\hƉʤ�5�����w�/����[i��j7^�t15$��% ��V��c�ԣ�8��ʠ�����K�_&J`Z���6���e�_��G�u��3I��n�؁���B�PA�OŌ.���4e� o���N���w#!F�lC���BH&�����,�2�׷�aj�(�򑼂���c�Rǘ&���f���M��G�ޅ1a�:�V����75(&Ҡْ��q����Sd�䡵��E��Ԁ�%�!U�t���a3.���J��=���.��x����q��Jzdi
��yx���f2�qG��{��O�c�8�	��gFI��Ix�oNb�Mo�>ۘ�>�8��:�"|�MM�ª�'YtS�T��?�R��?"�}'�jJ;�Wh�@�&(F> LN�3�Q�b>����Ok5���[4�_���q�ၞ
�G��kT�@��]i���T	������ ��=��V^�n�0�a���\@S.�]��r�F-� )Œґ
��^G����!�1�W�ƞY�()���S1u���!�Mi�!�T~=:G�8�s,�� ���c7�c��A�"�p���,j�� ���[mvz��kx�D��<N���S�vR����w\!���#)LaU��`�8S%���KG�[_�ﯰ<��c�X� V�eE$�Ӕ�IA
��b����	7<��T6�wY;#���_޴V��k_�
�U��ѯ�0˷�KtP���@����~oZ*W�S�W�tZ��7J�*�r?B��x}���"�W��*��gQB�Q���1��l�-膭3�J��>	�a#�l�`.U^���&E[f��v��2�gnS��]#���B�SՊ��_��ir��d ��]'/����{	c�Ol7;X>�D�h���$w�M�q���z`���1��V?�{��.Wx�}���&w�#I[?����cS=&�Eh��"��A��U�pM����'}� ^��?�0a�es��aK��G��fr��!t� �zf��� ԧ6Q�ʈC�@
���%��G��-���xw;4J(|7�1��}n��7+�X�~;ӕaȦ$�K���J�zV�$`jerٿl��'eJ���ti���i+[q���Bb�ƭ�K���a�K�~x�1����%qn�8��R2����>�%��ϣ)�'kx�\cV��v��{@0�ū�J�'4�&Z>~��~�?�O�K�6�м��n	9˯1~fv��6d_zJt���3L)ΰRݐ�1q���,Z8�$X�ֲ�<�ԧZB�M~�$,�t�B��ۮk�LƮ�@�7�݌^Q__gei��%*Z�2;���eX��|�jcir,��1�� �R��ҶZ��/�6@8����^^��
x7;n�E��{��K��P��z���6('���[I��i/����?��_�����H�/�1P#G!�+��=s1���x�Q���<*ʹDg�~�I9��7�	��x��d��BuΖ9N:��7�B��Q��|O��㚫��+�ngQc\ث����%~�������6��~A�9�G9������0���wrior^��DZXa��9���F5��8��TJ��g�����'�B�x~�^�W�����7|��}����Dw�`9���}�Tue��-�r�����������F�J,�RԪ�DӰe��Ё`��@�	B�"�5���V�&ZAҴ���P铛�$L�Q]���7�#�s@�I���h��Y"��b1�(�Nt3�S�)F�����K͛u_�f���ﮙ�ق�Hcb�0������+$�R� ��3qһ�����T�jB�7������GXI�&��/���˾č_��Y����d²v�I��%h��W�?rԄ��3.	e��~Um|���Mhuo4�:����}x���� ��#k����`�_�Ig潥<1W��:MZ�5KI����*�e���'|k�Ih�����e�p�Fc�����S��wG$2M` ����院�����@I��YL�%	L��������}��^�>��/��4R�H���Oxu^c9 )* pP��Q_�Z�h��}3��#w��b��3�5��
7�ô�{�o�?L��6��_�	o�^���AA'ㅯZ␾UJ���L!�5�����9�o9,�-��%
��[��bLI�$�e�y���r����S�}p<�&��sƀ$,x�p��^ߥa���`,aW7�|k�9�cd�䙮d ��q���-��ͺݙ8gpw��$�p�O�'�0�������/���>�>|�c?�N����3G�c��<\jY�q<�ʱt����	S?_�dd��I�c��=Y��zN�x/þ	a�x��+���v��|�!�	��	CXA��/�R>�M��:���bU�~��f�-��1�н�������q/���lчIpu�H��6�x���`C����j��<�\��y}�%�6
�đR���{kT����e��E����a��ml~�Dc�ҽ��/s���4�SR0*��5Ӟ�*4��S��ӫ��K��m���9�4��<�?G͜�E#템"�M��39��_r��:{&�;ڻIJ�8U,��J���J���畕3YD�q^v���8E��J��xzG����}���M_�ܬ��|ɛ����ƺy������� �3a]��V��v 
w�)�`��r�$����
奞M��Q���#�8i�k ��dH��Ya/h��椱� ]t<ɑeŘ5LnAT�	CۡH�ҫe����=��0�-ބ�Ͻ	����!ĭ�]@��Ӑ��A~cI�l�'�X|s#y6@��vz.���_�2.����}l��5|���W��c��W>�ۥl9;�` /b`��̮��g?z`�菥!t�yWE.��h���X�W�f��l�Q����Q�>�k!����v7L+\���&�N+o�N��n��J+s���]Q4��%��٠D}м��![� �9
L^�yk��om6)៟�dL{���KJހ���$`)JO	�[+�F.�ob.ȟ5VhBP��Xk��]P$��f++~4�)�F9!b�K���X.���d"2 �ҹ����d�^B�
�a�;�{H�D� �|��{Cc�^��_��5�Y���� mq����qB������=f���Y(��3�P��3����F�=A�@�t��d_H)�r�E� ��
���#��e�I���x�F�L CV�s~@酎(Gd�%�he�ʙe�zV�⣼J�ڢrl��U�fڣ5�����J����Xa�{uqE)	{r�7�l��� h*/�x:�N.u�B�9�!�a���w�lm��joJ7|�]��>����")����
��V���TE�5[�,Z�
�V/����fښ�M·[Ç�k�~��ˤc��8��;CPV�����!��*?�ζ�ܣ��R	�D]���	b�l�G�q�t0��/0�s��8�wp�n�m���W��j�k3S��:Q8H���������Y��F�YLޗ����O�������(H`�vo=�Ѐ޽O�S���˥�ެ�noDF��:�1��E����5l�u�pn,��S�(n�&9p��u�Y�;
j�A��|Iu�۟������I��%�7����E˓�;v3�(P�nNXԾ�p�e�'*=cHi�%���?��3{0AZ��mD�&+7�r"\�7�?�w��,UE��'����h�OT�m��/S������;u��IE���
�Ҹ#CD|(������?l�u��Ig���p��Ѩ�!xL�k �k�G�ioJZ�IM����J"�ýq��!tHS��!ǟ��H���W��2Z9��pH��eq�W%�Vp�Ҝ�J�Rc*�KnZ��7̠%�z�C�>r�8��d�ru��a�@�pg�:g�(�7��j	�Y$���Z�#��yq!7���щHIo�O�_!��4N~�o��22�|�	*�ʳ�Zy�Wh�ji��� Jʓ�b��H���usv�*��W���<�a(GQɦ=0@Q�VCHIB��Cl�(o-Fi��l)��D�Y���`ԘS�!�`n���_pz~�0\G����ʾKtJ0TEU&�H��k��j�(	��-�����g���>�y?���1f��g��;EP�>�9K�X#6�2*q��-��])c���s�1������.���p��YCk?D�:%ؼ��J&N�i�Z�ݫe��N+���)�,$k�]Y+�w;�����D�+HS��:�Lk-C�X|ZT����mr=�!��cSd8���}!�rk�o9�pmH��J`stU%�o7���L��!����v����C�s ���!�зY�|�j�Q�v]�o�	I�����SJ��1 �a8��8$��:��W�1Ȓ� �����e�q	q_S:���f�+4��T�ͬ��P�9ӻєM��Zus�g��n�;�؋��lA�j�����a���kj�Vd�T�%=e�w�;\�e:�$R|�.�Or�|a�1z�\KkG����+�61��|�7��������R=��j���pa� �C�N��g����L�p��n��Y{���@I� �,MgKmSX�����0�k���о����0�L$$Y*܍�=!l�L��x��!�=YHL'+Ԝi�
@�(O��3�L��R���>^��m���u:�e��xn�֚/$8��0Z2��!6?��/.��Ե�¶�3{� 6M�۟� ���Z>�ڐV�<�q�3��u��[��� ��R��J4@�S�D��{�������b"s?"!��Yn���6p2U*%�g5^k1�~�l,Jf�ܺƸ�*V+�E�@U^�v>�蟙��������CRc�Q�`�-*��Y%�&�j��|��:������0��k�4�l-
k.��:7���t��F2�R�)�5?N��y_�S8��9�TB��=uh�}Jن�9�7�b�,8���ED��`
K�q���?�/�G"��Yf��Џ���Kr�u�D�^_�6!}�ճ�&E�ҡ��xb��_�X�!A�
Sz>��J��$�#�kJ�2�������̜����Z�AݙZ��{���6�*dZa�K-�O_�a#��CM�&
�h��2܊GR1��2<"]���ZF*@\OJ��
�B)�ZU�az?�&�D�߈� S�vLcsI=�r�R��ޫ�ig���U�dRVq�Y,�^ɑ��=H1��̣@]8�t���� C�.�Cy�/�@@�y~�$��:����#38��1Q:��P���*�%�t�|%�xX�+����>�ȭ����j X`4���yGP�����j,�Bb�y��Wg�O���Cj:;iQ�
���n.`o�^v�m�����O���U�M�`wˣ���"�T!��|QSJ�����2&#�� �TVr�d� y1`Ng�&��bV}�;�g �;�G�6�	�P��a%�<
��@W7^�l'�Y��V��)�^<�+ /�9��1�j3���qS��I�2��O��M��x:Ϋ� s��C��/����^��;���OM�s�|�=��KJ@����	�8����r�s�Ajv�B�&jM
��̝t=@|�z���c��gY������1͏�VG��.<�߹$	Q6�d7i���.z��0�W�ԋLeG�G��O&���U��2f0�X7d?��?ޥX
.�.�v냅f�iI�t������^CG��x��.�.��(ڡ�5ƿJ�22���w��O]t(��X�d�x����U�fI2�{-_��0��߻�+�;�hp����0Y��(v�RENB�вڇ�R��e$;e�}��Ţ:�l��H�k��B���n�hC=Dy�����'�&rBc	A�b��g���lV���9a'Mh��|(-!�Tڪu,�X&��BI�%t�!���	-sF�V��%p��&�nb����線j0��S�%�!����2N�I���[F��t�=C�ք�q_~ih��s�ju-�3l�ҧ�\�5ï �x(G��>�����~�5�����wn��?/��IP��ϋ�*H}���j���L&���� 4,,/<;��AJ��.xuRJV;��V��υ�%���QӴ^[�M+ё�%��3���\�^�z��8Y�!����,!{�,ǧ~Yo��GM[e�?�{�зYk�=ԕ��i]���Q�mNJq�Ӑ��"�C���"���m�٭�eٰqQ�c(\_�Ъ���*#
�B������#$�U��J+R/�"�,4\xR�ZA���U3�'c�� ����I'��
�(�������&�x��Ʉ�9������	�B�hSdD��1�+o�-O��V[���8SVB�e+$0�2�1]}�!�~�կ ���Ng���W"������(�f�<��U�l���U�WV^݀>�_\%.>��h�6����$��ќ%�b�=nA���Nc	����?k&�\#�NÓ�|��Kt�����j�X�|���o[?@bUUc1�� �����;7^����2�����ϱ��}4���ȺIg
O�n�&9�3��������Al3�]�V�,�k\'�C~^��z�|�t�����:�� �ʇF���U*����V��s>�����;b8)/W�e�I�M�a�'��1��N��8D�	���x�߼�Cz���n|b��@��9>�4y� M�yh^��|F|gM�1��8�y�5��N%v-��� !�d��'5*	*Oq���J!C��
�;�J���C�SŬ�
��>�3)r
fA��~
]�HI�ԧȆ3T[�.��#Y�+OAzF!�j�d�H�A�P�n�H�m�O6��)��)��o���/���c��{R�������7Y�&����J�>�@��ء��� �dTP�?3�-T,*���]V�{�()g� M�\�(+�y�|�@V��r�3z�7��2M-���¥}KI��⃪:(�Q/ԁ�C�>f�����
�r��aF\�[Od��-,��6�(`�"�}plg�[���\��b�~"�u2�.��&�[�s�����?�1�f�gL�4�F������ыK%�-��j�&!*BKDz�8F�K��x�a�*6j��ұi��1S�Q�a��U��o厝J�����H���ܴ��B'��Ҷ�rjGB��4Y��x�H9|�=����y�K�r����t�W�w�>}uyK7���7��k��(u�>L�t#\l��e{>�`�l ~(ξ�.�ܰ�\x
I�?+4m�zή�0A�eݑ看�a�%z/�s��喹h��>���W��T��B�g{5���>[����q�4���]!8�' ���`4��J�����ۀLSH5�x:~f�t�`}�44n��j�LdW|L�Kտ��\P��
�i�)�ٳ�A
�Rc�/��ҲjL��Ⱦ벁=�Y�8�� $�@�����U����B����ǅ;"3��Ps.<��$xW=_�k&ӕ�p'(m�g�wC^ȕ�� ������˼���8�0#2E����t[q�\@ɂYd�e��L�k]�$�`�2}6�$>�1�A)��%0�4UꚂ,�r&��lC�e�M�Ի�����d/���4��G���ڽ�l�ׁ�cXi�����\S��%9ڪ��A���� �mF�]�)��{���;1��-3Vu=(у��*���8�F�C��p$<����?�1�\������ �@�d=;��4�-|�[m��E��G]3$'��5�K
FFO9`�"S�v��{YJ]�`��E�y|�D��lک����!\�2�N���=p��7��2��[�>����oe����N�V�U:�Ǌk�:������)�s&����$6��Hcd#%.�ɑSZL�0@)����"����}@�_��ZX�4)^M���?�ܢ%�G��>���1-�w!hJ7G�yӪ^�@Pc���vmB�YE}2?;KWkC�Б�F�PW��}	���=7�8dr��c(A�!�N|��[a����vt�jaE��o4m��N��9��C�@G��l�o:[��/�p�W�{K����j5P�ѽ�|��������,���y��I�@�s�|���,�,a8��2�iKaV��t�oC��s�����Qδ��6漆p�5�x�x�1����fQ�x��������J.��2�훔�
������*��\h���9�x�n|K?������$���+K��?�K�|'�:h����Ȩ�S��>�\,�����fȽ�P
?�u��������KRU�-��۠��K��(��;�O"+l��]��y�&~����4be�:�c�w9����9�������Z�n6�8��1qGY�dX w:�F�f�o)����|k��y���̿����U	�&�j:�r�W�~'��W�ǢR^ܭ��{����=�y�v����M�Q�zdˊ֍Y@�
�1��[��iV�.�{�j�l��Q�O3}���VD����&�����x�r�#L�r����ym��{pNl¿�_�z4���O��,�ulH�;Ҳ���D�Wđ`!�Px�P~����-4a�vZk
�7VE�.��kPz���b�۳��6u�.)X��z_nHWLW���$Ś��C����}VQ�$ &����+�ݡ��Ѧԍ�u���Fg
o���}��6?���O�pga����ot���)�T�SZ�p��Ë�`~=&v� ���=�J0�U��^�wD�4� ���oer_��z�����5�($X`�X�������cY�=�C�s�Hi;V��Ā=��<��zI��0X���eiM�����4��O�|�R��D���,y@+�0w�"	rׄ��5�� Z�J
b�)r?�!D�ҫI�Q/����(s�����1����+3�L$?��F=gp�=I9�Tcp��L��	�16Q��k��2Ť���L�S6��K�v�}դJm6Z�.��o�'3��J��q�/��>kV�z	W&)�2��[ ��3/<  ����^�g���FAj�5k�u��f`���Տ&?f۶�E�.��J"�p���B���>$Z�}^!�\��ߥ{��U�t7�wx% ��Y�')�)�1�=�?Wr�����Ŷ�ڰ�@J�tg��$�@��o�}%�H�u�2�
�h|�P}�r?��=n`�{��Ǒ��^�G/#��Q��2�~�)?rގ�����
)o�G���Uⷬ�������F-?���t-�ʃ T�\����7̆�m�_?�4y�� !Ec�c���"��"�x�/ո��p`^�}���\&��7�G�_z��^�Q�)41�^\�c-�(�+U�B,ң��ֽ��E;��VJ=Q�`��i� Ѹp.�,����d�2���Ĵ>�]�>�3}�0K��[��|�ֽ�
(��RNF�"�`�nf���!�i;���%X�=[�D871��r���U�u�i�%;G,
B
���T�\і�F��#Pf����ܤ�|��aX)��o�G��-x��ZQ�ZF��<퓜��H���ƹ߹HQ��dO��,0��r�����/ۦ5]����j�P�H���D�dPD�P�k��$*Z+������QE��2҅��i��Ɉ3�"���W�LV�ʽU�k[�K���+R˹��>�Jj8��䪴Y�^m��;ƿ�G(,{�|�P�+��4ߩ�c5�R��e��4�d�g��0�eo��}O��1Qs�M�t���g���lO*�"B:�8]_�c�����y�.��Za$`�ؔ��F�:Yl��Bv!A�f�Av{a&$?�!�����X���x��8�p+Y��D���l����]QҎ�~W����٦�l�D����C�
3D������oQrK��M�%�!��+.=�\�cHm�E XH�P��W���l2��*�΋�� �Z�y��,>�BA��� ��-.��@ ��3/���n�D� k���	�z��3��u���� BM*��4�,�;���|�ޫ�Y�J�<->���k����s�����sT���<�۴RP�M6�e�yL�p,��ŗ��
d�'�S(H��ޅg��7�4A�I�5��cR:�D3��q�<��<n���Geo��y���P�Hg[`{O����y���ƌ��\�v�liC(QB��
�K��URJ�p��+��w!F�]�ͩ��r�P��d�Ts^t�B�����յ�&���L��֌@�(u6ݢ��d8�i�G��+J��TH�~��$�O�����kC,D�C�g�g������L}�
�*�Mf{�4���GϺt��Al������墍��Eh?��bl	v~0+��@�-w�����I�`l!�)	O�_��"�G�z���ʴ�]�
�e(!��=۲[1_]�jՃ��N+��b���0�
��k�W�l׉��|���,8��l ��_�|8E*�_6w#���01�/�e���3��R�i��T��# c��E4���b��C��Q ����O��dQN��m�X��
���\��񷞟��㘢4��4�7�8��H��?'G���a�{�Rfc4$B�ӽ�����A(s;(�@�~Ғ�j5�2:�;�3ʸ'P�^�92Z"��H\K�ɯ��֜��QWŞ�������[�F����9K��]�x��з�4n��-��޴z�˥�[+��V�|�4<lq�F���R�(_�dR§oy���5��f�h��$FLZq
�\_�!E�S��\�eQ�P� "�7����s����Wv�E��*H
-��C-��8G-��ʨ~t	&L�{4�V[.P��JQ���A��8Tߞ�a��]_���S�t�WrZY�~L/ߌ��;�V������w�=<ƨ�N���D�U�E9[�U�&�a"qk^��S|���jd��yG�U>W(%��d��s(H���ݟ��7V-�#�u���C��l.WO�(��r��� �ܞza����q�:�5#B���J�V�!/���������?���役\�OI��t��9W�D�a5����d���'u�p�)�k�/��&]o/���i]�� 
�0�ͦ�C��7�Q:A�z��+p�8/<�CAҨ2���W��f!�rQ�Ҁ�e�|��b>�����ے7[r�^�!W���磰DI��ٺ�Ľ�K�QXa�.��lȭ=yr�m�j�w'��&�a]s��&{i��֤�E�Kˀ����#���i�@)a��� 7s�o��s��L- L隸��{�^��2��S���+K�K�3�U4����셜䒌Iy��Lz�X8���օ��iAqj���
=]GB4;D�t�O �e����C}G�䍕`h+I�ϯx�;9�����V�,�k]�{�vɑ�\����RP��#�sc���k6Λ� !������ڷd��#�Լ����sυ��S(H�����J}Ұ�YϺ��H��^��c��� ���K�}jl��kth�U{<_��Ap9�a�����,�� 3��<����睄K�O�"����$ ��$� �t�EZi�Ar��'�Z_��تv{b��h_ZR
Z?2�6��%e�}�a����~�
�p^�}wfx|	�2~d�=C	=����\�U�\q�u�ZХ�~~�ւ�8�s
Z�P=���g�3��ż���(E{b��{p������2G5�S�a���{s���?4ܣ���
����9��~�-�S����Nu*��ޛ���-���{ڀ�i����B P* ']|qK`�E�}m-��}��,�;ԭ�.�y��T����D��tc��D&ڐ2�G�܍
i ��Y(��5�'��M[s���ҍ��TV�א�e���� ��"�1��/*P��'�[��� ���.�`9���{BM^=��i�W�&D@�#���DI;���^qs�X+'ZA��m�x�?RF��6�a\{+�k6����e^��/hO�b��xWj��2�.'ѽ�T:�Q��g�#�N�{��-@���xҦ�ؓ��0L�_��i��˰�����P��<��	��Qq
)n�/0g�	��xn{�9D���M���	}f��_"g�C�H�I�r��؃�n��~c��[��Ͱ�FD[#�MC���N�Ԡ�Z_r][�Ӷr�쁰Kl��*bV	⟓�+�E=����4��!����w �p�Z�)��Yx��Y&��|Bi���M:3�H,a2���@�C��^U*��g�\�g���KM:6Ju�������)�tcC�����m�>q�w��L2�����`B����rG߂�I�Yp�=ݳG��ytd�T\a�����{l�����M5��gVW�E5��q�}�ԡ��C���(L�W�/T�+�5�z��)��/) ����T
�&�c��7 �'�_b�c��֪����K
Z�h�R�nw����G"���nR3h��.�Չ&I��o��ͩ~	+��E�+z�=l���%��F=�F3V��ɔ�[���@:vS�n�����U��R[h(����/8F�̐�� �Q�8����]��ھ����r�:dn~��-���xA�Qh����ݣ%�s�����o�E����R;&:��As��o��BW�i���cu�Z�#��ް2��L=�����%�y�z78p�<���i��W�7�������n>%��?�
�4���H�O?&�DqJ�g�(`crw�e�qA`�Ĥ�:�|m�3���v���<�����̙@���FU�3�HƯ�Q��&��
�k<rk�䈰֊ZK��`�{B��yÂ�1�������;M��¯����6���I<��އ� ����'t ���`�������w��sBc���4����j��/��ѿ0{�e/�T9���0>6��
�}�vS�ïM�����s��|#��B���C�i�u��|1�㼇�mԬsUu��$OiD/csp��)�4�M��S�T�-
��Ի�"�8��ղ~�=/r!�Ų(�C�w:��g���i ��\xv�5ƠA:��4�r���ި<����AϕW�.����t|�Б-��P�4,��T�p���G�mG�hL��YS�x�?wN���@�R��;���4Q)�
ׄ�.%a�5�4G���i��.�l����4^�u�D����&���DR�Zd\_kd��W
>=��016���{&�t���h�S���ʵ��@y���z,%bJ��a�M���~t��|�����o}�0*�`dK\��2LR�g>��Ę���.�4?��cU҃�y��pJ)G��y��|�p&��#�G�p�x����쬆Sr�3�9!�%9����GoX��(Ya	Ǣ��:KM���=��P�D⌤V�.��2�Qʖ&��7.!R˒�_~VCn�^҆Q�#�6�}j:���6V�r�x�*����̏D[{�G�P���$��mhaǵc+P�Y��@�E.�<!�y/�Q~��Br&<���bZ*��dy "�K��A���t]��􎈃�k]8=�_!�J��Q�q#S�Aܳ�?�k��jY|P�$�����l 6�����gFYf�+˖�h �G��pV��v�J�����M��[O� �Hd���.F|��t;+R(?��]��#�.5Z������pT�խ5���|=���ݨe*މ��e�yf�\A��փv<Yk�+9(�6�sӦ��]8(fR���+6zI���>3U_E�s-υ�8��y'��-����|�RAZ�Z2����W��l?)F�����K�5����d�Ĝ�:8g��&��@J�3�U}Ƿăxő�q�=H�������ù��)F��bɻ51��P�t��~�X��-�u�Rxjs�?�[���G��?A1a��`�������' ����ѭ�9O����Վ���ԾE��"���Ρ�{i����/4=����4
�7n/`s�:�y+?I�D���B@&݋7xf��1�6�)W
��۸�6Ov7�������l��6E���� ��[��qLF����-st�v1�V���}��s��V��R?�q�F�np�\�� 3�_���m�%|q�aY5������U�^�91~Yh*m4XH�hpē�GR�E�-�+��s�y	C(EzdG鴀4�̜�+1�*�T��{��M1�ك0ع�qi�.�}�IML,i���lRv2J�����J /�{p��a�
����<=堟;��r"�L�
�����.��ڪ�L�;# 7tx���ͫ�+��v���Z^B�:�ɪ)���$H�����q�f?�ÌH�rɒ�"���ଣ��y�����5_1p��i�=�Ӧ�U/q���/���C�B�]�n�?�_D!Z���T�=z��qE��~�
�V٫�N���w�K��%�A��<�(�|W��2s�т8Mh����g\0"H�ŵb�dPD�JV���׃���(H6�+CN�
I+ͅ�@������r{MJ�S[�V��ͨw�͹��~���Ko��.�2��<G�8��{��t�R����W���a���6R���r(���-����{Ay��kY���'W�JK5�o��~��y��(;/5�)�|I�ZE�3��N��'�!m�Y*�w�/Zb�;�2%�ͷ!���D��ЫΗ+�2�y�e��,��~���z[=z�Rk���p�I��
�/��d�GnW�o&9���x0��k��_�nN ���ң৹�]$�3�K3��@�7�1�x��|�*u��z&������ �!Ji􈮗�S���-������+��h܋@.݅<n���Ъ/,��`Ύ&�) ��j�Z/��ɷ�
'�-�ut��H�I$�j#���?��8~����W2^4[��"������H�$���� n;���W����)$`�1%5:�f1����v��P�d1'a]���`s�f��h./3A��w�v2��,C�J�~/��R�G1*�܌��3��<��ܓ|@_�aϘ":&�P��OS�ѥ����
5��@��M7����h���OTCMG{ubn�)+EG���9�0��2�}k�F���<N�*�����un� ��c Z_����n
�A�P��P}<��}�=�H����*��	���� ��(8yD�a�t��;_Ȁ�јԖ̙�L�3�r �����Xa�`;���y��-���&1�®Nb���T�����4�����o���$S��&LI;σS(Hτ�/�\�P��K2�<���Y��C|�sK���y�p�1-��o�v)E���!�J���J��K$x<��
�Oic~_=��F�����QO<-�KL���^�Z���m��(��_�/ȈS��Ip,���*HP��S�h5��0q)݅um�[�쐝���l�Z_a4G����U,���� ���E��D�&�o��cA�\:r�����=��lcm.}`�ۆ��n��b�)2tw�}*M
�r��V>�����i^��0� S�*�����&=��z ��[��w� �%Υ�Ɨ~��ũ�[���wi�~�p���Ǚ\�o"�U�'���!�����[�`�9��P��]��4?��01���W���A(�#��}j�	��^Q;%�4܈����]���V���G��A(�&Kxɽq�b�0�H�d	=u�n�I���Z�g�׼Vׅa�i-��d	��Vr.У<�x�q�%C�ݟ��i����O� �K�:����wq��t�i�@�}���s�E��vΠ$���Y��)I����`��NT�{A1���Y��F����8ƣ:�F���'�#���	t�LA����O~u	�H��Ԫ�>��G7�[)�4��n;���T��o4�pV������X�YST~_��AK��{"l\���B�FA:
NϷ/�H� N���DI��p4�1��Bl��O�ʥ(´ԥIȫB��
]+2�h5��lu��\�cRۏ���x�̠�*�Y�}�󲽊�"�wX��z���U5+�]6n��.��g��F�9�/�4�폕ۏ�)���g)�Fjl1��Q8Ԧ�zFXw� E��5��b���23	HY  .��|+FQ�����Ŋ�]&�^��C�ue�����BnJ�:����p��2T��o�}���B{�}Oh��O{`�(Ik����k�a��k�5	krٙ#T��{4�W5g�JEK��}��S^��W*K�: B�Ƿ�{�4��~����s�Wp��߻�Y[�l"��_L^r7d����@��XX�d�����%{=�LC�N���E��j.)�}>`p�ss����o�9�۽Wf.҄�evYY�%L�����
�p�+K{�x��d����(�"c�c��m����l��{N� �{ؚο�a����Z��=���m���Б��g�=������f���dU�l.i'����~�H���W	�R�Hԗ�sBk�9R#�F�g�MQh78�����+��R1�o�^����Q��\I�p��b��t�
�B��^��QI�>���y��y����&�'A�hI,�Q9A�Y!:7mIQ�,��kY��y�X��vRF�Z*Fk��vQi���鬜D@�1�ȻS�>~�M���+�U�O#�a�ˀ����6�x��B���\�J�
�j���rzρW,��|.�� �F��h�4����ʗ����:�k�ڌ�,.�~f�R��s��Y�=�p��Ie��ϫ e��O�f$��H��<�.��p�
s�9($N�/r�,�H�zB��Y�D���2[�^+��J�l%��z�V���Hh�J�d�2E�#$O�܅)F�2J+}����w��n1�#���6�e�bQadL�t��Y]�}+1E��9��P���  �?�~���A�]v#7N��\��{�e��su�d��眻�4�B����-f�A�`���K�����̼�	�4ݾ�c�?0� Pl�$�>��Kd�]kE�_F悸��\n��X.@�h-�1�����~�p��ò(������숭�*>�5�G���%X���i���釳*(�R�*v*�+V<���Ia~a7�I�n��7׎͠����1�ߍ�dw��\�av�/�>���H�F����X* ��{�6���QrkVCN==�tBt��;~�_y�6H�s�χ��V�ߗ-5��/R0�v������#N���WA�=���ÿ�C  >��L3s-���VK�=�=C�^�B�E[���%u�=
�FA�!'��R� ��GY�v)��jtmd�3��j�ҵ�Y!���������M�s1�7��ꄼ�q��h�_gi*�r�+l�j`���#�9���f$��WgV"BĶ4�V�j�|�%OB���@Cs����&?<{������0"���S_y)TT�[�Ke��-�t��Z�鄻�c��}NS�ܠ��`h���ǰ-	�
���|���ʤ/��҆J�� b����i�1��|�L<�}������>I+R\�:�����y̭�����ˈ�����H�Ĺ���b8���2&�f��mE�QtA�$��Gd+\��	��)��rN46Ϸ���`<��фw� �E��;�/H!�R��%Z�t� �R�_�ok2Hyhܥ{��a*b�0��슾kulm�_�~�����V4�1bW�]TY>o߇7�o���kO�w�ʚ�+��'Gя;� -Q�󴩰�v��o�4R6^a�H���X�u���i+����G@��ؘ)��M�c
|Q0 �k1ȅ���Jϒ � RL�̄�-}?� �A^�Z'���(�2h]�.Һ� ����[�$�K���$+f�1d���ۏ�VA�,�IM`����A��_�.�94�#F�2�!#r�bN��YLZ�,j�j��c)l�'4:'��Vw֔J�Y"��<ں�@f�2�"8�jur�(ղ��D�{-�U�9�QP�?Ŋ@!g2vt�?(��^4G��g�S�u�U��g���ϱ�ƙm�}}��\Z��Xt�d�O�N��|�l��\���B2_��NR��p`tO���~Z��-��[q���Dj�\ۄv�_:�11-��
������m1�o��4���T�]��a7ii�#���&�u��WR'#)I�
�\3�������[�n�0^�U��B�#D�G������AW�!w띪�uN��.dF`HM���`�����cr(�*ʤ~3R���el��y)Q�E6�Ƹ1�ʮS81��*��o�)#�ce{}��6�QWȖ��8F]�B>#�C|��V�w�=���<��U�9ߐk ��>�;�B)4���Y��ڊO�T���z�>ܨ=��R�mqJF!�+2�D����O�AnC�By]Zu��a���Dc��0���=C�>@�G��1d���F�~/����_�,�)=�_� �e��&����D"*�4C�n��6e�t.��S�;�P�uŧ�����V���G!W�dV�߳7�L���n��!0����a��"pE��J��6"U)I���
;И�Ѐ�/8x�OAֹpi��ܕ|G��+n��Y��h�*��wt�?'~���'.��p�-.4$�R���9����v���׏\<l?�����z��z�7���&TQ�L�r�q*ܡ�sr��]dpB�������'L�e4{ۇwn�ci[�AZ��H���A�re��i#��o4D�n��0�FwRύTYX�+�S=�o2z��tN/�L�|�ʹ�$�������0����\R��ּU{�b>z���>�����v�<HY�$�a�I��%P#9(RS��?�HJ����$�V�Zο��0K���W�.��A��GR�� ��&�U��d����֫ �Wf��(�uԲ�������V�:y��6�y;-A�PDQւP1N�&�o������b�om9�"��&���?)kK,{�=�kײ�Ds����R���=G1�ڄ�1a��6��GJ;��@�[o�s�A⬷�?���콉�庎 F(뾥���/��y����{y�R�I� P�Φ�J�[y$�;Al$�Q�Նq��ζ"t�W\ّ��M Z��B	��-B*V���K��)��)��"B}eeC>vV�k��,��mص���k�
��M#����q��s��m�J-T�,9��f���,_c������[%|��h�DW��򾭈�W��AK��jBU�Y�^#\�mV>؉G|���(�f��<�J�\!9�%T�<|`�sX5��ٹ"�a�u�|T�ժ���PJ�\�����/�miJҞ�`M����7�F#����x��V�Boϟ����۲��K����F���$�����o��ˇ�^��*�P#"�f8��n���W��Ŏ�7Կ{�vo=��ܱ��&Y9nf��rؕѷ �S����A�*�8�[521�n�S�!����e �F#Iq�0�/���k��
�-u�a������[߭���%Uf�K=@��NBHR����UÊGJP���y�0SR��m^,.���"W�"<�Ȭ�P\[��C���W�����W|0�d5q@k�ߺ���J�j�2�
�Q�,����d$[x� ��X�F��y�B�C<
I
�����"��:R��'���v�z,�n�A}w�U4q
���F�X�l=�4��r�6yT��rS}�.�k�e$Ɨ���
⯥���=%�˭���}�B�}��2<!��v �(����	?���{���TCMb��|�u6{�S�� ��@��=�;������j6KX[/Գ`Y�+B3[���_ OA?vMA�2ۄ�^ߖ���:�t���t�Ϛ� Q�- <��d���qd�p������dh�AE\�@d7ǘ�2A^�Jd'�k����=m{�x�A�=��$��埼��m2RH���;��u��=.��SG3wv��"N+9�*7l�`;{jJ��W��P�rU��*pa�@?�:=�O񄇢���D�=)�U��d������3��/� ���01i9�1$g���R�ÿ���W��#$#/v�I����%���
����x����$F��ʨ]+�lt�LH�:�d�PbU��<G�j"��/����U���q��s�З��|��-��M��\Ŗ���Z�O3V�XoŦ����K��Jǉ޶������ќ�Z��->�I��Z� �^�tΨ����|p�j�~�|�R֢ �̺��P(*�b[�K�:�Џ�����x%����>�6:���M�ߛ9�Uqٔq����G��x�H�>>Ɨ`�t�%�s?0��+hwB�n�9�{4`��@���￠l��/� u�-�B�&3���`�O�����hvJ}��c�j���m��j��_�� ��/�$e��|�hE>��\�&b����
�r�몒�ҧ�pٺ��^H0]w�2���������T�T��92;��5*�lD/�P�^�Ψ@[\Ɍ<v� �<�M%�	�?��n;9�r|M(�<��JL�� p�~[zE%�Ƈ��I����4�X�$wӉ���E�R��V���Y�FO��v{�369{^����N�\t��7�n(��}���W�X����A+ם�X���Q�W*w��݀V�k��/M)�ND�y�-Y#/C��y%~���R(��e��h�Z(Ӵhʪ�x�ݢ睵��-mA��/Z悮R��r�F���ſD����z��=�5�$#*�3A�c."s&%bK�;����6L�5�˃0`g���BL���g� '����y�&޷^������V�`S=�Y��rjŎ�4`��^��G�nW�Y  ��IDATsP!r�����2��a�#�9C��bYZ����?���$-�iyZ��E��d����h�yW�U���I�^�|n+A>����Y��-��h�6LY�q�}1+d�ݬ�A��97�C��5�G��ʃ�[,9�}֮)+eP��^c[j���۷���RX��]�W��U���7�O{k@X�+T��5���\WN�w�Fq$(!��n��[G�Ϻ�1�XH�1�h�1�k]Q$UB��W��� ��N��0�:;���U���8(������AvFa�1�|�\�]�Y���R��6�������3�(g��/T��:���=pޠ$�~ZWaH
>��_E����W��x�#����|��)����|��||Q���ǯEE|�WG�V�(��'}Ba>�������͉�&���u����5�о��8�+U�s�0K�+����	Ώ+�A�����Za%������B��mYo=�ǭ������d7Y�����G�U��E��&g�����P&����|룛���Ǐ��oI?��g������^���憏m\�Vo��CsHP+�+�)%�KI����:I�i���VKj���^�aح�4#��KVh6����~����3���߿�:��@ј�:R!�3{s�Q�`����;E�CS�m*~��bõ���}wxW,����V�WA�W����s�ˤw�0R�1�V��k��Ĕb�Be�O�����n�����e��\�Pޥ�/�9�g�{å7��Gՠ
~uW�c�	�5�%�P��ҝ;Ŭ��_MR0�M����"��˥��~%���4��{�/_�ߴ��*�*6���i[=Z�ǿ���#��76���n�7a�6i����e�'̮���������}s������]�qCmyr�݄����Q��M��	a��	]�>P�5����Q3L�`mi��v[	���3�_!���/i���ݔ��&�J�������:6�+#�J�8��߶���24U4&Iݫ�V���U���P���MX�4���ۗ�ߔ�:�?�X�(���/#[����ߪ4�/ى�?�%����5}���,X5[@)r�
�	�LW}���>"/��s�� �}{^Ȩ�ۢ��H��Ť�'�Jٜ����O�S����ˏ���v,8=�����z���:��M�v���{Dr�w�|���K+H<���i���{u�'�_@
8�pf����ȱ1ܛP���&��\�9���Y�7�/�he��c{��4V}:ϳBt'P��;kKٮ�2���>ѿt>k��~`i��m����(�d�/	��(����Z1�
���W�-,�z��X�����ǿ�-}�?o8���>e�
Њ��a��g�&�ƣs���Z�+<�u����Ú��g$+K�'P�"歭Y/����ͫ��f�H�Gk^�4o5֢�����.���K�?��-k��������R����/e��!�2\��W�h�W\R�{<���m��Y�.�ո�&l�Pe���Xu��hB:�)���1q�_����/�iTa<�x�,�9�}5��{�k�}O��4u��q�y���~�K(HV���+ �L��J�%����. �`!{NN&���B�[���c[9�Q/�@ޏ�.���� }6� �ަ�%��޷�,m���J�]j}��U���������D��(�S?�o��d1�n��'٠�G�h�ᖈ`Z$Q�G> �Y�ܶ������*�*�Y-�k�U��
���&�P6���� E؄g���qAl@t	T)U����-cKv���5�g��d'cM��i�p�(Gݘ� r�pgi5[Z�Ǚ��b��V���_�~@��2Xˊ	�[�-�N!��.m%ڭ@! �^����]wD8շ���+�����B+��@m��Y�z+Y^e��,�3~��Mn�+�c%m /�k~�5�@iR<�ТX��n$��j%k�$_�����o�<cB�x�fN�v��_.� ��ݍ��WQ��5��u���=����v��zĲX�c��[Z��t�M��w��oSA� �jX�@L���T�.��T=�8�b�y�BP?�znm^�r�m����]Ekr�-�g++� ���4�+�����xW�~"
���+ڬ���C't���5�g\Rr�\�V��~d��x��l�A��#!W+�E�����e������K1d��5�۸j�2P��V|;�g84��W������,Fܣo����أ�:�E��
N�lɠ�!)�I�}�X�w��MC��O���^exg���J�l�ؗ;JK��2�h���:�y��3}f/17=�V�I�ڢ�tJ�V��֞�4��۬l<���˴���;�<9	v�����*�����QP�]TԽ��d�R���zH)�~hn����+0�<,6�,t��GRK/�����PJ� c=�'+ɷ(��J��A5���n��S�g6��
�Ϫ�Y���R۫ϫ@)�B�����zU>%w��b%�]EY���jH[�JA���:4|Ъ(��G��y8N��n٩��6���i�)3-y�q���뻧�ᮄs�Jܼ5���eg�2�`e�j*wcj%:+����4�5,��`cZ,�~]C�ƙ� Y]څ���G���?��$��p��M��!�=��d%N��f�'_��޷'4�I��S�6 {�*$�߃#����'��O��1�U��M�_ N@��Ȉxʑr]��2]��%�/�����NǱf���^�#z~1�ޏ�H��~��$�/�M#��z%d�Lb)��^�Sv����
�KM�"�H�/���b*^,��`�i��\�7f��-�*s��uui�{[,G4=$ɸ_���"ׯ0��	�Q(?˦�(.">�Re@w��/��J� 	A�����JW�T�^���Ɠ�_��sD@�k�m�l�n�,N�=����:w�xd��"��!�$x�%ZI�s��^��1�C<1�G�B?�&~���mML�XF��˖�?+�K�^<T+S��cR���u`t��7ݡy��4s���!��Tn�⭞k�?oUYɲh��{�j����\RA��o�� ]N�Xۑ�Y�QF�En�Wd�sI���l�6a���g.�3h־�1��X��P��[��׺t[	b��n�|'��Y�	�����	F�q��J{5�4RP-�eP3�?tQ�8�$��;l F@��E�l>R�j��V11m�~�)��,N8O/�B�V�HE��F7���X�8Vçn!��!��B��]�QSZ)>���W��[Az�0F�&Q��5u��w�ox-<R�z���ݴ�,��L��	��5����c1�E�K��]7�S���Go�`�z��lυ"(:�V��v��^��E�G�EK-t�����֋���!�c3=�W�:�uN�˷���^΁a��C�L<��T�R})�_ĶZ)&�)e
����̠mc�V`�҉��#]���&|��=�Km�Kh������i)�Y�[5����ޡ3��O�`E|�?��ǖ�s(7�N��Z�Z}NC�:Π)��b�/� Y+�gWU�	j��Ni��/291�(x|�<u�`�ؠB�p�������?���AI�c��V	:zA��]��br��X�����)Eɭ�\Z�pU㊬�~Q3��^kgu�(�N���&�
��+�~��ːF�� ��hE�ս7��Q�i5USw��r'9}�hB�e��y�4�N�����ı���uGwLn|OY�c����Et'�c�,bq�W��Ƥ+���}9�[��5#�6z<
���
���ͫ��Y]_A:���|�����w�:�5��a�)��	��u�Si��Կ�J�+��Tc�ԇ]������:Gu=��q	Ș�����wQ�(�����?Aq���ώ��w����ӥFcJ����L�sê��v�D�>9��Z������)�F�=\%Rj�_[��l}����	N��A�n)G3J���W!�%���t�3mtQ�Q����^U�'�2���?��U��
}�0�	�������W�������L�u��w�{F�1kcj�����^�=C�]@z3�2�$�BO(r�p�]��*ꘃK3�A����>��) k&}>�M���@g,��D#�]�+�E+���y@|+��䫀�����W�W*�A�
��#����ѱ�T�����=�(�R�vo�;+N��v�#�#,���P� U�v��l8`7~uqn����z��ߓ5<���\PA�>��w�n����F"D�(jhN�5���į���N��Ȼ
F"����V�����AC�v�܄QLi��}����Hk��a�)IHkq$�(���<���F'��6xTD�!;i���sy�j,W`�q�;�l8ԉ�.�����F��\�Z~������LĂm�S:/��\�a�C�}�ݛ�K(K*oM�f�է�����Q'����O��30hp�>z]2V���
���P|��dX�kp��9)�n��@�;�Zc-�D����Pُ���N�:�)w#ό��O��&1�J��V�=NVZ�ls{�n�ڮGn�lF�̎ˣ=i�ÔԊC��"N<�k�<�%Uvя}��s�Z���>��s�L�S���0��S���b��$N����f��O��Nk/6��Ėڸ`E��Z��݊�eX�����[\�@ծ��l�\��2)<H�>���'I�E�v��m�����{ ��� �s+CU'a148�lX�7膽��3�dm2Ro�� u����D�Q=��r�\9�µ�����|��W�J'M�n �?����.�_��4��y]e[v1;Z�}�S`�vI�ky�L�*�Vr>^7�v���n�k@j�u}G�.��w��4��i��?�o�W�*�lP|?����S�f`�Y}�X��)�rQ�B��ǚ&-���@֏��3 �#�I�7d�K�-�����@^�mͩ&.p���%_ �2���Iaܻ�J�/��&9����;x���>�o���ƹ �6�>Mw�^],��E�\�J�N�.?�a}�rn��}��:�Vݵ��v�;\�F�����O9��)W1��C����s�(@
d�:���J����5�9[�(&�UQ��WQ:�Z]�-�@���$�p�4�)*��մ��� w�I��hO����,�����kMB�p���+F#bw��d�~�t����iueP%�LimL�
�p��j*]�3������R�k��Ȉ�@V7Q7��Tm��Uy�<��S��1�x^?�d*�^`�&6�ЪI���8��#�B�B�J$�7QfapȯR���!�(S�?Eգ��:m���.�0�G�b�:�#��p3!��^�m����	vS���-��-�p��T���y\h���DV�Ҕ���I4��)��w���{�mh&<�c>T*��2����^]���	�U�c[$�|�0��.���DƑ�_A��R]!���o� �����*�C
qy�*�a�g��8xd
=e���
�9��THHrk�=��~ǀθ3p�}~gAwc����a���j�*z3[?<f��n?�(��&�џle�UپL��K��y��;C���iN�_n�)�ĸ�M�CʐI>���׏��Ya��Z7���PJݼ7�â��)3�OӁ3v�T+.�宩�#������*�;V�C}C�++G��	Z�U��y9�:+Zb\�!�
`��H���a���'�r
R&� v��x���PwޭpHq�&1�� ��yd�!�|��sI�s�YB��`���v��=G�R�ЋN�z�������O�؅[�m�Mz*���L̉�Í5��d�����P�i۹9�j����J��K<|��.�T��r�x�{��8�����쎺���jV@z�]�3c�uE�A`i(�@|���H0Vr��S�-JU��:3]9��-ܿ�rD�"��_���3�ߩ_^PA*�iC�Oq6H�Y����{�pQw�����l�3����7�<�ݝ�P8&?�DKf@��Y3��ɳN���̄�߳�x�9�JMi�=bJj�|�������R~��-S�̛Ή���L!d��a�Q��;���^�0%�?�VgB[� �CFBeS�(O��)�Atq�Lᔟ�DV�uu�d	2��e	<U��7 a]ϯr,����R�$��:Fu�`?Ms��0�(�K3��6��K�p��-U���ڕ9Z�?�j�wDY|KMං�K}kU�۠Z�I��7J%r��;�2�̓�B�r���Xo�9oo��C����LP�ʱ�q�yE�8R_��Yy��Ӎ3�߷����㷀�K*H�B.����g���ʂ�O�`X�Q�A�U�o���8���X�T���-ɸJe⅚��j���$�̬�j����)
�n۝��p�����Kٟ�$T�����]}� ,��LC`e�� X�WJ=��W���k;�5��V���};xG'	�����[�D��&�E������H~G�����v��c��v"
~S����N(��7���F�
;���iH�_��1�|T�wd�n�*w�R�G�(3 �G�`�^0?^�vuII�$u�n=>I^���G.�y��6��"��|�P"%�M�x���*L-O֓�Y�u��L��Q�p��%�SR�K��av�>�v��Å�� }��ǧ
v_�:��G���C7��0��%f���6 �(ߏ�Y�e��pY��F
fn��J��oD=\�����aNw�#uJ��(y )Q��ty��v�@h0��mO��^++5�GQ�#���k:&� .� i���p���x����>�@�\����a�ﲵ~�� ��>����Y�|Qro����7qx:������:��}��-�4922��`�����|i���W"<46&�[h8�H����7�ɚ��9�~��21Ƿ�|x<�{+�.����i��b���/��һڞ9��]c�k�
�pa^}���Pa^[{Р�Qd���{�F+�:!h�Lyg�4b=*��W<���:*T��m��[����+0G�8�ҺW��M���J`=+��2ե���<�,a~%��}�����D�������c�rNh�zow�,K���Έ�^)(���KO��?o7��l��y�<$f����]��0��t}Уp��`J��~|����\RA�>����R"6���
9H7Lc��t�����
����+M���c�]�Ԭ�����|_��w��@��,�o&�#16h�������`�X�Qق �`ܙ��e� ��{j��`�Y��Voi�����x��![�� -=�-��[Y�w���@���D�O(�D[Ϝ�2�n��&���Q��O�85�r��W�X�*dݬ�k������. ��;u�O ÞC��s���T>A�\,��}��Z@�B��ֶhe/?�����K�[���U9�<���
�>*1�wkv�b��u:�+������0���X��I��-xG��
vF�)��t��(��w���xM���g �����,����f�Cb6�i:���pW������9��T���Be��'C	�%�"��w�ڌbv�< ~���g���P��d�'�]yMI�'��V"Z���gm���XJ#g��`�o{F�ਏt�X����/��h�O����O�H����o�iI|e�uE��=��1�\�{8���
}��9<�>ڙ@E�_ ��j�^P�Ŷ�6�w�����$[M���&�����qL�:st �g�J ��IH�ƥц�#+w��*H��>�O��%�ԃ�Y����L��Cw{�^Z�G�x��r`��gΎ���_7W]oc��p )��h����wMa��-�~c�aWF��]�I���%�0�!#��
�	�ޞG��׺�g��Mr�,�O����/��SZ���k�7&<��.� ���^�e)J�s�ov��!���o���Q.j�z�B����7��#�f�خ�ʕ�}7\zvJLH첫��_�d�a�hi��*i'w0`��u iؐ�����d����G��Y������5.)Oͨ.m�����#D���bh5>v)�����qlCf�$NT;<ЏɀtE���2��j������!o��2��3�N��l!L߸3�[e���N��o��� � ���3��[!O�$6������w<�Z�_��E
� au>&�5GJRS���!	���o�ܣ�4�(%�xt�>6�P�dh=�ٙ�a��?;^�rx��̨������� ��X���U9��$$k���*�͝]y�K��k�g���t��o�0_H������0�2_�R��r����l�me%���ϊ�G܃�,�e%��	̏�Br��	�������R�4X�P����X~�ǁ������z��5T%_1��l��ߗ8�%es�8��o�(�oJZs�Sۻ~~=8NA@h�Ia�g���W������yR;ʺd��Nd^�YZ1*T�������1ϰ&����s�p�'��P����|�Y�1���+��0Zz�)[���7�턻�ܠ/h�^?1�C{-<R�#uJ#Ԅ�0�UN(�Ic�Z���]d44.����	�)�E��̋ո�(J#m #�ZA�6#����]..��:�(���Ŗ�*�eAA�w��S���b��t����	�(/����h�߫G�p�%��bR�գ�:dz'{����W�穋0U�ȗ�paP�� 	d�s��a�}#-�
�{�*|	В�08%���n�u՟X�ǻ�>�@���&��5Ḷ�⽭(U[�0��@`/�����*ִ�zUtL�Jgo���%���g�<{������@0��P�^OA��w\}v��f���� le�K]�q��߅J҅���vi4��R؂_
��E����-�阹�Fy�t��}/ �$~�V0�:/��|�g�#�ps_ʸ���w�%#;�Ԭ��N��)���N�����U���D�*�mx,��s$��7)�����c�ڴ4�P����'�ʈ�����o�!�L�H��ׯ���m,�����UR�[�I�m�$J��޽�tY���;k��Kp��"�2ʛ|���0����	�=���X��J$��]U;�����	.�.=�q%�%���p�7kro�����V�
�7�+m^���������o+-�B�2V/��>z�/z�OtY�A���,h��x�C�!�Z�(2�V�<�M"�ZjK��Ot2�U�@��Y��j4c����L�)@*�0*[��+�\�A��YBNH��"L	~?
)��� ���{����H����;��Bo^OA"bS��X�9��H����� ��RS�S�1.'~�b;_~(H�wmЋ��9���@�����<A4���\�����.Lw$�#��������#�w"�,�����pk$v+5cE�Ke�-�<DJ�RP�AfKs}O�&��ʬ&�n�e�!���5�ʑ��� �N=���kK�S�2��~(�������|�(ג�{pVq�g���Z<
��d"�挭����/� ���k
���W���Am1yJ��F�#�����
x){w�����Ж�ԾuZ�$:�K�#f`�Y�j�t��m����T�c8W"�=h}�_�׽h�ɢD�=�|/iG������:ɭ�uZ3oN���!ၤ�)���Ld ]Z2-�cY�ږe���^����-�|^kݱx�l��r���j�}�1�^�xmۋ-�9��IW�����NA %x W6�1���
3������c�v�Ft'�;K[xU���kzd\pn5p�g���#H\B���T������3�V���L���9�V���MT�fܘ�<��&�SW���Y\�n�{�ajH6�����o�[��nůAwP�E�Cñ���$��NfA�t��@�ܧ�"0�c[Z�֘9��/<`/����,AW�$��s�%<Tg��].J��N�*G^��ⳇ�)��D� c�a�ю��ݫ���@3��V�!eL�N������ȩ}?�y�m�#����p���Τ�������;���X����,�5Ѭ)K����2�[�!��o%�i�]�˶@W�V��&��;Oq:�3�ݓ�-'���� \NA"<f����@�t��s��.���}2�hrhi���y��J�+w�C"wڥ=�q�wa8�s徬ͱ��Þr������U1�=_�T�s�~<�ʵw�٣�֣�8���U����xە"-��$[C�
ņ��k�e:�x'�F�HRu
��U%a|�0�r0_S��K����5�%=L�y \NA"��0N\ğ*�P|�.�wx� �� ���o�N�&Z)ĄכkZ{�R�Ҍ�t�9�d�1��e���P���"�f�D=�f���J���ߊ�{3�{�H=���%��k ��#�g��!9�xn��j��W��J�Ұk�ƞ����b̶�݅˸���I���bR.D��T����U�S��Ä�����*H.��#�\�y�O����dxl��;$D�mK����ƾ��^I�!�χR&#\t�Y��l��Us��k����MU���t��	V��=Y4@������] �����+���!�"5H)N�'c���P�":�,��5ɝ��Քo\{~/��WW>e0n˚��iYᑶ���y����X�?�4�|���䣽��>�d_J�t>�7�Z��o{�h/N{?�����H��C���o�������+�� ��Wb�0��>X3���|u2��JC����Ԧ%�ؑ��K������3��hT�]4%j���}ë@�
^F�p=��ө9G���e�:��zQUX����z�EZ�G..��6����e�喝���RT�]jש�5�fD������lڮ�9��H�m����V�b]s~���r��
��0���Ey��Gh ��M+׿�X·%��g�>	z�&]��H-I9�m�6L-Q���;p.v�tz�;��,AIy�dκ�Uu���mݲۺ�]�ܼ�9up�q;21wV��|�Ҡ�:��Uj�ׇ����d8u�X��E�B ��������\�����V�!8^9ߋ�g��܃Q=�DЧ������Dy��v9�dA��[+'��ځr��.�-0۹�m|����d�"��Y���g�= �t�4��x�HT5������B�I���7g;zp/��!�����-�=&�}j>\��_SA��Ȕ]E��y��/������<���.��.,M��.
�ݑCc؃���_`*
�����K��4���R�f��3+�3�e����_q�"61���Vq��8�MN�_�w�����r�-�D�����I*��!��<��б��2��lź���VAII��:A�9�g���lh_Ѻ�� �;"�hn�~D��9��t�]Ɩ.q�U���3�m/��yk_0�?��P�}��?���dCz��^(��2Z��ִ���tW�1���1	�)�sdH_��?vX��p�ʠl,S :�}ζ�� טoYc1*�^:�q�*�H�D�@pE�4҈��v��w]6{����P*�q��
z������-T�RhXx�@�ë�
Rs=yHIB#P=f2�� t�u���Z��_I�d˧-�HA���}q�Z�+�)��=x��nƚ��r�0����)G�^(_V��ߞЫ#G�����z����O��fw��C�d��1p߳���i��(�z!�^��3l��1�9�������?S��{ٙ��-��m��V��۶I�I��(���ڑE��Dq�<���xKCЇ:��\���6V��;���$�J�s,�Y��G@zv*K��`�jN?V�(�P	Q���g�==�;�%L����_�N.����c����7�X\�l������Hس���oz!�i���r�	-�:�ڥ��h	+�>�}�[A��RS�H�;5�@�ձ�E�81���ߜq��L�@�Q���%%����"ȝ"����s��5;d�@Yuڑ����>^�DH���}��C*� D���{��1��-�膬���ekXw|P}��@o �JN~��yin�x}Ok��l�,�V��.����< W�^9�ghP�zJ�#B1	�9�_�?���k5�U��2�-�R�$Y:N����z
�;�ę�kd��eׯʘ��ï�x�����΍�=��4T)>��__΃�͞ȫGmN(vi�KM�ϧ	(�9�zoDig*=Ů�X���ǿ"&��$Փv�U�ӕ��$.��shx�T�{J/��ݺ��<\�"�HG`�Ǧr{�I�ۓ���ઽ�Y#�����#F��h�Mm�K%0�.� ����`���o��=��`�N��������1���I(�g�5ge`X���h��c�[� �?`��W���"��}�pr��� o�滰m���}��l��UQ��la�.�N���=\����Amdp/�Է���r���K�ɝ�&JO�Q��(4�@���&��:�h�b��7�8��c*��3iğ�y7���=u��ml���o5�>��=/������ԍF��qJ<6� ���5q�=U��xB��Ů�l�HQ�M9�D��7�09L<� 8��N��ǀ�̃K��(��҄���n�vvq���W�n���Tv�]\�)r�xD��Y���r�׎F���N����qI�e!���������v)�UY{����\=�䞶��"��ţ����,�3N����#z�����ᚂ��1rJ(?�[/L,/� 5(�HC~ r�\��=[����us�|��v=pb��-vQ}L;�[�f���W�V���[�V;U���|Si&Q��Â:�((Yt}�^�q�'��8�ab����b���3����K�_ۀM�;�(gS�]<�Kls��r�\�iN^�^�x���^�/��x�O�V�E\�:S�4/����zgArZy��&/��6@�ޭM𦌞�y��P��WI��s�M�F���מ�c@�W�d2��n�jW�޽k��
R��>��8+�3�lЍ��ϳ�sBTd��-�r���&j�eT��,��xg�9�j��g�z�XAۿ��a�\fp�#^�0��"�i�X*j�u���c�}e��֩*O}��,e�����s8{/���6�nw�?���:3�Ǡ�5+ƪ��5�M0	�{\�+	f8�x��sܾ��Ǡ�d���qM�e�4����������<�̶���9b�ސ�	g�GeQ^�.$^9�V�����,ߞ+��l��~�uXy�`�~��]���$aݣ%�-
@�h�Od$���2��P@�����ʑ��|�Z�!^��=}��"P���P��嶝C���Mg�Q�E��BJ����b#� ���FE.A~Qa2���r\v�Jm_QP]	���!�dV���>�[YO��6(�%��3U�#�H/��t����1J\�*���&2�\��
�@+�Ra���d�휊Kk���mj6����潂�1�ψ�x�*���Nϫ������x��g�HT����h��Y�qR������A-��w��᠂Z{��|�76��^�Sv����=���PXf۩q����8:��ײ�V��A�]�F�}�$rT�
������!�Oo�FE��l8�V=��w`x�'��f�4���(y�=��9��ɰ��V�M���Vx_���ڽ�%E�#����"����5N���e����(0?Ɲ�p�{��Ӝ!��6IX7�a�~tt�z�k�ُ� YΕ�%�e;y�@0o���x$Eq�$��S�����f7��U��@�XO�7I œgҪ�'S6G�<������^����/�R+8)Y���|�d�|�����=����
ĭ0��2�nZ7�֢b*H��L�s����-+������+����V�U���/%�V���b`pi�h��	z�%�ͩ��/	�V�+1���i���"�5�"��p[��k�ѡh[��]�sC���y[�䊖{7�$���(d�����;E���R<�ǟw���*��X4\HWd��*H0�b�7F� �*W!/L��{`x@��#B� ���� x����6����X"�{
j$	=E�p:�%�ʌȩ9�F���ZZ��w��CXO�ĩ(q�x�6R�S5��1\ ѐy��d�In����w���bw��x�ޡ�%hqfk7��.��e��$���o�a����x�
�+��ؠpJ�������?/��*�|	�uAo������iyK���d�1���ʷH�Y��lNDNO^k@Է��P]���6Y��~���
s��	p�Ph�U��=��R��$7�;�����ǁ��$q�g��Q�L�(���/� 5`K�
���1�h���
�P�RJ�i��˅�
� d�Y��\��>�&��'�e'�E���q���T��$���ě�{P�,uG(�3Ì
N�Iܷ�E�7pDV��H��vL���c�=GϹ�zOa>��C��!4aeD���%�
�a�e��J��V��q�Z��+|GE�B��p1!�S�X_0:~W�al@��6!Ȱ�n+���:�И��{��z����-Ч��%��W����W�b:"�r�v�+�2"s� ���*]&dw%�:�Ӭy�b��.9@_3`����T<N?R>�"�9��>j���?�4^<F_��ٗV�vaG�{V9`^2%}>�a��z�^���?*b��>O��;0�5�� ��ݐ�����>o5�x��1�%jھ^�A�����xVp���Q�nXHrBz��SU�6�5	��4� * ݃�ߗ�S�olx����X�t���qxa�2�qQk���n��:5a|t�*���pˌ
���2V=��| �GO���;z��bʽpQIX12�[��-����b�eV	G���X�^]xUs:�����˴\�'؅h���;0�8�8s�AP��4[Ѻ*U�{�D��),�H��~�W�X�`���ꮪ���Վ�0���B#�RǌU�	��<��X��BwX��G��ytq���̢����^�����7s{��T>AX8	�S�@Y�=�o�$��d��L#�S<�*�P��G�C[�E���z�*D��D���zPB\�V׵=O���2�g��:�Cۢ�X�h47;�@������4h��#?&���*�o���N�<	4m̨5�TV�)rE�����涡G.ivA���������+"zX=����X^*[�Z����^��
����T?Ѥԁ��ܧz��l������	�jOx�l��O�Y����oBXH_'q����	�8��`�>�q���q�`a�:�U���s��\Kk_~XӬ�^<��ц�o�E�%�F�~k]�e��ASF�|z�ƩyU�9���/UT�Hc���`�l�4����J�ì�	��<�?\!��Ϯ�t����6�uҁ�w����m������=$���ǥ�y+���n߹�~_��[�{T�6Sf�+	�0�r���^��k��
��c�\��*cq��^pB@!�i���s��\1
�/giD��������zt�~�jd��OA��#���@σӀ�{�c����:�1{�K*Pi���E�=d���=�wp����O;�V�B�)����d�.`N's7�P`U�x�x4�N���f�˕�U�ik
MD9���ފ��:�v �
��sL��8G�l"p��*�u�Y�∉��Os��=@ـ�TɃgpc��� ��K��^)�髢��:�-���,������p|��#�ݎ} �9q��ߋ���멠i<�t��U>ܥǌ
��L�5=4�r��im��-�[�3!|\RA�gO�(��.v��9+�<��{�mŎk���֍���啄0+7__N3*��ɩ$&ɏ�gĝ��Ŭ�@"6��,C�����Mv������)��$G�R�G^��H����
��IM� =L��8��/'H$��q�u�ʢF3ފ�}<>|N��s�
�Og;±Q���6e�K?�o~�|���|2�ޝ*��U91#�*�nz��3�[�T�8a�U%��z��y��~K� l4�X_@�L�����9䎘�?	����>����v��3\RA:$�=j����k�捒��hj�y�����|weC�_Q�}V�N�����M.���\�����@�����r��K
}�PGW��#�ˣ?�J���6%鬴,���#pMq������^y��nF����*� +x��V\����5�)���ڕ���й�G[��H����`\xX��ڛb2�����.�\Opq��:	�5�1�L�"�"�$������o��'�� R�i�A8��O����(�����w�[�zZ2!��e��z�Y�T��mÃ�f�#cG��o6��
��#�B�r���X.����E�0��7��mi�<޼����6F�9��P� f�V.���X6����l��j�[�跹(|��fPrdq�����ҍY���L�&�� ��}��WZ�$�Z)�7��<�3��9ʳ�k�ݍa��
JI��i��3�[�(wk��l8�T>����R�B9W�@)=L�I���5�8�4*y
�.E�9E�k��M2���p徛�C��2}�����L5F�S_�1�H�ް��[V{�A���+����ȢQ��WL~�+�bW�������-pM�8O�{[?�]��F,v��?��`�?�Y�^�q~�	������d3A���ɏdЦ��U�H�YӜ�C�q^
�f�X�i�:��!��50ٵ�q}����K Yyu}�ez3���.�}1K Y&���31>D�`�iմN?G��3B�{\�8��$8�kV�ųc��Z��0�<���o�����iM\���2:[�*e�(A���\��TX�M�(���Z���p�	F'�e��%�d4%x���C��)��ؽ�X�OwB㌄�ڦ�b%x��}M��I�9! �	���Jy�� ����u��ǩ .�H����$���xV���{�t1���m�����J�Yʜv���5��t�U%���7����ΗT�8�����)�"�͢��KcC_Z:5�N���@�{<i�'�(�]��#��.
�U9ef�mp���])��p'N��Fj�/ox���Š��o�jtX�240T:-�p-�� �qB�ӌAf#�u�
R��/,�"-[O]#���J���ʎ)�S�Z�h6������N��������J�ϛ:�n����������v1�x�4N���H.	ܠOSO�t�^�Y�$z�]r5���_<��]�G������LK�:�A_t��/��~l���[��B>wK�����
מLؾ�b�K%y��x�Q`��w�7{j�9P�.�S��&�G�5$$6�����H� �X<�М����x �m�[��M �UX�C�U&��{�c��d	B# R�}���
���s��3,�2d�X�e��K�7���+�� �6 ��#!�i�ϭ]�dI��$�v̌1(�C��e~��+m���bs�JyMC�?v�$o�t�s��M�|"�`�S�Lr���ҭ��)Xa!����4;��}�M��EH]��y9�x(Wb�]FB=I��'|�]� a�u�.���AU��;�Y�Z�ѝ����KP~��̏���5�j��QT��)r�%�o�3���;�G�"
v�L���pII�T��%�(?i�I���0�I
��q�7U�}5�.��y\x�@�E?�	�m��)�%a�"��(N����T6�V0 '���� &���Ê�T��y�j��r��8*4E�=#̰�]�a�}��3�k�*<h ��4�9eR��*l�'0���۰##IR��Ƙ 2tF�c�]�9Ϋ%�ꝑ7:|�9�Zݫ����o�mW7�����b���z�tx�^��Xu�N8p�$z�����W/���>u��C<W�$�y�U�d��Rz]��
RCj0��m �=IZ+��~E�u�8bHG๨�PM1Y�w���MV֒�����<p=q�������ZM��~C��L*F�!oC�זA2v�s�N3�H5&Av��_؛���^�
�q���e�mà묾��S�틕��`{���_�I�S
��=r�����#E0i^4�s9XA�zwǴ��[7��m�I�ֲ�Ɍf�"Ep%������ [�J�G|>�8�#O�,?��6hË^v&OoŲ�.:����J׽=[2�A��]�~�Kˑ~Y���膙�Ȯ 35T��E8R���'�cX-O�<�u9�x�"	�D�d'���O�� @r�¬B⛎�70�9���=X8@w���F�G��I�8R�W[�9|�w��P�9�c�~�&�#�cY��aq����L�S�� ���0�)�3�d�p;uX��֥��:�|V�	��a�}k��^� ��n)jt,����t��ZMe��Q׏ae*���@��c:5�΄�]R"!�)�+���k��ø���S���z�*� � �0��X��+��D"V�����FD�8� ��.X-R���y㳗�r�J$b[�ה�e�}�������G�сJ�Ŋ�|��kS���/��.� e����	#H���?;T�&�����D[�(<P����x���#7��MD<W��b&>�ϼ�W0��g�@X(U14����Ԅ�@([雱�d�{}^�1!d�,�{|��k��M��nYs0y�~�w�=�>*˸ۿ\�>�7I˼��QHߒU���JŠ^���|��U���n}#��N]����/u��䲤}le`�eu4��~"��}�Dq$OP(c�ah�T��QZ(�	�r��UsA�����bզd�}�����,�_5���`>p�W�ࡤ�PW���ќ��,˒ֵ]�L��e˼:K��K�7�L�N���j�!H��?y�r�!#X����쐎<��e~L�F�E*��9�7�[���^��xx��c"r�g�)��)lm�XZV �z�]���K���]�E�;�fjS ؽ�{�����x�?�r�bj���e��y��؀����)H4��_C���»��fp�d�;���� ��~jL
�P;��1��!������4C���Q���db����/u��f���W�<�0���5����Yq��l,{xEbĭo�	�C%�Q}�ey���<~;u��'N��H���RPwxq�)9�e��؉��U�Ⱥ��I`q�,P-�> -`�8a{��8��9=vQ�]!��-20=!��TbO@A'T�������$�ҙ�Q��z�p�m� �9��D���y?\}����z��@�r#�]�!T4_���gK{��Q�4�o���3ؗ�f՚ap�[)KR�G�{�'����}/�\� �IN�x:<cD	��ak�V�kf^�L�]E(wo��}N�/� m��@mY�ӱ1��� ��0����:l���W�rQ��5����C!Z�
�����Mq=q�:��mWyFl��FN��"���k�������d�>�K�0|u?lM��&δ@��$�3�{��n%C���s9�QX��Xo��|���_�L��2 ��$?�6]Oh�|�P׶� O��DO[��*�D:
[��od�����!G�d�9�S�܊u����k�:��0:a����Q`�i$����)b�¯��sB���W�b�`�u��ܻ|�{JM9��H͔߃:���:��������l� y_�Iz���l���F�W}��$���͈`�|nM���d�e|iat��4���q*�f��%���~��
J�fZ8AbF�)C/�u�:ȐNX��y����T��%����%(� �m�1�3�t��Xv����"�X����e�&���;�������m�g�-N,��(����f���H��L����[�gW	��@�[_���%P]��C�� ��I��k"��qsJ!�&�y��b���	�wX�e�i�<�4.]ͪT�	��9Z���ҽ;�*g���p�Y!-h��#����ŏx�zP�-M��Ȑ� ����hۘ�5�����m �T��1\�g��i��>������f*�;a9?A�x��T���Zݢ�����5��]�D�j#Y�L����������D[�]�%���5,+ ��*�A�,7)sE�E8\DH���'�pW��ף}e@~F��®r��K,��P��Ī��D�%N�W�E7�u��2�}"�;1��Z|l�F+�=��^^�"����a��S�c=*b���]^m���K*H�ㇸ<L p�ԥ�TԜ���!�L�Q ��Q�{	��G�^@�-�(i/�'i�108��*
K٧�(/�bL�r[ދ����!j� �2
HS݄v�ё�fۺ,�JMkj�X�ߡƔ]�y Z����)1�dm��M�$Le�R	�������M&�I�h�|�>��U���CY^m�k4���_r>��d,���)�LJ֕*���C�1�3�Lc�L��
LC���~jtJ�7R^�g��.�"^�8@}����IH���}��	����Q!�=�W�Tn�f������H	�³��c)E�r�ў}r�ۿ�]]ς�@@n���7w�Z��8������[���s���wj�U(��ؑCN5d�d��j�k}�V��֮��#�"խ�W��̸���#������	��"(�i�g��I9ד9*�.ࠕ���u�5)�5eo�/x{y5���,?Rb�0�*o��)HB�)��O��,�wzUU������LhL4�lp���1���.HO՚ݚ����x�����&t. I��z�C���������3�|$gIl:"��=��]McG|��	���w���m��!�V&J3N��,yO�g҇�IP[���`�hj�C{�L0�!�:�L��{1�����1��7ՙ�6�=�$�Wsi���*V��?�[m��a�Oi�F!�>�M��	�e<�;TD�K}d�4O��"����<vk��O��������*�tH��rf�Ҽ����caU)�L��˫Kb%qe�5GO��8�ಮ��@'�Ml���:p#ۜ��4��\�(��
�*�k����֗aċ!�K�_Ϡ���Xx6V���Z�����O���``���%i�rݙj���( ����m�5y�8��f%���b���mV;�u�~Q�O*#�P�4$��d*-WO�'r_��Y����-O�Mc�;n���dC���ް�����}b�u�������d����l�2�o���I�}�9gg�`�f���/�~�h/���x�"�|�C4x�Je��%Q�Mp9is�����������X$BK�(�L�K�4��J�0�~ ��UL�M�����S�]@�7�+x)Ȳ��Xb���K�v����#)�������k��uT�k%I�G�
s���r2�HHL���XWE��������Y��gf&?�)V	�f=�ɪCޓ�_l�E�=�+s�T�9��8C]��Vޠ �b�&Qpwb!�P�ń?~ܦ�G.�l#����11�&�Tn�-ʞP��S=(
@�b�����V����g�������s�mf��q���l�H��Buk� ��(,Hâ��>�|'���ۡ�!�7o�fЖ�5O��[~Y8Y�g�����Q�u�rME�싍�,�N;�fy�OKJKd)��6	U����2j���NZq�t�2�����SԆ[��,Є/K۵A���+�Cn��������$pփc���s�k��D��\"�Vn��.�E�y�Y>n��Аm���4�Uq*꘬ N�Q������ӶK6��m�T������6lxԭ ��S2_�Zʕ
~f��ǭ/��ٵλU��>2.�y�ZG�+�ͪ��@P_`�I�	����=�1P��>L@c�^�E[:�(�#�8�q�|cg�o�h\������.����~�����2��#��	Up�N�!u$c�/��1���SMf��$ك���q�Zh-�G����.�3)�[��m�a��2��?%���Ҧ�"V�DV�m,\�/)&��H�������9h�����'��L��g9�dq)^��l� ����3�� pq�="[,�Vj+�A"R��C!��_��.�E�g)e������f��	�ví���i��_���,cԾh,�n���C� �-G �C�-Y�+:�Y��M��y�׍���g���&|l^��%��_��>H}����{5����!�����#x�+�4f5>�H@�+ �Ig�pݖ����uɟ˟i������{��qb,Y���3@��L�9 h$w'�t���dn�G�xN	ſlo�+�������n�V��
x+Jn!+�M��ʖ7�@;�+�ᦪx�c�cO%�H�h�)����ꅕ�m�n���r��G����ֿ��M��P�{=Jo�ț0z�6�S<sR�x�F�B�j��Tn
����GJ��3+H�� ���yHIL4��e6>���H�y����`h�zUI��Z��)�Z��2j���N��1���NM��G%�ZV<�J<o����k�L�n��_�=��� mց��խDY[�����YC!rѡ4�3�����U��?���������p7�]�-�^?� �,<��l�ӟ�7Fpc ?n�����e)��|���+���]�W��鎑���8E����dh����E+
��,?�L?oL`����~���eə�Q�UqQ�x� )+�}. �74��!��H �|.��Y��c�f��U��MF��s��gV��������O��������uIf��`�˼�t�CA(���䠙2�n��*{�$��MЂ�G�����)��?*�Z��`+aM��Z����� ��P��ͩ�:Mn�S+p
�y��N�}�ʜ+}"�:ou�T$�y���y�aU��_�K�7�ƫ��ʲ_t�^��o�io���$�=�C�r�6򰧌{���U?	{���V�'�ɛ0���O���%��f��|$r�XbU�k� )��]�w�#�+�0>Hl���D��"R�*�BX��s��m��#��x��H���O7i�_R�[]ݭ�ubӶ�R�i�d�DB���~&�K�e��eueH����H�R  o�[n]�Ͽ����ۭ�>*���l�Jc��Ea\K�o"c)���ܟ~�[#\�&��W�1���#g�K�L�Lp��'�@���)a���h���g�Gz\OAڬ?�Xo�~���ۑi#��"��_��x'XK"��/A#T:�7C�m�$��+H,�Iwpu�}3��7��&�Jy��������L��m�����	�:�������*�g��G�Gj8ԗf�[��jF-��;�ޔ����L�o7��?P�1$�ͳ�^h��&��v�ǂ�y��w�r�n0D�C2_Ȋ�����JHY�@�h?s�kb����L��ςO����h��нm�xn�F8��`��¼��u�����v�{�;��	�y��ϱ�=�[w���5�xQ�iE[�O>^��NJ �~PK�L$�������|X�Te<+H���mm߶�݄������_�W��ˢ&��Nb;t���TPqxڟ\�,���U^� �$A�A�$H�,&��g?���y��}��g.��̐c�,Ou˵%�����T~���U$����N�E�y�"�u�|s��q\�٤�?�\�z�i���&�7a��0xg�ǰ�!xW��Fi��N>��.���N<r��V�or����z�$�֌���ھ��	{�*֢���z�Q�O_={Tg���i@ �N�(&�Q��)�	`Σ��t��q-�*��S�n}���ָ��ǖ�?Rw��m��H��1?BX�_�+4��Թ?���G5�hؕU�V�4}�E�VJ�}J���'�q����������p4m��(�G�"~�ʑSZ��Z]��k�Z�?u�����-O*��ⳎW�6����ے�1�J4
�,c��q�;ԵM@��zpe�!Nq;�	A��#j��ό������L��ِ����6Z÷���:�Mő]1;�ă]av.����Z�GAh�.J�mu�`��e)g6��c�H���>�2��!��0�<y�9S[r��Pz���ܭ����n|ES�Tψe��Bj�O�9
���b�*����ٜ����6�׵�L�-RV(e��փV����֫�5h�$M	ss���#t֑m����/[�����Gں�s�9!�6����y�]���~]�>+o�����*Id�+!^�p�]]!c
E*AKm?�kZJY�ضQ�M����䡍7|n��F�ȓo"�:_,��Qm��By�/�����lZ[I�[���,%���R>�#���g�e������-�!�#��%�V�B��
�E�}�LG�RAgID	��pD��~�ա�*�|D�-�Q^��TD�ϲ�V���܇Q�N���m��C�KY<��1�ڷ|�@J����H|��U�`�{|���a��A�R)�@�;o�a�k�~$'ܦC�����8	�y�>�	3!M�>�[	��-�UC�#��yz;�m���ʪ�;�� Rh�&5�%��Mx gXW��B��mh�l-�Ǫ�c��Wn���:�X��������YP�'G����ϓ��:n���Aͤ�߄�"��s1��Z�R��}������v���s3_;�E5x"���+������got����1:G#.�z��^�	c�u�a��M�kS��	�}R�[�:��I�����̤v�;�բ�J��*B����EЕ70�C';'�pc�d;��N�L�`��m����۶R�I[��N!u+/���$�n��V�<.R�*h���.-�`�Q��Ip,#6��.kV�6��)UsY�g�V�'�Ħ�A'���K�(����U���NeG� �̕7k.���aʹu�\l�����D��̨�I�X��[��ru'Q����J]!�/�	<�ˈ���B�LMY;�B���$��$�TQe��X�;���G�� !�Tw�wKl#��Y��������wF��6�S
N\��Cqb�]̒������C/w�W�W��5.��-�Nd�@��,@�.nB�BRW�_��R"(�`����,��+M��Ll={(����(�sT��<��u���BW^9]+s�v��sJĈA��QSb���
!5�����u)t39e|�zV��C8T�9 lg��>�	ե�Z�C��.
F�bu'N�&� �����i <�z���vH���R�j�5��Ua4���T]���e.RDs.��4��<K(�4q����b�� UW���.�>��L�_o�?R�hn�6s�mq?Ws찗R1�U�G�em^`���;�cR�!A��6=t��J��E,�p�r�.�q������9��bƛO�� �DyH��&�&�da��4���X��ve����D�B�%������H�Bg��"��Yr�
��<G��b��}bx�5�m�HNp�R~K?=�2��t�f��JS�p��X�'�3G�+��QG&m� k�,�� ��6��y&V���t���Ox�����4^Jb
�Fe������\dQl�76��w�%$���/����P�8�I1�+�c@��;fG�����g��@�$��GO�0i�,�0R��!��w�@�@��spXLk�&
mDߑv�PhBWG�'��QЌ�;!�D�}P�ɑ�CUD�@RI�L�Ax0J�%$�]
�І�aZY6��[�-ͰA�,���l���
V�K&XW���k�����0���I�G���d8fr���� �`�]�H�ܓ|f��s�����$bq	EM\X1l>Ƒ�U*�t.�&�m;p��٫��r�>M�r�R��
��A9G�!��_�H���k�LΖ�^�A�ʳ=�1I�)T�]҅���5�� y2��jۢ˽�m�o�Z���[ɡw����({E�2fP�={(�&a������N��xP���+E�����s�'�Z�K�8�;���|�5k�����3��$��R3�I�<#,��FxjJOxyo�iM6D*lM�5"�׫�����jp8E,�U�k��,a����S%5f�����������Fy�Y�&:�4N	�}5�4�ɞ�$ɡB`��<��ш��/�T��~K�)8��5��υ�u�x����e�.��|��w���PJ!��%���ף� ��P�k��Q?��	�P�1���z��n��*��0W�s8K-�V��= �֞��{�<F�٬)��ڧ/�����?ʎ�Z���I��Iq�����x��!��sk��eA�B��rƃ��xiB���l+�+mt��VV�%>xN��U_��+����(�j�NT��{�S�,u]ywH�/0Q?B�#9/�~%��W�Z����A��x4k�3��h	�+N�\9�������a��	.� !!xY�nV_A����p�^�NJ���0����y�'�Ǉ���T���v���)��HB�dU���+�F���F򚰬�6��y��ј�ԍ�Z&g2߸c*,�` R@H�b�,�U��@���Y ?r:xl|e:��7�ST�c_�<2ݝ�
G���֠e��t�ka��|l�U+��s�W�>B�x=�W��.Ȃ;����3%A
�(�~g9U�x����LW��qFr�nv�p�����l�6-�KKs/��.ˀ��Կ���'څ��b�]b�
g��1i��6�A|��;[׾�05Hz����s�e�ٱ����i��L�-�R;P:��;�O���;�z(�r���7�G���9����K�g'IKGdZ�8�T���mR��j�dY�x����{��n��k�ks���k۔\�xHp����[1I�;�!a6�	1�E.ؔ��*�;
HIR5�Q*,h�! �_G����v>r;�rj��Zk&ˡ�]�XճkWY9�T��X��i�WM�J_�x~c]Hg�w���KN��皀�g�>��BmG�b2�u\R�3ӭU��<�P�QL�l7Ga&DyO���18����*%���b"�wҨ�E3=����p�(��U�ag�<�ǂ��S�i�I%����R�ߪ�wh2�l>�ڑ�~�)�T�p�犷F'��^FТ����<������\"����qf���+��-pI���q����,�'����; �LG�i[�8U"�+{t�}[��]�`9e�������I�F�~ �<���Y?�s ޶K�����E5���@FI{��@S4�qósh��Wm[��C��C�ذ�i���A���"�XbWJe{N�@�Z�� ��\��I�W�n�Mt���0{X��9[
��U�g�xO�P�}��.��ĩi{���$;bqi�����ЯmE"e��5��.���Z�S���h��C�*��:^�8�IzeŤ(�li�:�ծ~x�������E��yY�E,�h�j�z��k �6U�����Y6�x8�F�|I��lԽ�Z��UC�yL���ʁ��܍�I�ep|����֮��.�`J�e+vb�%t;0C}G�%��mİr�j�����&
&ڒ�jML��Z��\jxs҇m����
���FŹ����5m6���e����D���Ue��U�Y��Q_g}���v�&S<l
�:�IBA�ܸ4�k����9��D���P��r�ȑtu��r$�cޢG�Q����U��Gb�<��V�ٵ:H=M�F��s�x�@�R���@�P?R���Z��m|&���زZ������!q@7W�7���c�hi��u��(�|[��tZ?��֘8���W����Zh�+B��j�v
V���qU��w���nO�����t�?%V��-g?gG,oc]�~u_S�	:s�d��X�[&�fMh%� 9��K�!�h\�)d�c���%�H���"��Ѣ4S(8m�J���.������[[q?Qmt�7]�||d��r��n/<�hD�gq�ɳ:��ʮ�Vwvv������
�N��	�S ?���ɟJ;PjҡNK��"�_���� ���0�����%��^����\!�P&��̈́��E# V�@�	m��
R���(=��O�^�ء&�cûNk���4KRc�^N*��#��0�5 ���⅜��'ޭR��O�ɂ$ �R9 V�t����8��]$��N�x�Sa�<Zu�B�x��a
o��U����I|�-��]���=گ,�؄��]���Eq*�I�
p��Ą��`�QQ�"����xk�F�Iۇ$N��3��z��J�ؗqӵiu*
.=�*d�(������g]�<XS:���I �8��~�I��bAɑ��a(�Do��8�pL�r�1��KS?�&`���Z&�%L|#F~0c���nOg(wI+J�/;�9��� �^�e��6v�tܩY$��t����h��J�Dʷ�E$MP��1Y����<��-A��Q����`}�ϙD�����Y�JJ�B����=a����>��{��J�����rAW�̸�K�h��eu�Y������_��ME�Kf-�yO�U�l���*I��j�|(W���DY@�ִ���A\���ЕO������#��=I��n{��(}�����iq-C�ʶ��gU�����Ww��R�I��NT�X	\˂��PH�<��R�$�ʓ35��bu�� \������*�P�-�hT��''��Dt���#�����YRB��@��t튑[����G�_.m�e�ve%�B�p8N�z���jswA�32ґ:�{��&����G���&OC���"��r�E$�D|H�;H����Yl�حCo}d6V��¢&�q�B3���ATy,��J����Rh��['�.@R[��Pz"�'"OS�w�4sy{��G'=�&�`���eYM_|c	����R,�&��2��ZA���AG4o�AG�S
�/�6��V�!��C' �G�=[G����w���}6���i�3���L
l�׹��4��wnd��*U(�CF@gT�:�ZO��5��%�C��[V5�1�!ˮC܌#���2L�7k�@�˚�>��~�\p&��n�j����\a��#�k(H�d�u�R�w�V�fK8�R��^RZهr4cn��`�K��8��fIh�*(��=��A$�	�F�jV#�G����(^�$��O�r}�?��g@�?c��{�E�P�қkt���ȱ9�p����id��������'̉�0�W��,�N7~+k��� ���kW�;HQKW�EGN0`�{��x)+䭝ԗZ�ը�G�|I����u�����`o~4���ڔˀ�]N���I%�.������Ao����]�mĶm�-��?'��g��OoW 6H��`���-vN���x<R�ɧgi�6̉���..��t�{�&�6�E�H.���-���m�� tV��h{�LQ_��㈰�}|G�-ur�ߕ���A�"D�^d.�c�}_ o����mJӸ:&���)�-.��ll�A�"Άā]#�Q�X��� �m���\��l��dm{'7�x>
�}��j�;����;�0I�)Z�͔$��i)a��^�{�R��[�&����^Q���ѽt;�l��Ѱ�틖jw�1�i�ah<A���T�:��Kۿ#�~�
׏dx�ow4��@��>.{�[e�]/GǓ��W�u��#G��>�k@;�s4>?%xQ���C�K*HP�K��Y�Ao�*�7�z�M�6p�j�X?t��d��gu���O�J�Ӌ-��{+�	
��o�޻�遾���,���J� �y�Z�E1�,aVNYc�����եi3��X�Q��ڹ�Yk���+���JAdy=��{ϸp{���=���z#�V�U;���5\A����z�S���uD�`����|E����R�����n��t�ֶu�����R]9��z�*\�#aD���{[�c|�LӐ"�m�z:t�L��S7�I�&�G��M![>{\�߷�$���3С��~}<�u�z�,�8��s�Ī�?@J�
Rs����,J(d��6f7b����1��3H�)�������qS���R۷�k�I��]!cd����O᝟��.UI/��iD�+��2V��ӝBy�5�F�=��T�f�kr�>5���{�
��ڈ�gc��b��C��>M��a�^��1n����#|���M;�fd̗�H�BV��٘���[@!9X�J��
����<xpά@Y���"3m#�����\&A
-�#�����2�R!��o�	ϙe3U;��0>�CF�:��+���o~��b���Zʇɬ(�1Ž2^>~T�!��aCz� ��L���GкQ�~Y��G��@!W�YC@�O:'����rlp"N1B���+O��͎�w��1h���L� �����\�����9�������,�w~u�j�%U�P'e1���W�&�;s���5��K����f�zh��k���}9�K������p�p��vV��l=���L��a���D%G�1Q����g+Gn��oyE���r3��u��ּۏ� ��$ע$љ�Yk�^�=Vڹ���C���Ug�O;��g�M�d�q�@BY���=������s�0)� ࢐"y�uSAQ\Al���������v;�@�qS@kZ{�s�2
�x�?i�|�s%�E�	��4j�Af��ɸ
���±)uO7v�+C������!�5������O��Hķ<�������
T쫽�����#"x/�a� �{e�'���Z��A��q�EN�[z�z��kJcM�<tzߋ�z��;˯-��y��t[I�s�Y�|��}Bx��ϣ�I���B�Y�*}�u$o�eF�W��[q�3mbG�k^���*�_.����sf9z�cf
\�r�ټߦ�J��پ��-�vߓ�t�A�o-��Q��)V34�ʙ۱RB��0x��,F��a�o��a�����J����#;�.��kZ(���-�j��ף�5b�ׇJ$�G�aW����3qo=�����ӴG�Ytna�=�^��S�ņ��m�Ā�}�xцj@��ӄ$��0�LO���;\�욀x�gi��)���Eq~��a���ϙ���}\��qsb7O�)6�p���3&�n� q<@��*����m�c����ʾ2g��P���.)�1�$t��M�,�Ytj�\���Z�a�	��wZ!"|�(~�qF`���eg�4{p]OK`춵!؎�0x�j́W�ʙ/�(Y���O�Ȍс��R��Y�M��iӀ�v�!S�	G�=S��,���� �H4���x��tK)"x9pW6x������3���,&N��up�1[ �r���K\��Y�ݢ���t*c�ڗ%�/����Tw��(�pm
W$�WiX�#�����/糮5J�$i����MM�/T��=7��ͨ��w��0c��G��ѹg��N&��c�f��&�=�+���c?R��)vY4H���SvO�C�[��d!\!��9��vZ�
��r��;�ߵ��ַ��F�k�`�<�_&j���XPį����;(鬴��� ��"7�B�DH�X��߂�܇�4b����#ޔH����ɒ�����<7����Й�wOt���l��$;�CZ��Ft�W���m�Y�BN�v�B8����:��s��k�o�c��;��;{����L\�(_)g�z�ϵV�hk�wRy~ ���W�(�������Y��yl�y9'F����r�D��E�"�X��Lѳ��f��)es
�	_��/�$B�5J�X3���"� Fe\.I���?c�,�2כţg���ݞu��-�ݺdy��Ϯ���������g�D���6-�N�����Vz/D�ʏzP����
���?4)NQ�`�I���u�*���ߥ�4]�mȩV�C핑o7��rIL�!���߀�g�j_Y	�J`a9�e�e�Y-�;�G����RsgU�F��ȳȑN5
~e��dg��]������
(���YG�,�9�X_�"�NA�CM�o��68� ����3o���a��6��Ev���8�9d���H<��?`��@�]���Z�Q����ׅ([4�w\�?R/�o, ���������5ytW�8\K�x_�*�σ:�\9�w������WY��̐₦ѣ4�F5,�����K���/ *B֋�c��q0v����f���twҺ���O)me����W���B::�q�P��d3W���Z���E^�$�|���qy�5�QW�GA�oT�}���*�����܉0�n��l��M.g�M�G����z�b�mPVSN�FO;M�oG0efbY�@�0yЮ��)�yg�c��g�czUZ*���>hlRj5�g��=�!����i���u���*?	�Q�bJ/S��( �E[����[+H�pW�Ђ��l�S�Q�����D���@��xS+K,����{exCŧ���ÙH;���+�\�[��upW��8��\IsGC܎�n�� ������23]u`����s�u���5����.է��^�9�*g��)�B���j�;�#<�KT�r۪nh�u`�'����,�<��x���|���T��#�B�ߢaY�\� _��ζt�z{���#ְ�rF�T������:I���Ax/��	w�Jkޡ�t�\mC<q�Ze���L��q���y0W!g�5��ѥk0b�?�>桶����l�cT6w�N%�PaWW:m"�oeb�}���Ub��|�`#]?�4�a��n�M�!=��˽\����� ��N��Ή���M��#Eɞ�Q-K�X���(A�a�gAk�,�=C�l�gG~�F�W�Kl���@�{_m��-�����]�V��E(�G�� |)5
!�%_�x΂���'���瘀���	 ΙC{\o���`t�����twx$��{��Am��*����,������{̵Ƀ}�v�ρ��h�)Ե��+�wd\�PLP=1a<	,� n����U�b��\;ĈrD�W��e'%�2�d���F��%�o� M!����_#�t=O�ǄIYFf¡�-���1k�g�aM�����]����l���I�k�Zh�E%�޹�1|8��3;C{t8���c^��9�H"E��D9鮢]��]���	��aTX2g�V�+5���s����1E��㎩���1�����.ׂ�� �nг��_�`��Wq�G�`�v��P�4{��l������\�V6��>?�4�Mnr���^����;X��>�6���C�m�u�C� ��6��£t�IQ�XJ�
S��ޮ�l�}�hS�H����nܠ�{Y��И��̌��Rh~��i�O�Wuh�4"��X mn��O]w��sjH����J��}�Z�<#�=�ȫ[��ݘ���;W=R�ǡ�F@g���
ҹ����>]��K����%0�	�d!R�'�n�\���ϫpj�L]߆ą���xB�6�G�uI�ႎv��F����#�pŷ�X���1�/u��_�}I!�\}+{I�V�x:�v��{8@��t`�"�@��i�����z@���ݿ����v���~%�م�U(�"�^K3�XJ��#+�	��qJ��^"^X�]���W���[�0��~�yD���n���ݜV��|�mT�U�MPL�wY.h��q>6�nO����1[�n�TmŵF0 ]�Sq����q�Q ì�*��eW�1$���,g�iAi��^_҃�#I[�v�m!��g`*D����=�d���jW"���܉��:ԋ�_�=�%����>F��g�����,����r�g�Z���ٳ�2�3n[
��ټV�gBo-��ﭕ�;����
ҙcB��hT4��eQr�$�Ћ��u�r�j���ͷ�ML� �?Av���ar�~o^-�3�`�V]ͦw3sS)�#�2�!�P�R��w��t����$mID=:&��6
�y���A%<�Je�!Òv>����'�Y�������M��֭!��n�|-4@Qo�HӭQ㍟:��r,�Y��i�	t�T��<��ި���h�=W5�z��W{x���Y;U�EnV�kɕ�:�u� Yp�y娟�+ʽ����������3������8@�ߊ�!.r�Q��o�|�|hG���7Z\Ҏ��?`�
��۲��O���ɠ���s��ƪY�kw����(���k5����׹��w����O[�n� M��fo��X[�=��<O�\���h�x�͟\j�[G�K?t���A�6[5�>pOl�S�F�mO������Ʋ��]G����I��{n��c�:�G�h|֨�]A���W�H���)�8�?w.wP���	�������Rx��F1T�qPܪY�l@�\\����x�ȏ��ʹm��`�'���X�[(HՏ�w��k8c�tԭ���=�R9�NQG����O���cL��2$�n�)�ֆ������,�CD�e��NXZ{Be����}�z�%��i<��@%���/{'�!� `�\���R{�$UĪ�/�����r^�%8z���y�:���Y�M�)����	R(�-t��4�=^<"G��&��	+r�.��R�e]�rF���{SYt�(��������k��&��J1��sow!����z5!ҷ�^C�|�հ���M6~�.@VL��E�̷X��s����f�qk��ΕX�T��㒾����q���ӇD0�R��x����������x92���~�o���"3��:����6�C��,���񷿳�9��]�]��}cm;-5lg��I�˳H��yw)Z��Y��.v�q��H��f��������� ���z8��S'+k���ׯ��D���7��W���)���e�V
R��%���K���p�^�4J�s^�`/p���^%
"Y]���)D�7�ȃ;�u�_�t���Z�E��I�����pSXA������?��l�e#@��D����x�#�\�P��w�G�1m��JK�[5��G�5��Bn�q�}�+8���Ű��2W�^��ص��)���>��]Wpdo� E8F4����z����xɿiwB�$�	��~a:$��� �ݖ��B��$bOJ~�B@�`�9lES6�o�x&�Jo�o�a�}D:Sz6��Y��A���2�H����,o� �[�Fb��\H�E���J `�;��h! <���7:ϭ�Vz�� 6��"~�$�v'x�=K9����|�e�Bt�9�mZp�l��!��N��w�:�|�=/��t/x+��*Fx@ړ�s �d�w!X9C��mf�X�����W��7�"�=���iȯ�q}��t�=YH����Z�ܭ����?�����������RR,��3���4z>��4���G�*�ց�w�-�[���;���1~���Ƕ׿�����8lqs��U��KX��WH��V�g�u���XtV�g��2b�7;<x�f��|i+��u;��j��D�9�ra�+��7�hLn\��_Yn�\>����j o#�� ���M�|��~{%�c��t�j�^>�Vr�ci݄�����J���nǿ��	�G���?c�.{@D�oKX2�G��꬙�d�Q�1��*g�M�6�A�Q{�� )b�0�H�Kz�w�k�J�TE���kI�Y��x�l �(GO���fb����,�j{X	���P�������χ�i�6��}g�½��)������^H��`yf}�z�g4w ��ZV���yeR�e�dߒ8]��S�u 
��*r�`��+���$>6�`�� �TQ��q�{4���pc>�&
R�|>J�S��(�`�}��<3�����6-=5��u#Y9�͈��;gS=��J��)r'�,� �8ە��(xhx��Ρ�դR�Mq�S�F��)t\�>��s�R�n�c�CA�M��E�Z��N��cP펄��C�^	�5�S��.Z��5`rl��+��[=�n��]m�`Il�����0�����t���7cI�T�9��J��Bt ��q"������=Mo�!�����փ�S�ӟ�e���QW4�>P���X��d�Ÿ��gT�F�[�S�L�`�Ϥq�Pzn�O�PzB[5�c4���f�p���� )���1n^�]����b�ܔ�_� � u	�
Y�i�1hpB���� G�c8/�Da�ԗ��9`������i�n��E�L��B������N�����[AbĽ4���~%�4<>6��dy��� KI��T`��utS(͒E�yh9���S��j���T����MY0|�̟H,Bq�Cyx>��H".�+o�pa��V�H[��"��"��ɁD ű���:�G���M�� }�Yx�
��"C���4~�7��e���/1�ĘE�E@�5G��#,a���Ŧ����d(� [�U������Ck���<[cڲlȾ^q���,
�F��@��6E܃�$:!v���+Zᗈ�8TG4�pY�%�2�0�;�Z���b��P@f�CA�7?�_?K��{��.֜��O�����n�=�����N�����k��]b���D8~-�3��VTw{��RA*������o��=��w p �?�^�1r�G:+5 Q	c֮��P�<�!!������o`��Ĝ�1��>;�>���� �?�ii���6��}�m?￦>�{��z�n� 5��O>nv��2��^�4����ƣ
��S�uA�oݯh,���{�{.�ZD��wa��֝�
�j
��_��2�,�>xւ<:j��)�kG��'vg�NA;��<��O�pq^��
3F�;"�+NZ����㬇�\�<*A������w��N(w�ϛ������p������	���xֳ�p�E% q��`��� /�^��7���v_����H�:�M\���n� YF54���t�ⷀ�3m"7C��"�`�j�&L�E�4t���N�F���yh�s��N��?q��Q����&$�V��3f��,Z˥�!�R�)��cZ�̕p��lA� s�!�]�C���4���r-����v����r���³���ȇ�U[O��+HD�g��#��E��&��������J��L��߆/GA�Qmd��	��Jm� �OCN�Ư[� ��� чY�aE��C�n��)$w�S�?3(��F��BU`Q���e�V�L�V��x*X���Ľ�R�^Aڑ~e˸
'��!������[��H���^)d�t�A6��Ĭ�>�������'ī)����l���Ӗ�a�YN,2р�j��d�p���𐻭��w��q׉D���)��_����k�1@�SPsH��aM1bFw���9c&��K��$����W`#hy�<�������Ͷn�|����h��Z[�9�l�Bh�n����������g�@�B	\er��W��|����u�jGt?���:�؅�N��-�۾0��]�Jih����]���)����'��RS*kI��L4�He��,"����Ш녤�'���n�r����
�.�	�S�� �rd>�T������v�J��I:6�?���CE�v��<$�j�<���
t�:V졹;Q`�EZ�T��0�yG���V��t��(K��6yB-��B�2� +1$8�O�_b�#m~0vx-�	`�GƇ�c4����e�p���"�n4e�V���R��gZ,?P2�͙sJ�@��%xg�F��ot�{gx0��B��B��-c� @�9~�Ţ�Vf���4]�)��L:��`�a�`�l(w
�1��W�����\O��wͺ��k��k������P�8�Kc�eA)I��f>tX���uٲ�vG|;�{=���=��Yo&�u �}v��Q���ڭN+O�e���ل!�� @���*�1�
9W�%�r��m����=G+�����u�K������q�)P�Z��{/!Ԝ�?�Ÿ�"T�ͅRr1�r�o��w��0?��E�s�ulr  �Ħ���}Y�����H���-$��,|wKI������?���ƭd�0˙`��P�N5Z�YZ�}�ȓ�@�!�s������H���P7l���J)��1�~=�Ũ~O�������6���9H8bu�@�ɦdeO�Z6$��]��v�<\�҂��HY��P�#�l7��Tv������� �L]�	���..�0���>�`�ٙ����[�*��E
2!R?8�`h��2TL��ݮN�~3�3OZ���}l^P�h/�_#� 3��m��nm��!�`oH�,xh�����T<а@Nݑ�
<+�^��z�cQG>p�)���Dqq��dt�"��-�_��`���]��n���,ǴMI�B�|-��A��
6մB�j;-W�B����Q�����L��T�R>��"%w� ��u�.x�����SX��Հ`Ҫ7|Zv��Z��
�_\����w�-w�>�%��<�����k����@�J�(sz��d]e$3�\���^HK��z"z��?��}�㱍�l�����E1�
E�8�RA���^m����	1��O���*L��i!E��'!���8-����-�w����Ϊ�Xr����#�/C��쨮�������l�� �jW3�2�;\���
�����+�~
R�Ybύ���}�$|�@2�5�bg�T_I�8��g��=	��c������AUjf⏘��-K���"����Sޓ��h�OH�;*!$xC䇝G+���+�?�X�W���^�[��U�G(�q?�3����>�.��)�%�cڮT�d�	g��9p?�cM(<����Y6�dI��9LoAz��VM��M�����,X:�[��P�|��W��9o)M�k���N>�dY-�&d��%����: �2ULߖ�?~0p ��m���~����j���!(�z���ZG���@�'����|'P��u:��]�/@�k�R��!ò�����zgi,|�|������ܟ�r��|��͈��$�����Bl�'/�V��&毼���q(9���0�D���5�nKx9�7���h����B�w�z��
Mn�����Ȕ�Ao�����\QVG0�
���K+W��v\4N�qo�OB�D���Fn��?�2��v�@����^���e�RIѼ�z`��0�b���S�W�O*�D?W����@����^_a���O���e��-�D����!R�ƮQ��!#�۬�ă���~�7OƷ����V@��2"���>�QijA����	�����<On}24l�SKp�΋�難��_ ��U^�ȣ]�W�w>� �4�hA|��f����l	���η{ �ؑK� �����\A�!����h��x.XW��_�M���r_i���
<2����> "��\~�U�1�[����P�����Y�b�?Gi����7*V`��~�a��"�Ve;��X��T���a��T(�d�	U�Po[}��g�k��QvU\�0���J�{J��g�`Xƈ� ͟͠�co/���*H-l�Hg���v�4ӳ�3�Yp�`,�ZvM��Y&n�FL��(�f��G$c��V]�1A����h3�~F-��	1��Ӯ�ӽ�%�z�|�iۙ��	�+]D����.0��xd�eYķq]�I���R�a�-�X8~ra��sծ��`�!|�$���[�~m��Z��������ݾ{)I-���BJ/�d6zP�@wX¾n����H �{ѮQ�QE��JV�x�h�	��q,�p�8k�l������m;�ϋnt���ݾ𱈪x��eB�g��,������9�}�v���;����a'E����4]��?1+G|w������O�����e���Kl�!GF���݀&�v�2
��q��T�7���K�{*H��E8ꕱu��?��vo��ߝ�[�U�e����=J���Hĉ<O���`�-�T)�v��i��~��I.�m��J2݈-��E��Ɣ���L"3����[��<��Jd�G�.���7��-�,r��f��E8�s��^��-�6~�:�1࿡o&6l͆"��j�S.od8m�1��.�Y��
-�<�j��v��4�)K�:�Ў)�b�ׂU����H5s=�X���ɹ�T2�TBFQ�8^��nB�~1x)S~���9�~5�SA*f����h�=�Ty������;����2��������* $�ǲ��,+O�ƛ�����4�-v|���Q
�K8�hYW(��?srZ;�N�fXI?�X�F"�q�o}�הl�Jw�HAL�)^��������k頥��4�nr;t��=���e�3�C�WbKZ�\�AI�Bx6�,a�LEJ�2�[�nk���n��	�!�W�6��,� hF/e��>t��Ꮂ��
:Dd��t�'\�r�{5����~r�A�ĪM���'��i�~������8ZC	{]}x+8w![�I\�;ͯ�4�2�����
�j:0aT`�h��uN+��*B-�;���J�.��SDAh���ը�B�L+4��� \E17��� خ����m`�-��oL����;ͳ�yo�OGW8�+��
�������gɞ	�T��?�'g��ڕrv�΄�9���},�x=?9����YwvAG?��g�c�k�7]q�P�44~j��)!}tm�F�� 3�r���{T�f��J����R��VDʛ��y:�Ĕ� ����\��ZI.��c�v0
aZ�j-�jr�_\�9�������y�D������ZnE���7�/BƳ��P>GwZ�g����{]�Gd<ɭ�N#�{�+�t�o� ��"�̾'$�*��*oԵ�@���8����s�@E�!�W���� �|�d�#(.n���
�����_���ayO�D\S<	�^m��k�<�Pр�^_F�\'g�9���i/����?�0}���4h�q����9B��4rR���$y����d�d��I�I��o���0�k��u)��
��9WAO0�;��8�i�1 ���oK*k�v��ff�52�4�,Yn@�%��P?
����x�t��v
�&~��X�~�[�{��R^�(��.�D,Z��ql�K/��W1��z�ҳE��	�o���6_�N�oY���;H��Q��~�7!n���Ǖ�<���{�����?Bú��/kbl�Feqe��ߢ�l�(c���9Zx
��-���}:��W&�ƴ�D_����}�ϭ�?�ǘ�����۟�a+�m���YiXޔ��Y�.�;��������i��m��m��H㱄/���e�ʡ���706==nf���:�yV~v��Ϻ/�!k69�r�������W�`2�Pce�4��Y���r<�hMQ��a�|�*G�D���?]�7Hk/e��Rh��\���w/�k3`!*�C\�+)61�F˶Ȝ{T�]i��LɸEt��8� pV��g�4��d�r7�;ݻ,�߄�{�P��$S$:�|��W<��s#����}�$�@k\xpC����#�W�f�����@sS��;�j�-/��)H�㳄����=��'��J+%����֔�y������H,4F�3��u5�q~T�}
$A_�xX~bu���Ԡp�BxO ��w8��]����|��WjPg����sa����AaZz��<z`X��Z�Q������1Hf�����&hhL�H/�8'�u��?�&�A���T-�xVO��	��ā�4�s(J�TX�09�"W�y�4�̟H1�۱ H�~">``��/HC~�U�r>�5�)�!��1y�bDpK�iM�����b/�"������D�C^+�K1������b�8�Yإ]�b��)�ӻ#�/���63
�Y 2����i�EZH�\��GX���-н0�r�Y	X���Ҋ�U~��������~����
*-�����ؗ���D%���T�Z��8\����k��,ݲw�883d ��­�\����K��af��)��?�y��,%T��%N����.��uU��qʮ|>Ȱa�
��E��m!����b�-el%���.Zwd>�U�H}�}C�����ְҹ�d���u��2�Z�?����]{��=x�Y���B�O�뤢?r�Q#ʋ���
R�6-!�KD�^b�s�;Z�%���M�_Ыx�n��;W�RD%
R�*��ڲ���+�I����ѧ���A��+�������&��`q=Qv���l���bm}B�t��@����A�Q�a��@�U����szn�������uB� *�:�rp+�"�M�uPxdDR�6�1������ͦ=����ot��z*�r�}���D%	����pF
����X����ݘ�����0�45Cv�{��sVmGF1(+S�W����7��ٳ���G���M��DV��%�oW���j��ҋY�=$6	�i�-ʒ��a�j�Ma�}�<Öu�ڊB��=s!D�c��S�\Ƹ�"�e[8��2(p"�kK���p?� ��_#�|QqO��:mC�	�"�D%i;G����z�Bg���n9-�x�J3�<�,��#�k�v�����,�}R�=&�ƕ�R�?dl`g��?q�(�'�k��"P*�"[���<�c��5`�u�q��O�ux]1�j�	!�p���=dI��������m��I��Wu �1l��F�3������7cūb�wa�2�t�5��������ݕ<	�%���<n��fV�;6�D��%�퀽�Ǐ��Ih���%��f|倾ׁ1�ݧ���ƠI���M.+��z�so��O�%�����W~#���G��=��50��e����_�,O�̤�rDs�&�15֢�~��6s�,U��@�����6	$�4��u�T*u�M�d���,5�k�%�3��w���)"G͢���, �g��r�`������1\�#xȕ���щP	b)o�
�� �Xo�hL�$J	��m�_h�I��&b��5���������S�(g��l!�a,� ��`1�d�N2{k�@k`
G2=�ZX�����X�G���Q$�ۼS�g,��qr(��\���?v���W�vJ�@��p�i�ŊbmŨFu0+egF_9�F�OZoܭW�8m�ή�3�&�/L�?E�1�)~�K�&���n�f���5�W{�_(�Y�&����]ѧBQ&u�g7���� e�Yu��=[�(���8FH�~�a�Y��%��fI��/^�9ӂa	��+�*�V(�JPQ��:b�Ĕ/]t�p��t@���5�9Ft�s ���ӖT*z�	2�T�*��C�P�ڭ�fä$����F�'
b�����������kr��5�`�(f6��`����A-쁑NL�;2�WX�/��+)?E���r���^�-�?��&��P��t�!�/.L�A=G[���l ��*a�[�gAԡ>Pe���Z�0����fڹE����'�8i[d�U��N3�qM��ָ��Y�����C�z�ĨX�m�����qL6��,�����ks_�\&UC;��|%�3�z��0���p�� .]�B�����;���|�д�W���{�F���6���u�.#��%�?�muoudDF*GY���XT^� �3z��X��e
Қ�7���!l;���39)2\�����s���Zf���G8��gqqt�D�9Obv��525������ǭK^?��^��5�W$�ew-�i�a�w��9�k��k�G��.��в��F������H�Af�� �����N����D�䐋!	�ug �9D�Dt��[�vТ��0��G�Pjcb��V�Lh��q�!3��� �_`
͍�|mF�u��-�p����Gxx�Gꬁ	���
A�����������`�pf7 z,,���Ϫ��t����VB\yWw���}��B-d�H#^r?66$\����m��R�S��c�k:�(1���T����]�~����W����.�n��?�����#+�T��	y��O��^�����s�E !�7���{���e/b��wV���d�#�Zp�R8@YQ<��N� �	֝�ű��ԝ/���楄r"d��o�PcR�j.i�sR���`<�y��Wr����q�k+�|��(�&�l��w�v�.K��I�3�U����2�/��%&Yo�������73�W:%��`!�l��w����\��A�R����#�!gB#4Ι�ݠj�w
�x���K�� ����S�v�Ms)6�׺V��i:iad��.؄BsBڡEpo7C�G'+*n���_� v�@w�%��(LR�v�5�:2z�!���!d�釕lB�f#ޱ���I[3#����+.���(�@���o�	1�����*9@���׾S�K4ly�w��*�w:��{18���V���I�嘍9r��,��Y�b��]C�?C���4!�ܗb�k���+�e ]0� o!���W�B�귇��Yra��̖�,�.$�U�-͑>}m�]"��no���v��+�>�Q$��b�*P�������o���Y��������� �3EH��������)�_?b��_IX���N�T4�B��x4T.j�f;Ir-UKACև�3Vѐ���������nt^�)����]�8�$׺,�2_���u.#��R�8ީR�a���@��r�<C�1��-ߛR�W��]��w1��[���e�mys�<[sܚ�
$fs��zhD#,��=�C9��s��+|o��#���Kg��nQ���Ȁ��GH#�i�ȗ}��N�'8('2�T>gT�_,��5�/�z*xU����`�G�clg)�g)Æ����&�&.��u�O�)�2|�KB`I��R
1�ǔ��Vx>fFax.*�ǋ�J�i�9�tk;�������e�:_��3���y��_�Hl�YG�-�!0A��5pz� @�Y ���mɲ��ba��e�#��@�k���*nc���_�&�M����1ɐ\W�҅�񲻿�h;�!�ш�0���SPΔ����tsd<�F�ߑ	�t���δY��+S6fS�����~�����ߏP�{��]ެ}��^�4Ğb��Z*}�XxZ�h]8��5�[z��ƿ�ٯ�����?����Z��M��� �̕)�YfE6�)/Yikn�ndM�����d�4�\2F�~`1�Qv&��n���7D�'��݌���!��_ѝi��T�70�85�\���H�N���&Tϝ�$=�
)�s�]zo�W�為<
)�������ϟ��������=�ܬ�	��K��"�2�<:��Q9y�r2Nj�ĝ�/����/�ݜ�/�m@�ya�\���}���7}��_?���}�b
Z�D��ej���R�`�c6�L[��Y��o�>:4�*��D]F1��]����f�͂��+��_���&/.��|R��i���yTEX X�0P3�\�{7�rA'"�-뫭�h�ߨ�Y�uC�۩����g$|N��H9������$ج������������\y�� ~1�<�Z��D��9K�y��Z��x���@�ʹ���4��)й���p�L�_\gat�B�n�?����__{J\0�ŝ�dqS�2�
=	r3q.i��M��+Y�����0į������-	'7A��J��eg��:&8�>�9@�.�������J��2/�ٟ$���P��"�m��Tً��~����û\1�zr�ʮ��1�K��!�5�D3&��^/\nۇ��|�|��������?��?�c�y\�,G�Ҿ�ϻr6�ͥ@�}��f�R�@{�5s��E֌d*�Q��m�S%�5
��������!���g!��i�F5�93;P,��h����J�w����G�3��!Hۙ"�������
�?���	�-�s`��n��ٛE���Ab.� R��U^����ҡp�#�K�4��}�g������m���3��HT�X[��=� ?��De� ��H�!{��ؾD��|;���������Yw��iw�kH�Kt
�:\��HC�+H^T���aiY;�����`,�.\Ϫ���>�-����L�R̶�A�èEҏ��'�
n� m����������I�9<2eg1rr44Z�"A+�I$��@���'��I~�`�JVE�Tg��\�3���Z���1kq~��?�o�<9c!W���Ve���(��_��'UYA��}�7�B�W�R��y���Ͽw6l�u������1sJ�A��+{�"Tf��+�Ԃr^ԋ���|������\Z��&!~��~����|��:�h<f�C`�*��8���qbT�寿�_?��W���KD��Vq�^ˠ��v�Ҹ��Wa%���3�E��:�v����f��l�$���w�4�l�����uDM`Yx�녞B��)�˿7��������-y)'�C��GS���͉/v,L�R���dZ�ϝuT6*^����Y���\�K�ZC��@�=��{?��k��w�h<�a*��"��0��_�a'/V�뛜�?���_��H}���.'�Z�\*B�62�QW���=����\0�"�}<%˜E�<r����0SB���o0�7�|>��/�:����������3p?i;��o���K�-���5�ܪ��F��j�'���xr����eWj���φkI^	l�r����Tx�^$Q��V4�ҿ��$bm=@���]�"���6@�YӢjCnF�J'v�RD7S��d��/l��хʉ=?;���3����F��{����СDc�1ځ�G�������.v�2�����b%���idK_q��=[�$cbh�K���\�s�L�?y$��DXG1������y�4Μ���sG�B�@��H�n��_{������V��
���1���1����x�V��b'$Xl���LarI(݌<ٚGJ�(��4��+�1OZi��
l�;}����B>Q��1u�P�OS���S
	[1�Q@i�Rh�����{
�aa�����o��Z�X�~�ە�zE{�5ݱ�GQ������g�y/"��ݗl����Sh9b̷ю�Ӛ\��fl0�qUb�n�z7+��#��A;ү�cb[�K
ڳ	��E��r�W�ɝ��h��3Z�,��L/e�r��]�����?V�Ef3��d�~��L�^B\'�*�9g!�I雯�2����	����A��oeIYm �}O ېx-�e^�Z}`�&�^��-�Vay��2HgF^8���o"1��b۰�I�O�h�%�����n���@��*���g�,r�-��J�p0�S�.kq�ךW�1ܻ���g֭�L���m�Q�H���{&����w�X�D+��]b��h�VV�3�Z��Y.�l����<^>�{G��w�Zt{��������i�	��v�������>N��6��� =��~p�����q��|�5�8�n�e�Wh6��^ֳE����:�����p�H`����n	9ȍ2!P�JJ�¦&������E��Y��*�@��X����B��4�C� /ӑn� ��x�����4C�FeEy	�Ć�u=��Nߓ57B ��r��A^��:Z���I�X�&"�m�����������V��RP��Ufb�'�#b�0d�[ͅ��z��u�cN��� h�j�}>��Ԥ�0�tےXv��ʐ�]�~�b���{��ne���y�d�����a�R`w ��R�2`)�.�gmA��߾�ܬ:8ك,/�Z�[SZ1�&��9}�<��[��?|��*�Hn�)�c�q���r��ъ	y�r�!�'ڗ�`r�<����+j`�H�x��m�4���;p?���Y��AbM͈���&%�K�Sʠ�JrJ�xZ(:�x��,���!�w��g�p���a+�n^�
)��Z	D���Kg�·�d�se��bd̃Vv@S�u��vm/��̡����5��I�����t��T+4s������rw �zeM� Sql��W|$[h˨�D&�_�򐐥�ZjM�!q�@��+
]�C'��|�]��ago<^��C�Jg}b�Gg-�31���NO~�/����Go2�W��� �v<�2��6s��,x���[�}�9A���U�/���,h���:����ȱ�>�;�j�DN����]Um=[�	�$x ��5���P�H��YW>�lR����q%A���5�X��a�����u]B�9zZ��ʰ_Թ��)b��!���t%�B��!M-�ּ:@M}P�Λ�&��,W����p�R7���i{��Vj�m��'���P�i[�~PZ�pe����C�΅ʌ?I�Hc��tGP�b)����n�-+�Ţ\�"��]9hR�� M�d��t�鏴�~��H��'�u�-��ë�W��G&�'�Ѳ���)��$,�@�g�VJ,��^"h���3�GP��(�>"iS{
<x��3&@!
��U>��rr$OBP��%����B���sID��Z�[e<�|3ȶk՘:��X��ڍ	I8�4�|�Y�;C��_P聴��[ �����f{�'�1e	��^��0��5��^�M������ ��"3_W��	٨�{v.�\>�gꆍIcc)l�]����k��/e�҃3���d�i6-�5�)%����X0�2Ϻ���hebT\���I`�(�ή����R�T����l=����|
��ݞu-F2����c^��ʉ�4��n�/g.���Vn� E�+Or�q�������@�Z� qVV�m���N5��������e��)R��.����pe��
�L�\Uª� +NLc�㉫��)הN�v-��Q��ǀC�ӆqY��;�� ��JCQ�l+�t��Q'A�⑃� h����v�`�9�Y|�4cp��Z��1�^���+��N8� ��Ra�I8��p�+��F`n[��f�܆���38�l���}�n:�Xm��v	�d��""Ж�;���4�Yi-�=Ŧ7�T�܍�~�w�j�;3cSs�2m���wN�A���JQ}Np2>�!Q����ց��ί�&-K�m�_�bzQ�s��NTzJ�e,���!S�O.?c+3xp��L�B	�M�UW��NA"A,����@��JFfGYC����M��"J��'>Y����ɄE�^}�Z��B!pܒi�~4��@#���^L�]k���J�\���ԏ��9�2���u~6�F�(��c�1n�2Zp���T�myC����~C�d7@:T�~��!٬�i�k)f^�z	��*�ҽ�]8�5`1�T���ئ� ^�������`bZ8Y�9I��pM�	��nKtϐ�r�IO��k%Nh>�����.����c�1�`pwi̪/v.��D�2)D�p��c�<��٣xBK&�����o��v���\ϱVy��VF�$��9��@�Ĳ<���t��~��k}�#��W¿W�\_��o��>	����s�G�C��ܯTcZ�Җ�!��A9���ma8�(Y˗zo�,b�G���XNۭ�J�[M�-r��X~M�8�;�)8���7�'4J!�l��M&��Ӽ5F�]c�U�����n� I E��*�5z��DS�UY��"���LX�u�T\{� kp~��8�=| v�f|�,lu����k)^Ē��s ��,S��^��[���CD�S|Vl%�,E����	�$����,p!_�]T��زrx�a�Ā#�3�J�рm��#X0��P�����iA�����59�<ES�Z<�$M1eD��P�|OF
&�^�m�ÃB��4�;����I(��8�t�^,�J��_��d=yV�HSQ�G �N���:C82<<�p5c�V9D�J���Ɩ4�\0�um�)k��$1w!A�!�/���5m�j�+�C����g����ɐ�
`�E��>g�sb����1o>��J�k���/lY�DPc]��uj�E�#�4���T�#h�ͨ����!��\����T,0�WM�0l��������->X��w,�Q-\�F)�2������T;����&��3R_!���>�o��I��)rUOAh�A�&s3�c�M_S��Z��85r'�[8t�ZXkf������T6¿���_E�����Nb�$��q���PC��k�AY�U���o��aG{�F�֒/�2�ۤ����y��^�>���/����d24�}l�qč���M���>~��v�@o��P�g�ŝ����
O�w���(�+�8��i�4�a`ef-�o�=��[��F�:���D��f�X����3Eb��]�^3��L�"׮k4��a���k�Ȳ���لJ��Y���� G�"kS�����-`����V�	�Y8�'f�����GS�X5�Y@��ޱ��\W��mȋ`�?��TYN�õ2�:��P�!�Y�Y0���t1bs!�ڱ�mΙ7e��L�Q�\�B!��I�I�-!� ж��?��3��Y<c?��M1�幹���/C��A'�[Y�1�yh�c>
���Dm@�/���5���M Vo�X�ݻf�+�ۖLBh��WK�O�3;�V���v
��*�m%������---�K�ؽm����]��鷵�A����qve��+�)|T��b���74��\�5��ʑ*3�5qB�߳���Q\�ra�;zd����A�wa�2S0��	y�r�#�7N�a_�w�6]Zo�	�zi~\��Eijd��pM�et]@'	ϷZ~���|��:ˉ�I)M�[Z��M���f�+|�)96�+E���6�Љ�iۄa�*C#�v��K����X��}ֹ�V-�}�7�ؐ]B\ ��2��Ha��*�UC<��65�hQ��.d�����ժ���5��@��c<�d5����[*H��f�#cK��s�,(So1TK0$zX����j��`���_[ػ-q ��K���s�6s5��@��?�N�f���Va�-��k*�Bh
+U����?�ĩ"��z���ZߞH��5V$V��t�ÅHp�9��Z��m[��-�ٟ2��D�
(���(h�UY�s���H����&_}�P:&�RݲZ��|V7��#f�c��f}���e2T}�Hp:ȍ��P�	�y�Jg�a�i;	���.#;u�X�6��i����)k�k�{o8����=$�hɢ`���|w���veI��H#	�Z����,����<Df�s����S����,?	m����g_sϖ"��|�e����>���ۛ� G�ˇjSɲ
Lo4hT�n=��+1òج�I��-�0-��G��c�(a��h��ںv�#B1�|�s2\L�ޅ�����v�ܒ1f{�Cg9��P��3ݨs�)������ǃGz��8�iݤn��^8�H�`\�9C��  R�ҩZػ�r:�j��P]��I�_��F���q�]`�;�u-ް��Ь�=`�Y^��˸)v�곶Q��[X�꛹V�o��3�����s��l�D��Ǖ��H����0sza��=Cy�R{�P��z�ʅ��=Ç]B�x��h���G��A.��mz�@��eģ�������]"�ū��'&M�sF���W���5��G�N��+�
�&ΨF-���1��z��x.�
����c��J<+2���weѹtZDy*���Z�E5�����K�Wj8��=0�Ǧ"	�+5�zE(>]�-	�x�q��ƣ�|���Q
-_��W2i^�8Ny-�_N|�}=�e��yנ���l?��?�C�o)�?�37�|n�;�g"b��� `T^��}k��T��J�w�
q:�����i��6�p�����$)�yH��/����Qӫf��b��9����wb,�٩�b#�e%*@/0�4��ʽ��_��e��,�8p�����J7�ʇ�B��P�mN�|���ġ�P�C��Ԗx��E~ �ɚ��X�o��T�Oz�rLC�?�ƙz�?�mi����J֘�����w�]�W��í V(H�S���w��t`�[w�a<�����d�nyρq�k�� �J})�,�.���p[SJ�B�/�JPE��uԏ�g)|��U�!�9 C�{��<��M�B�������a1��n�M4�۸P�BI�AH4�������0��Q�A��i0s�S���]��-�<���`/l�Ba��D�������ZRr���S��{�8n��B��Dp�bn9 ��N?���Jy�\�=�=��+��"x��
:�lt��*<0�̠�\��@fI���Ϻ���M��m��d�,
�i��I�����Q�% 3`��}��1?<
.���6����|F���#gLᵌ�
�Rf��=)����KZ13���Z�1bT;��W��ּ
�Pނn�?��]����%V!�#�$��� ��FK�� ��T�j�o�n,c�ի�p�8���n�:�����/�"�M�t�;�,��j���$�0Y�N�q�{wl �8�Q�|
z�%ѹ�t��ʛƗGe���]�*�k>��$|�,��"��U�s�`�� �ƀ�����?&�/ҝNA ��X�.��Ck��e�������6�d?����
�8!5Od�F�9nl}ڐv*�7pQ�&k�jOq��_d_���r;�~ǺSצ9��֜�qI��\���es�a�lM��\��K����͓Ç�.Y:��]Be�i��8�VA�[R�__Q*�)�(��^i9m�)�Dph]��Ԋ���,bnPcz�Nj)��ŪP<o�캮����9��_/Ө�%�\p���R�����,���Hcd�Z�1M�����w��4NJS��I+g��"���Б�ՆO�޽���(�>��$(�5�(#�m�]��Y.�P�\��v���5��E��|��xU��o	���������;����i�|G�Ƶ�����������Q��O��u.�4
Kx�o�S̿u�K���*Z%ѓa��B�wp@.�2Ɗ�V������\N(���z�����y4~-`ckS{�RA�B����w;,����/�x����-��b��/FZ����N��,e�ǨE[4�o��!E�n7������Tv��ʰꝃԝ��=2����&7+�p�����DDta¦:9�'┨���ۼտ0No�������/v��B�'�g%�n�m��k@�҉��Y��5ź��'���_�Թ���웝	��@|�(��[�� s8ڞg�-�x;#�tx7/��4/ג��ƅ�Ɵ<�ǃ�1z��T��>f���G��6d����rt��6X���@H`)3��'*�j�B�A'��n� �{�����A4N+�j`<]vc��6Y�M6�m^�8$�m��%@�+�	�05�H<�j�Sy�0����ѹ88�L�ߟPߨR7&���Ya0ٳt�:R.p�Zp�e�Qx:.��iѯ���qh��r
��gҌ+�_y�3?��4�>_ˣς[+HY�|�p	��gN���}�0����*ȮO�=s����x������2^�Ɉ�}E�s�i�����vf��3VK�k�ӫ�ׁ"�[^�<���=qT!qݲ9�IN*�&�u�m���e�y:�p�����j�a�b�	d
�|�/0�	N ��X����;�e=��P���y&��J��l]aѯ�E��Ĭ6.��b�"��^K{�v����y��$���w���
��v�����q$$����	F�{�=�}�{�  �E�le� �ߏ��+�) r��?W@M.ז{KR���Q��d]�7�Ұ�?��k���{�n�~ǝo=ܯ��DoM� ��"+$�,_��y��Fg���<5���R�,�)��*��B�쀓�{�lٸy��ےxJ�&{g��jh�w^��-��T�n�8��w(��S��W��r}9����hh�08s;H�C���N���
��4��,�"5���u�(.�-q�e�~˂= G�-�y��P|��co��a)*����8�g��g�ir�H𧠟�k2�����f�ϟLg�MgT�Ɨ7��-��w���
ꯡ�[7��\9F������h����&h��#���P��c�P�87U�p�F;�fw�4�GW�q���J��[ &G�L����ͨ��ʩL���!��wa� �>-��I���~�b�y#�� �߿pg���=Vv`�e�Y4=X�;�IK4�^�0�T��b��aw�?+#��qD��|Q-��m}��jW\*جk�������"��}Gܕ�|��4�+��i/%Գy�AnmT$���>SѦ5�#o4��A	h���@��L�w����'/�l���p�#�vKa��G�;�����g�Ⱦ���)���M;K���e@����o�Y.���)x�q6�L�Y�y�<��8��X�A|д��N�[*H�������-��L�b(�*;b�1�%m헊ޟ=}���b8��O���[)�
��v=<h6�rg��!
�RQ��}�r�߁S�G����^A�ƴ��4�}_u����QQl"�1$4T�Q��]{��)ǋ ���4vy�ߏ+Uh�wo��WX�h9����7� ���#�}�j�e�˭]�{���&SD5����w^�|�E��8?|��*x���ν�\����od�ԃ��9
L�{�(3�6<8�,�go� e�6MUNׄ����Z�[`
}]�q{�I��[��Y��d�_F.�R�H{��=�����à%����y2��S�}+���7O�A//��MH��;*�j�:�����1��֙˗��&յl��|��s�9[P/�+���Ľ�J���WhyT����#-��M���W�60������o�2d� ���O��ai qb"m�-Bh�i�FAOU=I���#�>l�8�n�Q:Ey~=~q�����Hhƕ�;My��E�jPr	�n��@[��G�!��	�È�� �Tk/� .Y�z (Y��׿�;�C���=��
��_�� ԗ�=
�Т����O��J�ƫ�˗����7˱��YB>���д�=bTحʟ:��K���I�=Z�@���!7ctJ,��]����}�zd�s�[�+(��_�Y�l��r�&.�U���j� ��<���t�ؽ&dSNۑ?iK�֗�.[� ~p�?�y�2�L2��݈�����a�z;iWod	��@�hW!2�PTL͸�܃�nO�BncqVm���_������`��<�]�^A���W��.B��e�Ѵ��ӿ���:��!zA`����KG�e� �H��mծgɀa��t�~N|#��d���6�̊a���H���������%��/^O�U�Z@���,hk����J�)	�Lǭ�������҄��M�r�������C#��6��&4o���A$^�݇Ja����b�Mʤ���F�ZK�����|Γ��W���y4���;H��n����F�H���h�7�����L;%����o��a���(��%�]��n��Cvo���&w�|�U)F�t.?H��xAY�P��:xC�4ʂ�������#�d}�}�qC)[gLhH��~�l��Sy�#mѿ� D����7n����0��x���V3B��n)�
�ZT�Wut�#�Ln������!�:D����2b$z���̝"�����(h-���e��C$dʋ�m��%��)��*A~_�a�=����,ů�BAB6C���C���Ar����Ms�g��j9Sf��Co@��ߠ�~�bФ�31'2e{�	�5]D�o��:�XS�Gd.�%l
n���b�/�(�)�p~������o2���w\v���d��z �BAj�f�X!$(T;L�$PiZW�!���}��X�����j������ �(㋷[=
�e�����?x�{A�굥�t ��v�?=*O�Kwԛ�Q���O����G/f�;۷_J�tX��}pEe[����.+�
R�+k��K#�"��Ů��f��Ǡ���lb�2"s�1�>����J����o�^-כ�
�� ��C#i@�-+�|y��j�0���a9T��oo;���k�&Ísy�������x�π�[����E�ub��X��ߑ��Ĺ����X�STկ�AZxi�R�%���N�/�A���[��6t�>��E{O����m����J}��?���*:H�\(*�$5q���) ��-
:xC��n�'��Q�C�X�^�3�1��F=��y/�0�ߕF��㐅+H� ʺ���7�4֜j�.��\U����DռY�t�G]� oDX�g|���RA�092bG'����|�C�)�t��ݮG��)����X>p	\?�5�[�>p-�KC��?"�`��]��?,��S�u�Ȏ^S2~g�J.Lbi-Y����.מ�h��?�6&L)M�"~	3�
ņ�G�(��Ɋ�V�gK��� ��n�W��b�!o��0��ٺx���G��[T~'�0���b�x��9�����rA°T�W��>�~ShX�=��`���.�-x���1�{�Iց�c���N R�e�k~
tw��@���֓VTF�	^�=��ʾ�5H� ��+@[��7~�ܙOe�p��k�o�J��;�����l�]�	���&��h9��)f�|>o'iƫ���k�v_�m�hF��u@*� ����92�My��M�54�	rd�;�X�j�7Y�=��[+Hڽ���b�[0Bh ���4�̽�:��':�F��H��(t�\z��N����c)�
���7���\�(�K���%��m\1ۛv2�����0$����pX
��o;I��²���S&�/�Z-��Ui�
����o��{C�˕�N�ޙ�Yu��׳�
�� �hǓ;Dp�z�P�N���J�1�ϫb{����F��a��-��#T��`���v&�xL�"*�r&��M� �����3aX6q��׈���]D�w�r$���A�������D���Y1����9��w�(�JƂr֡q��R��(g��KѬ��qQ8�3�P���k(c�D(��ǝ=�p<-:̲���<�n� a�^��a�*]Tk�Q�E��y�� p��fZt�U��0}�J����	z#��Xz*�jm� wC��� �īQm���X���D�1���j�g�p�� SV.���ڄ�\��]�7�r0�������@���nk�n���NA�0���F�4	'�+n	c�H�i�l���玾e�E+���:<�������s�����a�G�@u���UB��kl��H}���s��#��,_����ȑC��}��zT�hHہ)�����<R��3��W���5tZ�`%��:���d�BZ��?�B�s�ܹ��AxC���#(\	�;�oii��e�r_��!��� ��7GF&�}F�Ѯ��CX�FJ�{[0\��Ȅ�=v/�s��/ ��p�)�#H;�]��ޤ��wΣkH@��v[�txI�-�H�����v�ܾ����i˖g�r⏗�&��t������n<���Oy�����R&�4[�vL���bXg�-��M��ӧ�7���sp��e�O�s�������˦c
����z�<�����KnX���3��e�B�m˺��k�M�X=�;T�]��`�_��T�\����u�#௤V��6�N������|�U̧S�_'�����-�vdN��02���AcGY[+3��6�Gt�/��6�UtЪ��ͫG��p�������>��!�X��Jx�tr�F

���ￋ�"�@�rvy�߱�h��k*���0����ڙqw�T��$��x��TCI2>�2�!���#�
RL��ty��by�I�z��d�@}�&�|1s��~h���9�I;P�U�m_1�є[C��d�T�U��A�1<'v;�1��GX��pPՕ��qT2:%�|��c��&h��::�k3��ww��V���_��<~c�.�G�SKW�TP����p��89HP�tc�9�:����ok���C��5��,p��#�
2}1�wT�|��x�n�P��y6�b;���g8��m�J�NA�7���^"6�
ѧƛs����@�$�b���BT���=���}����T�G��i��ʏ�`M�ˀ|0�1_\�s�a�Ls�{ V7����BR懚qKH�_��o30���:VS.��9��b�%n1֭�� �x�(��4r�-��9W���S���ڢ
A�g5��o��NA��y��Ѓ����*���M8fA�y��<v4�����`�z�b�w���<2�sA��`Y����0�342?$�gI]U�7ffO��X�����+��48��/�bp��C��3`d܍)��p9�VDH��rߐ}��^Sn��q�@�;j��^)I)/�]�{و�������L��iϣ����@�=�L�{���)H�d�T���-W��������T,!1�D2���(��u�o��cs{���!˗d���e��V����l����M.e��-e)��,��5جK�l�2㣝�$�e����r*\�s��)��m�M奄g�+�#o�P�w4%�(�p�w6��t���`���0��k:�^��O�:���!K�~ɝ�
��U��e)y�sM�n2)K ��R�ʧ?���Wv�r��wI���n�l�����;fg�*N�&�dSb�~)�9�}.��x�����{ц˝P�o�S�v_D��с��O��sq�xbr�[�]�iV�ɻ�� @��D�(�c`�T�*_�ǩq4�����占��g��T�n��A�Ԕ�G�d��O�,���1�0���Pl}�2��R7r<�)c�YX��$��#��W�sV���:��i��@56����A��z�'�b� b}Hk}[�י��=�˨�r�+w|i�[�]�=�'t���65Ux��ŉܚ�Ҽr'ں?�PT]��8=����<i�G|�������(��=/�}�r�I����w�t�b�8=�*�P*jWg����TW�m-s�W�Ao���z$c�ЋT>[�Mb���-j&�8OwF�p
M�q�/�A�r�˲i�y9e��w����i9�$<��M����#��dPZ�R�%��a.����	��_G�7^;��*VIsE ��d�Wh��ަT����}4dP���GZ�����4��9-i/�M�������qA1���'�.�a��^+o���'�Y|��5�a;?�O�}�`���.>���w�>�Y���542���J߶��$n�	ٲ�����ٝ/�[����yT��^��.?��]���j��ϗ�G7��n���z��lXt4.y�B���q�;�};ͅ,$���"!!!�ȡ���Ȟt�AT��g��"���;3d�|W�������@{[�����p8��aW�b�,QG��G�/!r�@�$U�/O��(�,g>��g�a���k"��+ �Sab`�X%�Rc�>��s�����,4$lf��S�*�߿?��p��� �Y�6��*F�#��!m�8�"Nڪ�w�S#m�d�I[�r�LBN�gȀ��h4u{�U��{��y<�����eB{��iF7�5Qg�ZE>G�r�~
��k�y`��fyBr�q'�,�mٯ?������3}��M|�:۰E���"(=?$�4�=3�HPV0��������HuЅs��Z�߾�D��H����LO|pK�����)k�Z5t��$�*z����Cf���M�R!E��b�=e%���B�v�d�ko%/cXtI���$��`��hq�����w{��Q��Z|z��U���͏�p�Fb?6:��$�}�v�ݕs)仃˴�{H|*nU{ښ���;y�Z� M��N�u�Gt���������א�݈��.|.K2
�� å�JCy6��l%��l�e��uԿtV�Om��c�y�ߚ��G������^Y���HY���p���r���72/����s#6�p?�`p�����-`����b
�R�vG@g���3�[���l���jq�7O3r��P>������#.P���,\�T��u��g���������t�>�go�'�>W�r���Gv,>W����`�5����[��+�;��-��h�0���������/B�o������D�&=P���t#(Q�K�Z��.��hco������_ڹh��'���V��&��ĉ�X{	��[5��$1���Pp̭Y��m��6?��Q���C���ټ�O ����7�&JD*o�$י{����y�Q��t_i ����SӁ+�Iy���f��V�����j牷�N��Y�X�S4���-�{b������E	��I����-�Bs�pe�����Ox6oK��'G�a64��p3��ehf<y��!hވ�;cf��쏚0�M-���p�O%���J�bĨ������.{ �L�F�2��2���J�/#d����ǖ�ԁ�~�>�!"15r�%���l����Y���jio`�lu�[F߄|�}8	���V���7��-41m�ބ`�E�|��%������d[�'���u�0%i�Z�qv��[��!R�l�ļyn4�(-a�\};ܚP��$�V����P���	�V�9��xY���
kj���Aj}�$����(�h�TcP�l��`���{A��~_�Piخ�1�x���0���5\r�j��	��P)�#����w�\s�B7Gw0�3|y��-߫h�Rp����G�9�"�ց�Q�9��^i	(�2�>�Bk���k�K�T�V���8+�nQ��Y�;$�3z�n�E�w����v�Z�'	1�k�K&��%Ary�+F̠���adV{��_`?�&Q�?g��L5|��ҍ�2�Z�Ƈq�ԊUj��
������:D������L�!��{�v��UVl\���&׊�o��#YF����*3_��w�X�v�c��|"5����+����s*���t6�^��7�����5=�#Y]����	�j�n2�eQ��O�����DO[�ֿ�t�_ U$�﫨�lF����0\�/��$��Z-�{d�+��tJ~��r�o��c���b��uGg� 3� 
�6�Ad�+��0�+���S�0�߃���4{�����q�a8�A�m��/�D��ӷ�T%�	<��O��sf|/�{*H��K��[���[���M02^]C�+�<���q�^�)Da�s`�%q�z�7�
��N�fG�t�`HL����Q o�`���C;�Wz֐1%;��ε�쩂�7���S���h2F���+��%K��z���*~Z�i��R�s�L���#HBlU���j����2 ��И�� �Ta���I���]|:�?���s���+���Z{&�5u��yC#�� A�u�p)�ii2�-��&
{ƌ��ş�Z>@�J�4��[�vs�ć��@y y��������K4wU��->C� ��O	z����bޠ~GI�1�kN��S���\�����Q��5f_����2��ꮬ<�&�rq�Q��|\�|6�㍓銎-ti/,�����w�j�?S��q-�]��<�D��j�v�	�cl�%��WG���"��z�5�����O�Az �L�y@�.���dYG��V�̞F�G�8����W���y������^dZ�=��t�F�w*h\���k*��u��ݠK���g�a?���8�y���Ss��8��rͦ3�J�yMV�����-�4�B�ڦ�'�|4�b�e����m�NA�+����@Y�v����i�g�Vʝ��P+�E�]U���Wéuq"v
�Z�cg�F?��TM�-;\ը��-�l�#Y�l�?���S�&R�
���ӿ��;0���p(%;|y>���Q\���I��6޵(EȲ�(R�N��r��d��JM�6�l��cJi�!hkJ�-|�1�PJ��<b��e�����p�����}%
oƩ]	Yۆ�RqϳcJ��Ɂ=p��F<t��t?�Z>�V�}_�F��}J|�n� ʙK�8*J���y�o�t����;0P�sp���lGG�<���B�@��l�՟�2gr{�Aͷ�0p�)��G��zY�c�
O�+����'0�a��X�m ؿ�`	�E�M�y�s��apHs�c�*&��]S��')Z�@������!��0.�	���ٝ�=��u,Ͳ�����oZ{3�P(�~����T}��m�,b�VxDa�ʇ�_?%�x9 �̴"o'�J�룵�[+SQ�{H�$�������D:|���<�!�C�Цu{��Y$g]�ux'g���c4�(ݐ�M,�y�+������
��h �0��+)��弚�U�����$t��G���aJ`�<,����>���'�e?�rp��"�΃��yQ���x�ܐ���)�Lݣ��kU��\�c�r�?��.w���4�\�:��p���@�P�8�9f(D8��[M��q7��yt�.����{M��Z�=��p�8\%��D��vN�ߐ�o�T�.��)Hy�NZ�ia�$�o͂6�L7���)�=�35����fDx��0��-���w��@����Y����?�޴`���GZ7�zL���7��3p�Hcj�Ӥ��r�rg�� ���� yhꞰs���D��<G~��[J�`%�>n�:E��ѾB���ɟ�y�x�(�*Y�tf#7[1���ע;YZM���4Y�AMe ��D�����2�7j����H����Y�y5:Z����}6:��s4��-m�ؙf(��z-;�輋b��H[q �Ƞ�|Й��~
Rƿ8b�����+�O�[d
Z�e�מ���
��a��E:#0�o������˦`���`�����!L/��J(FyH��� d 'z�~��l�9b_T������P�2��
�`8Mjo�m."]�5�|�LP���U��E��	X������h���:�c�%k��Z�X}��xV����M��i\��
G.sO�Y9����z���l	�s�.�.���;��5@gyi,�2��;Z������7��gy,x;�%~�4��1����/+�y�0��ZQr�߲�D�#�&�c��yؔsG�)����tQ���gM����N�a{��-�M���m|����l�%Jd¹�(d85"O�ﭝ�Y�-�qRi8o昼��4َ�Ⱦ���3�~
�`��n�W�q,i۟��T��GV�5o��Y�U��g�Ͷ%�u1B��գ�����5?�k��ꪛ�C$1��PDh��8'wH��Dچӕ��|��o��K����=�z�W��C�J�:~�TsZx6^����?F����k������;|	��=
?+�h|�s��Y�Ӄ���C߹�vtL}�=y@?
��@��]��gW��]o���s�)�^m���o�B4:}o9Ϸ'����{ʉ��+�y"Tt�:��)(de�~yU�D�vͯJ�y
�L>����<��d�AU��sh�0���[\��#�E4A��s���� %Y�+�ҊN4�3/K!.X$yBj�l� ?t��̷�l�ڌ����6e4�#Hv�
�S�Vb~,����E2l�j�֨<)���k}p{ˌ��+z<ےb��Q�ه˛J��{ʋ�=�!3I�Ѣ��=�<��Wpm+��p�~�_yQ�ٱ'�/�W�y:'c�nj1�n7+nH�3�v�l����}OI}�s�7?��i3C�jr����St�)7�J܂�ɭO�@�W`�cw�����V(zq>)k;�m�dq�ݩ��6f�qw��N����T�x�p�,?������#H
��S�a?��:¥�Y*r�-Wd1��nW�X ǝ�r<J�����6�����ZK�sr�p<�W�Qܹ�ul��fC�MKz�AA����[�X�τ�����a��}��ן�zW9Z)n%?���n�wN�~\��9�����7���S�6U�&έ�)�Jh�����1��.&�'�6�Y6��&�ff�o�`L ���E��Qjǀ���֚F85~o�0�]�#��w*����Е�Q A��+�%$���ww
�kJH���Җ<g�0;�����gp-vۺ-��6�bh�vt��o�smK[�����:#�FG�-ѧ�_#��NXS�"�����~��!�l��1�荩��3�$Ų`��*},�>��ڋ�ҩ������ku��:� ٹ��Ǳ2Ti����d.�"kYX)3Zh������5m�5����g��O���<.d/.�:K��A��n���b`��~����OuW�x���:�'��=/��7��g]�!"�6�Z�������ꐆ�Wީ��~~\���(@O IAݾ|X@���T�D
���4���A�g���mꚇҧ ����/��A,YZ�v�E���,U=k,��R�>� ���8*m@?�X-�[���z���u����~��~?�hͻJh-
Dp�e{�x��M�GLM���+��GP��9��
��ڃ�>E�9x �v|���xTݒ����;�!�)���N&8��^\��{=V�5N����ߑ��-h�U�UpNI9��h���q$��=�������]>,o>0�}�*�uI'�&�jH���g��n��s�˯�ԻWF�d�Z��F�+ʡ��eH�pX2�W�τK*HQXh~f,8�/@��2���A�(�ӗŷ|���^��3c�1�H��rS�%�n��rF���
t�(?�L>�Y�~s0��\En5~���k���1�yіH �a�T^�4]!! ~�6��/l�:?H-����W*!@!���Z4PO  ��IDAT4��b��>�,ה0�4"��������%ݟߣj��J~��5���򹉤Ƙ3���t�_�\��{#�!$e�f3�ȳ�V�x�N���mD;���ڃ��n��{_Gz�H�Ih�UŴ$�I17y��_��^i"AԞ������$�jw�B
��t���w�Gf\z:�ب����q(�6~m޿$-�z��{;����Ԏ���$���MdD-���8�j����u��e��e-Z���orH�C����;�J�3Bl�-Y�%����˘QΐM l�)İ�^|T�۶�J-i{�F�W��gu7}'����6D�lJ(ҭ�ʁ�a��@Əz7)f��X]�����q�ŕJ�5���w���f�r^Z�F�B�8˕Ʃ���B���qJ1���l�"�][wVq�����q:�D���S�V��6�ҩ��yu��6D��@}	Ê�(M��ae'Fa��h� �B0F��6jQ��(A��^�}�ot x.|���w����~�>`���\�;� �>�j�?,Y�$)��Y�pQ	ՠ-1�g��-�j+�XF��$���1C�V��}AUC��
4щk�t�\����Д�;��������G
�!�`_Ȕ�ǿb��氊�#nj(��Y��׿w !�CW���+ia�X�k+q?ʿ�b*��T�;~(�¬-w�)J�;�N
#=זRϰ9�7��n�����X �4�l�ou3l>W���v�z�̶������׬������#�BhY�W|@����(���m���Z�~�#�y���o�9�&�6W:��:{�� ����u.���ߐ�k6�7S4I�c�&[ �P0�'�v$�,�Q=���`?p�>�S��^�͛����A���)���Q�A9)8b
��/� ���ܹs}����h��沏�#��z��g����-�b���ܗ�a�i}�+6W���&5h#Ӛ ��XW엷<�"F�)^��9���Kbw�g`o{Š|8�[��n*z��b�>T�k�¥<&LĕpAQ�9�u8���&cxBŉ�.�kM������^]N��k}�����Q3�S��:i��I�W�B(�����-nm\�Ͻ5~mw�U��(JA���u�^+�{ �!%D�S��tj��.�me;�74�L�9FY�k;��uxC�~�A�+E��-/��r�X�W�C
^W�
�T�.Jz]|+H }�/�?U��l8[p�b:D_S+��Sb��{���&��Ը<���˿FJؔ���!�����ƦV�b�ez:}pg
,�e
�(���*���NS�SU~9����e�w��s梱�����̵�=k��~����}#�L{�V��j�(ҥ*S��&%d�K$�Bj�f"��=��1��L�4)� ���/��t��<ީb�	�����T(���M<�n�U*�N�9\[��g:����t-Qv%t���S���:��>�aa4 ����5l��	]2��Ҿ�E/����=aW��5q:���ts��ƴ�����ـ����T;)�&_1c�Z���>5�vmԻ$V��O���&.�2ne]��!��4����=�M9v'�������.X������)]�ǡ����������\�u7\TA��� �і����g�5�ds��qb�t���R��VGˑvb>q�"ԃ�ʏ��b9���VWU�����"�}��R�B��=��@y1�iB�P�);� G��Vvk�jx��[-r0_rMԇ��R�x�5~iK�?֜�
�\�
�����ۜ����hMF��MQ,��Z��	©��)%|C�+vkUu�4o�����t��v��5��3�C۠�~P��oB��9�6�����hڠ+O��M�� 6����O,�.)<��G��g(%{ `Z��V���l4ib��S���>D�PE$]]E��(P�4ΦPYP�74`D��V�v�(�ibbzT���Q��#����� Ȍ�k����nZ�{��O��W�H��jNu���Q������^(��dr�����(ɑ�*+�%��)�0�lo��%���5+XB�}�)L�_�)�$T��}�"�cly����a eV���7J���4��h�S}w���AQ�r&?+)%��:Q����(�w��^�gڄ��mP��k4��e�`�c�nu��y�D\>��,w�!J� �]=-��鸺`���JM���ѷF���`«:�Vգ���Y���S%i	��ӭ�a��j��0��t��cS�Ȣ��OA�Ǻx#Mی\�G/���0d��.��<�\y��U�C��˳)ɺf�U3kD@�n�ѹ�����);�6#-�Ƹg��
�� ����͢b*4c�����1nw�gbF�/�1�����Q�T]^�A���"5M�@�` 
N�w���� �̔R(��΁j�Q���FSQ��x2��똫�cB���{�;A6�ea��6��h ���	R�Q����A�Aq�D�	��8�ι�J�K��1��z�f�@��[B��☰��ny�70��Gz�s�"�
O��ĵ���q�;|��Lye��#�m2?`�i�c��[�>��\#���&О�:�P�{����`"���Of�
ZL��G�������W�\OA�?����K�fa��(塬���L�,�O]��b͢��*DIcR5�d&~��S0�l71�d�UJw��h�� C��J.
{��suQI�=s?�������@������k�qJ�^��k��'�������%ۭw��<C���~O�sN?~RR�0���J�I�g�������G�q'3XCӯ�5.��m!���ۛd��T�¦*�am�"�.\q��!L��R��GV�Y(�C܈.�.t�P/`98f�)����:d�vwB9�����=��!�NZ���?�0�(�����\*��q�pv�G�4 �<#����<�F��� 1��K\	��
9�P�v���;V���G^� �H�o���_��1��,-B�Z����F@�=���cMWvA#�����
�!c��ǘ�z���?��Bt�4�E0����$�+.�q_F���y@���
��R�<��Q���w��:#&Ã�|L�J��x��C!����>��a������L�׏��!y�1_R
�hzGM�k�߈����_�$W�)Y���i%z=��_ҿ�#M���Cv��� Ӳ�M/� Kk$�`7��2ڣSq���*�zJ�y!0��Ƌ�皘�W$r�,��b0(���s]���_ӧ�z
��{����O�(K^h�$˓xj�	�G�+�l���6Y�a2#��в9X��I`�ؖ��fT�}k�ܗZ�	�����nv�h��u~0��!h��M�����~���$����"���z҆-�=e����W}vh�ה�	eWn�����������_����,du�����&��4-g�'���%LA߱�"T���w�"�6E�l1Aq���Rc���L��������=�ǿ����CA�#ݧʘ\ŭ��L���j��V[ ���[
��?�cMD����xH\�o?����%�1>�:�&��s��X�nA�H����]R��ߌD8q���b�b\!ަ�E�^���f
�i(��B��s/��=�J��i�����~�����}�9^���߫��3}��Oc��R��ñ��*N�}DV]�C`���T�c����4��M�����߳�t��XAz���9�v�*��(H����%��Z�1��u��t���U�Tu�P��\������w�	\#�+dK�h��e!N��%�oI��������ӯ���uo@
�M�k`t�R��ě#�m֔�1ӿ�J����d��B�6�,�0+B�������]��&%<-t�ђ�nV�h�Ɛ�k�������w����T.v�[�
Hؘ�\�ob�n�o�@��$/-Z~�����=��)Hˢ�ǯ�P��&�hّ�]cMX ��B��q'N6V��@�[GA���Ҟ�����*��Xۯ���!��_�*�ڶ���#7���g~(��JQ�"cƝ�Ch��hu{0��_$��L����Ep"��E�\�˘�����<I�(�tAK�k�2uMz���s<�#��\��j�Yg�_\�*S,B�_~%��!��|В�����R����u��+��S���Ĩ�M���^�t.�Q���\�ʚ+\hɷX�<����� ,�n��-r ���}Fh$uMum̎��Ż�<ڠ�1 ')3���C�r�Q7�X梨�*o+�=��L���tO?��1~����[�D�a=Ck�^4������n�J3��}���h���A:��چQ <A�ݣ����2�h�_�x�����B��if�L����Ί�w��q�k��9���e���(g`ǝ�k��s�nE&-<�ZR��_D/��\�.v�k1 ������2v��L;؝�H�N���@�a�V���:��N��9;h.d!Ӑ�*��-���c��g��Q}�]_����{���MtF�����A���
��*�A�&:�))�\��|P����W�# s�-��|a�	S�Q��){�|
�� -D�Ǐ�8Ayq���%A��@r��R�4t��}�t��t1��<e_i�R����2׿�V��݇k,~G'�u�%���Kr�	����H��-2���l�\�t�D�H�t7B�Қ5{2�j�φW�
F�k^�H�X�dq9+�If.k��_Qm3_Z��@ї��š���{\�S?E����=���z�m�Fk*c43�+�Ҝ)+�˹,��X��y��G���7�M�-z0#fWDܭa�̍)c{���nq�[�;`Q�ss&Z.% ��w4�oVt��2od�ם�>���^Ǆ�r�P`�\�v�� �����C2��I�;V�7���@�Թ�d��` HcD�����
"��SZ]\M]���Qp�]�RIK�3����!�/��m.�E٫Zm5��"��$\�^ebұNc8���b���3���@S��l��"���$̫*B\,�Z��x-�go,�(�)�NT���J�,�dǠ�'�˓��k7&|��h��,����7Ӹgű�e6��H�<eR�1;~���^G�fA+[f�U�zc�S�!�����R�<z�&5\��2QY���Z��;ؐ_��ȁ�Mp=)b<W}�	�$_��R%�@ؐ�Lj���u�� _o�q+SVԡ�2��JAuM�K��+]����I�=(7�6�,�H�o��-��c���L耄l���f;ƶ��zi�D���1ʠ��\��`Q��SJd`"�@����@w�����A�l*+ #��Ʋ�@�\��ߵ�04�fc��V�";LQvaDp+��$.��r���[Y��Mi�q��ꎂc!��h�B4�1�$�Ն�D��s@�(�FaU��1�qp���n�ǟ�|�+[él��niVi}+�9�t��Ѱ���6����)�����q�Ќ��"Y�a�߁�گ���̹v/�vg,kp�����1Ns]S�E6���EQ���jp42�Y�R��>7YD��>_k���5�U�\�-_%�N5��r���{��a�,�hԜ�E��>o�׹ø&Gwt.�4��|�� hƂ~���b]=��TJ5���r�Ӝ~-׷[vS�1�.0�3�ͦ�7I&��$�!8�Oט��=*�\��c��� r(�c�'��,�^�����^��'�^��Q�+M�z��8.�v�P~�B���\2_%��E�cW֔؝�$��$�%�2$s%�B��3���<IՃ*�[i��(;47�B��T�oӗw�6�&,P�1v�bC���HD�=�Ft3$�L��e�����Y��$��=i۝��C����nBԖ��f*빪�:���]��%""�QH�A�������Z@Oc����bTG�=SD�B�7�E^�oФZ[0��E2��#e"�Ф��
@�=��p�pǼhl��[�J[��D�U1,�y�NМd�a5��i�%v�k�Ȯ�~7���Ԍ�:�ܦ$C�+�"�c0&����N$�/���򓲾H�G2Fi�$�A���a?�P: Q��F�PL̥
�Of:K�i� 2��M�5� Ub��@�wk7�������W�*��f��j�r	�G<׼i]����������h@G��^��k=��Ѳg9�k��Ǹ��u#}�]��$�q	Q�N�4C>('�zV�*�A�D�RK7��i�Z��O/�Fp|CZ:�^�K��@r��WT�-r	=��b�;1��{(ㄪ��3�J'|�\RA����r��i^Et��z%�k���4��%�ʐF�^�-�rZ�X�}P�Sa�=Q}ٲ��|�xT^~U�9W.��B�K�,N����d��J���P�7	��#b��\|�K�'0�O�@yPT��z�����e�:O�v�D6#��}Z��E ��Bu���+��8b�)�h
�g������Z��~<�����OWY��$��,�	�4�s\9\5	W`w	���j�첡\a؊<jS��$�X�g����m�7M�9�Yx��2���,��
XX�i��Bꮜ%wJ����@��+-��w��5c�5�j�n�JS�\(�R�Ր��%d��������}���Y�rb�	� ��ҫ$H���HC<C�r#D����������&�~�dw7(F�9�@�/VԪ�*�E��@+D���6����_���Β�%�tNM�E/���o>�FsD��:���sⳜZ&�e�/���h�<�u�����Ѣ����F���,�ˋ=�&<��?K\������9�$�e�&h_Ʈ4���G7�B���Ԥ��^��g�ޥ~��o9U��5�(�B�_ǋ��:C����
�YW�d���m~�!ˑ��%�<%�l�φ`г�h�*���0���/.5	�a�Ze�����σMAF�30���#7;��L������u�B���V��FLT;�2�z�H�J�<��uk������Z���5���Q�-�� �~��t�P��5�D-�#��b�=�X���z��̬�����
nQ�ړ��S�%�+��Z�v�E�\�VH.��@�ړ5M^/�>MU�KTv�Asz��BN�BcYO튂&t$g�~B�����a�gpJ�*��m؝I����%

��<5Rm[�Kur�Z梏�`���l��`�Y����wl�����,H�e,�c����~�1c����gz=5��Xp����%ڍ1GO��A��l��@?�U���
y�ߛ��М�R�&�{mA�iO��rX�����/�ޞ�&�.���G$S�%�aT���`�(�]B�)��]/:Z���)Ҙ����h��?��̫Ԑ.� ��o�=Cd�yAe`��݌�w�Z�s�ua .n��3T��J��� >Ҝ鱇J�C���*��7�ͼ~]�x�Y�I@_�;$����(3�����X�HM�p�Q�P�k$$Ǡ�����8&b�}�� em֌��^��	������E��`4�N�̖�K���?MD�3�A1�}[> ��)N�T�JVS���@�W}9#�হ���ucx��k_>H5)V�\��-��n��&.��8��alG�X�v��qB4f�KI�ث���ɺLN�Չ��2�>�s=����P��ʛR��1n�&��eY��P������Zi�ҕ�e3}z2q/C
��/�s=\SAR[��
R��$O�P(V����w��0h&ϖ�2إ@ \;@/^B�M�ͧi�6�a���@�\��`r.P��X�%b�W�<g��E	���ϛ�����j�sn/��,1�^��MV��|i�28��Dr}�ݷ�*HQSL�	�ɖ�3�#��bԍ^�L��0�Г�O��ϏG*h͂�X��ٛ�mѮ�;��(]�:�9�Gs�.�zE���(�mE.�v� ʗ۠ܗ����۶q�נ �0�^#Gu��O����s;;�#�=R�:X�`k%�~���D}%AW�+�`�ʹʡ0��x����긟�o����j�NC��J]��W�5G�8^�Z?�!��)v=A ?�t�#����7�YI���)H��*��CM^����+�+\�/U��(��y�N�N��Tq���Y��()��h��B��!eDf{m���L/�:��]�g���M�C���?T�`��_�N���>K���q�L��*��J�>��h�N+�پ�L���}cS���= P"�������M����hXa5a[]/�9�r� �x��E�b�Ο�M�3	'�����k�U뷅-��.�Z�xU�H�H?��+��<O�B���V�C��ZCcp(��]����)r���!w��M�7*c{qj��ٖk�A�eTd�}���F~a���[��<q�v��۸�F�3_V1����zv=�tzS~�8j/5��JfLm�=��L���~�+�=gc����P6�|9�H$iaQ� IvO��|�����)��B3�Up���25bR_J:��'�C��������Ȋ�������F������Q��#,W�K�KI_ %^+��-��\�z���e60��q'k;)�j��]}�E��#52�^�������)�Q��i<iΰ�k>�SNR]���]��5��{ R���
)ER�^R8i��Ul����c��I�8a��
��Ɖß7u�"U����$����n�%�6��"B)��LLo�*����:!/��!l�Iڶ󴥁ʄ��V�B
T���H�c?g��oGU��Ou��g3�ֆG'��A1Hې/RPTyhߦ�����f\Q�ٵIj�p=��̟�e>���!Q�:��W��?/�Mд#��Ӽs0#���%H5x�=U����+j��*�г�l��ǐ[:���e��6#��>���� bb�tV��F��hߡ��.��&!͕�|
dQ��n�����ȷ)�ŇT�{��G[��_tO!˷���M�zc�Q�-0�]�(n�D�1}h�R��+�MOz0<�T�,̏�>��%�=��8b�x��rg��MöL�Z��E/�мg	F�Ӯ���Qc6xꀡ�-�����F�C,_��̪���d�_�
g��#Bl�ZT�Nfd��Lp�--��g��K#*5���6��^���]�()塰�v||��Ki!ig����s��ګT���F)�xTƎ��Ua�(�"X�ѫ"��m?RP9uN��?��2Ft!d*�CG჆Z�v�pm?�0l �r��	St�Gۜ1ɾ�k�&Fbl�8 MyO�nI�YV<��\k)�����%��
=S���2v��Aq�٧���e���,^!���[$�ڒ�7�N�Pe�0�Z��S����HXG�z
R/���k�P-"S�a��A\�S�Y�:H>�޵�~U���B����� �C�H��
6?Y������y�4Dt���� mũ�If��<S9򂈾���
2|�lI�V7QL��9�u=0~�İ�޻�����o��Yp���s�l�E~	��vuN>ˇlٽ\�%��u��e^I����ײ'Y������NWx9P�OD� u�\ڰS��w���V� �}��oɞ�!#�����j��~���Vb�>1���q�ֽ�}�"#�"ߊ���%��S�q�l&*����El*��гX�gK����$DP"���(
_�� s�}��4+�:9v ���j���iM�n�n�V���F���o�Zm;+�`�k��g��i]U���DBK������)<�}�ޠ�1��7�"�@��K:�Q������w(��N������<W��˯�T��Y��=ؐ��t#�X�=BO�ٺb�a/��l��or%
�SH�ZT_��=���]p*s��+���iڍ����6M�j�i��)��Sئ�kq[b��C��m�U`���׳bh��,j��R!Ry@�uE�o��I��և�Y��.����~xQ��5̗��5���Tݤmc�d������q��'������$yZ[
SUNL��m��J����~�
p<�Ӂp�sQe\Pj��
���h3`����Ds1�
|��Z�j �|N[`T~��J �����%;�L����;��Y��.s���q��7��-[�V��Ͻ!�6���16}�uxӹ��?$�*�Q��O^dMi���\�"��Z{�O�\w�j<��Cؾ�ig\�Uxd�W8�z_�W��4f)��.�-�2���`��{n�ޮ-�5�Z3�ޱ�7�EOݔ�#d�k�B����{�,�?�(����f%�ja8�fy�����$�����D^5Ç&L��pM����4��)��4$�a*��'^b�F4<��"���
}�)�[�r~͏�2Vb{	���G´��o��d�w��$��#�`L_>�m������MgD���A�����l�[B|�+�Aj�G�����ߚ���r�婝���/� w��LF�Ĩ�<���E�Y����|t�,�%�=�n����v7P�l?������n>�=�AN�������?��b�)A}1Կ�f±аE���bW�ǻ=]#���(�˟�[�SN�:�K,��p�������wvk��py�7�#�p6��d����{�rH��j>D�̕��Qw�ֱ'�s� ix[��ٽ|��Sˇ��<���Iu�5������Q�I�JUI�䌉����|RVE��t?h�餰��b��ոD�DE��l!gs;7#غ�����n�+�~�zk�ܻD�-��Z��y�9O���)H��<��,Κ���"b欅<����v
�h�	�G��>"}:7���@E4ru�J����I���v�B KF/����F�h)�B�'2X�$?��%�砖�ԤH�ڢ����-�s��(X����D�|���?ò]@A���w~,0�guT)�����r��|�QQ�'M����^��T#��WA4ͷ�NJ/D��ٍL�G��tX!y������u<�{譏��%Kծv4g����&m �k.&JU�-֟��Pg_�˴���
�\�T���{�,�g����)5�>{����LOQc�1��DK}�ʗ3�8F�(�r����#p=s�e�[�W���=M�υ�5�Mq*�&�XV)���n	iw�g$�R��&6z(�P�#�P�9�J��`�����sX�|eQ�u�܆�ڙ$$NR�|�Q�u8�N�/�\�{t)���H�t}=��V:唗�J�F�$%�K[����]y�֏�L�^�g��r
�wz�ˋ��i2�e���X��|�����듩O�E
Ym�~�$��sݴ����cwG ���uT-�;�q-נ׀��� }�hlŸ@��2��_�^�/�^�_�,a~����aآ3v_�.1�[o�A2c�UE�݃e=%��"����S���7�è	I���:��浹"8�++���2hh^�7P��z����y�mw��|8������ny'k�S)꺉��tNކ��y1h ���SNS��=�P�����o����8Ш�
�)���$�K�剟�O�e�fQ�ґ�'��M��h�k�|���4#��ndU4�Z�{�ma��� V�n~#�vZ�ӿޡHoC'|ö��w��S��ƺ�oY/{A|#�)[��@�,�������PU6?�`PS�AD�B��4PD�iHsbec�qg���-���WtZrMa��h�ϵ�' ��n<��u����eX�n�:�~�r9>#	z���+S�ۂk
f�,�N�ʘ�8�n���~�Qإ�F�8��>�{��i�xx ��x������}o�kZDD7��ґ~O�}ޥ���Y�՟��*H���\X� G��g?�ny�b7�Հvԅ�1I�m�+\��k�m,���O$r��-c8�ߚ�S����m(�+�������(J[�$/�iv?���>Xf�gWY+��vY3�rU��ٵϚuUdFsBk���L	kc��飴�(+:WO?`=�H]�'�`d�<�����5�`�LM��f�0?Ң#bP�MS�������Ź��~C�T�>�dc	M;�ѫ�R��`<�Xmi�(�(\ӃJΞy�����
�� %X:�Z=�q�Oz&Ҍʊ}���zGBq���u)Mި�kc�g^�*�×S�6�:D{_aF����ǈ	��K�o�.���|V9B�AYq�\o�05�G�����F�*\e����ﯷ��e6x#2J����QK[�
Z�n�X�G��D
�@y	�tۢ��rf��z­������"-6�xq����;�[���?����ե�t%�x%i+`s�v�����Jo�F&Y��c�m�#�qM[+��:KޤwC㪮/�k���F6��Q8�T�zd��Kc�x1� �3�g�7?�p��g-Ğ��v��52�j���0��0�a��4�mTŭ�L6ϢX��D��_+���ǽ�څ�%Nzx<��|Aẵ�.}ϱ���#��i��D}�i��u槦���[���h�5�D�Ej�~���$^�$�=%�����C;�$��8�ڰd"��V�K�ˀ�n"��O�����ϐծ��k���՛}Ä��W��)H��T�4����<�5gXz�ѭn�ZXݓקEy��5����J;	�>R����&��p*L�����0�o#�'>��;u����y?��bXw��~�[�'zu��4�ނ�[�V���aI[��ㅨ�����]��?��D�us>P_��� �i�T�
b3��*�Tt��ޭ��K�dAV���4c��	e}8rn�=�V�)��s
�/�Zѳ[�BI��~�r����D���ryH�3ZG���;�E�9
C�%u�Q�2鬆ʚ��*�&S�E��s��X�����8��fT�N�;��c-��f
����e���kT/[���}J; ʌM�̌Y�}���<:�A�%Q©Os��M�ɼ���hw�z7��-rb���q_IGkE��"��D��3M��d��$\NA�W�����{w����C	J#`�e�C����
��=c��v�6��j�4%�����]�9����� �24�:\�C�Τ2����/E���Rz�8z��S�0"�?{��k��ɳ(�Vf�wi輈�u��ʖZ�"�o}��^;�����~�XwT/$��lRck׊.�5�<8�|u�:m9����w��$ ��D6�m��@�:���^]*�h�nZih8]D�Z�F�;�!���;�Y8ֶ2��5�9SC�\OA���F�=�B�P�F�8k�]�n_k��s�u2,�E6���v�(��u�i�r=��Fg����>>QȦZ-��5 ,i[K��)-h����IE?\;m�bLG`�Թ���wD)��c��H�`~X�v�M����͠�{;�?9}�l�C�$uWw���׺2u��٘!b�fKC�G�������g�W�{�7�{��m8��.v������\�쮍��$*?}����ZKTt��H����v��-���O�
��b��u�y�q�" �h#�C�y�X�z���_�$(�s��s���~c.i��z��n0⢩˚`&�'
y��(	����#�ER���RlIߜ��������u�G)�[n$�����%3O�$Fy��~�ƅ����6����9���\6j�	�x�i�΂�ǹW�3w�ϳ�o	��O���³��i�ph�(�qB�uBz^#WDtk�"�~��^�ښ�o1���,�#�,/) 튜�ԴG��_NA�tם5��7��[`�SU��J?ڷhק�(Kc�L�}z�1? �Q���������(ȃqCH�6*C%2?�oT�H+I�ϰ֟
;�;�f P��;k<���T^c�ªtk+fI�:�4Vv��mou�����@�\G����<�{�z�~�<���2��t�P��%)�hgq\e�N�O��y�Ycf}15J�?;�_OA:�v�صHm�YZ�ʑŃ������'��Z�F��6�藳��"�j�������^��9�Wl$e�vk�v�:��c����L��ַO�9�~s;���\HTdL�r����/6��Ca���Õ��CmY��,��Y.B�poZ��1aZ�<ɀ�_XV�y�r�ݙ��������7J�`�����
8rIi	�:tO`\��=��\o��F��5��#�����Ʌ��"}[~��V��{M�C���ŭ}������h&;��<f�Z���w���Gd�q�ÜG2���w<^>s���]1A׼�3q��_�]I$�"O��	�Y�/��{\v��Li�6���d�{�n�u��.��B���U��L�_ѵ�d^��pO7��hvu�8[Dޖ|�]�HZ��xk�[z�N�0RVJa�/y5�V��}z%e�:,C� Y�\�r����Q����2 �}g��[=�'�T�qJGB�o�'�OrKi�s<�%�/�]a�,Qʆ����t��3qiV�a��]�WA������s/=Rl :�{�"����\��׌��w�����d�Iľ(a���Eƽ�u$r�W����kCt�{gT�hq���@e��@����}H.P��-�Qt@���o�M��8�@
��]-���ѫ�	��R}Wa4�ޒ�j*��č[a�C�*	�/��E�Й8֖��`���yl���F��9>vt�T�O��Y������_��z�ՠ�����*�F?Ӭp�5�Hu`FIQߚ�j?d2�-4sKP�Y�z��v�mq���{��w�Mq�|ֈq"�~F&�Z���
��S����8�>�/� �Hk�X��)c� Y�w���r���zD����:�:��?|ן��eu��/ȴD{I����\�ģ�c�ex&@G9�Cض�<Q����E�J]K+�Tc�
���(���l`g���9��J��`$��5q�V?y�`�ml�w�V������6�*)}�1�g,z�7FAa��Op��K>����2_=�G��gwu���N����G�K�Z��V۾�5�9ZzI	�b�䞵�rhg]r{��ó�#����z�Z���+.	��u"'~w��!�3���>�w~��٭?��W�3n9�����.���g�Cm��a�n7E��i�f����U?����R������BXsE���'��퇰��hT t�l�@.��}N=�ky�0r�|%<+n)S���m��B�?)\RA:�����m���u!�������V/�C��~vQW�i$�b�{]�+�	gǢ���ҙ�z��Ka#-������⟙�5�nu�|(�r��
 �s���eU2)I��z��Vܼw��wi����7VI�Tۡu͆hg������{����ْ0���0�s�������{����V��	�h!}.� �.��2�sI�H�-p�,Ԗm��Ei�����X_ɱ�9��s/�O%�ً	;�>yԑ��:u6:Lw2�w���*C��g
��Ç�����+�m���C��ƿ����s���T�=k�'���Ϗw�}��xޫ�����q���J3���h����~dw���Q؟�t���;�w\�kCO���)���d�c�v�m\�]���4�#g���?:fP;&D351��&H-={��2�y��Sn�K��5b�E74�_�A�B�2��)�o�`�PT�kQ1��O0W,�kD�]�dt@���X���\lR%,�3��H�n�:$�Hptel;H/�gPrs�1��e��=2r�*�v&S�o}�,����ZD���WHQ�A��,��:��s.�"����tƲ|ͻq�V��
16�0\���7���i.D�����E�E�}��>�)��Y���u�}�Q9z=��1�W����ѳZp���j�\ᅵ�Y�C~DT��yԽ�S@|�E��T<�i�u�p=i�*�xK�ʫ!�ӯ�����y���K��EY:D��^j�!ɓN��Y�R$��<�Ze�Usc\�l{`�ȗ��N䀬����.^��SWX#���x���@��J�/g3��Ɍ���V�'Iۄk��Rә=[\#�(ru���߶xz�sI`�>9�3l��x\Ͳ
u7��NZΏJ�����9��ԹUb�����Bb�淴��F㿯��>��Ҵ�ȸ�����7��Vw�(|��J��u<r�������4����W���g]�*��e��p"q5mU�hr������z7�^��N�:B|y����*�窩��"��SOY��G�`��Ƀс���=���c�\|�ee�kO��	C¤foCL~����@(�Ԣ����sE��i�	m.;��)�w�U����s��Sn�@���E���8_OA� �a�������@^��}r����g`qDY��%�W�K�W�>��<�����V?�����YA?�0����?o,���afG7��k�y@♮��kߩ�^��K*��'%��\F�Q�?��8\� |�pO|AQ�r
lH��k��(�'U���x>v�_�'��=��AzP���������ie�S��L�G���q��2�Ҡ��oR�&�I�� ^ �{"���o �C�~&��q��f��b$M�ڼr��f���3��^�;���_a.� -������U�>��gdȣ�$E~l� YSZp�18��?�L��2�݋���� ����1����F�$�ɳ���A�����a��)VI�.,�=��x)� �ص�4"�aK)��Ѩ�ѫ]��оM���X	yy#3�<�MM�4�G�pPN�ov"`�zH��ׂK*H��P}�~;	��iA���kD%CŠ��?�� �i�=.��Ht�&
���bDJ�;h��� l!#ᴉ�v`7��
�Z�/����v�J%����լ��4%B_3h��Չ>1�T�T���G ��g� �PY*��0=�X�̹Q0��Q�Y��/�K{!cU�"��ax�]�3�k��;�r!�9Y�G��"+�!S�uZ�Չd�3��>�Q&������E���8h���{ڋ�~B5t?!��9��E�
i�ME��G�G���-�"��.���5��	.� i+���� ���{�����%��Ʋծ��C�W�	�0D�Fy��5�"p��P�	�'�@2��X�M��4^�_W��
^9�,wO_���E+//)�'��xc�O߰��*��p�2�g��ލ>H����9�q��o������
Rb�O�٥#u}q�cKB'"E%Qi��o��;"�0x�dx1D>K/^������X��i쿷���4�v�fٓ[����Z�}���@�����E;L���9��H=�������^��x;@��3�yO3�������hG�d�\RA�rf���/��EH�]A���	N�]-����>�y��$E���}-|2�%ӧ#�)�G`3�s�Õ����/��-�w�C�u��~o��$��޲
����~k<W�-�vqx)�Dܽ�ui��A�=�8��\RA�e$�H���U�>ÏJ�*I�/)�'ږzy����\�Û��-�nL5�ߤKVFN�3���MGA<�|-����r���߃oCTܐrh3�3�kgKv�l77a���W�_X�.tav�'���m'�v
����h������K*Ht��L�a�k��7l�]�Q,�+����ld>`È(�)ƍ��F��0t���	V٣O~�z�H��T��r��w�MO�&y��;/��[�R�M���U�u�#5̉��,�a?\RAB&Ɛf�JP�f�H99�R� R��~#$����|��<�er&�42S��D���D9ʇ�ge�ZfP�9��H�fMlY�/ƐI��f��F;E�?P)��:��c�wG��C(A���D_N$2�;�|W+��U�z[C�B4?���9��5��-}������,�JU[7��X�`^AT�}��)2�oUY��tD��tT�٬#Lǂ�'�����"�j��>��	��|n�h��.vN�c����	�w���MTk("-EwUydLl�>xQJ�۽�$hι/I]O.����pI��:.��^}�D9z���N�f����6�h����=K�g���ݑ��Z�Z섺n��|��
b�c�vw 8��o��s(���r
	�Hs�Y"��xN�2��~���U%�e%E�ߒ��p��y������P�Qa~����>�A�ؓ2|�{��l`-�y�-�I˻�����S>]L6.���r=(;��{*6\z�-�_�.��7Tؽ����o%|;�#�7���ɫ����~� 	�<pB�����'n���]�Ow��λq�T�x��@q��ݏ&~p1~�� /`G��Sc��C��\���J�����è����%֧Ke՝��%��{� /�n�Nb�BƷ��> v�E�=iSXxj?��3�%���[ٶ�<)��>��;�*xm����;F��s�C+^���ݯ�7έ ���_3~�>��qI�`�U�{g���o�0���)����S5��қ���ih�Z��cJn|�A�x�,���蔣��t�Z���cԣM�9݂�+(�ǀU�U
��Ț���]I5=�1�T}�Ř��#�������_A����$HLǱÕ�"�ւ�o���?��:�D�x�a�~WCA����v�*�le�1����Qߑ�=�7������o��%1�2��`���w�\��n�oB�?	6�~I��o�����1&�~Ҿw����%������o��6�LN5iݙ�A�&g�ڊ��*.��V���@���o$�:	���5=# ��%���{=�da����K���c���\���ۜ�H#�nB@��hs�=h�������t�8��d�zO|���i�V�����@���Ɠ�uN�3���S�_���ހ6iШɂ%���z.^S��2�ys�3tw��h3�e�f�2d �3��=�c{�R\�Yf���c�z�ƞsTy]=���
i��Ȝ�lZ��N�3�Q�!�՘��#�S���n~g���J�M�C�"���\q@������-�˃�*,�9����=�0	=u�*��7znq�zc� ;�_Dy��lv�J�DZ�"ΟY)Ҡǅ\yP	q_b��]��h"?|���ۨ����v���
5]잁`>�����Ӗ���ДR��P�����VЯ�S��F�;��t�� Z�-�,H ��;���6]l���M���x��+G}���O38�1j��j����-;k	wg�k� ~D�����Џ̥U��^�~���Y4��.�F���m`0 ڧg�i��<m;���w���]�P��F���3b��A2��Lk���:p9)1�l)w;��#��o���!
@��(��V�Yx�\�4T�� -z��]�}��碉����-M<R�e`��RFz�{����~������>���"���r��Ƚ8�<{�|@��|�xP۠���Ʊo<�]�Y{���5x�%$�o��9�ׅv>�1����gHy�;�`|q��8xB�gYL��>�u�|�������V>�����m�r ��E�͂��\(T�O�/���<���>����`�$Z��-�U���1�o\����q�s%&�ŗ�)H,,����~S���h2�^�"b%0�ʾgq\N�8
�u������Г���06+8ݛ�&����o��@��/�<���o%�όɚ��5��-��������F�%k2@ǫlz\NA�{I")-1.�����Q�\�7|�L.Q��	��=���������g����~.f3�P9p��������\�Kr�L�h����u��o�)şz8el�t���HI�,�z�F�մ��w�<:4�t����a�\�֖�x,�}���u�<|}Q`\~ɴ��W�y->~���t��Ud�<N@������^��_��p�����}]�!����2���_���T�&�vp'Hf�������~&%���feg�8�D��ڝQ�p<�/	�,�o���q�/8�E|�ӻ���ۍ�S�i�Tv'@
G:�Y�w8b�и�D���o�"���\���#�Һ�VǕI?�o�@�.[�EyM��O���)H̼q$���ږ�)B�֧kA�}��{IQG�jʣ���a�m+?�������UMcĪRO(�Fk�<N,B�B���������C��_4��c�wm���Y�����Z��3�#U���q��Ќ���Ɫ1T��� �+����S����y:�s÷{��ߖ��œ��iZ,���&Zvv��;N�*ƹ�����M�n��ŧ�ú���r�%$�!�>�>�L�[9�"�458�#�Z=���$�����8ڲ�q���٩]!-`��J�r\^�SL>�`�댖F��fl��7��[�VДtgGtC�:Ϲ����/|x�=Β�E�g����р���g�>���gc;�m�?I�������5�<&�P��<����|�E! J���T��p��^
���^{[�d�:@ք���͎�D���� x#|N������)����p���h���mؐ}�v7>�\o�#r��;����vSW+�2J�y����ʘ�}j�ĄQ-?z�;��@���eL��U�D�-j���!���ox?�-I{��u�;�5��H��hV�l_��.��v{5~X�;������(�i����V������8	C�OD�A)E��r}�W��v��+�l�M0�5ͣ7_њt��$����,�cD��ǈ�� �怖�;9rl0t����gr���K����p9	��G9�Q��r���E��B��|+K�&�4G�P�6�!�(	!X��ۦ�q�����W��eK2�� Mw!�< -�]���D�kc�%�G럯F�n*�6�?;6�7^o�Զb,���6[��g�S�m�_waaD���(��`9t8��S��zRKe��?߅��h� �5��![���dW�2R��4 G��J��Y�䆇m�.�OyE{})]�|��Uܑ��sa��6W%r͏�M����w��9�[z��?Ss�P�h�/�����6�5�E��5�[>|#ĲW�j�>�S�2��uK��e�=G�;1�(�gl/�K�ߋ����D�BM81������x��1�S�j�=M��e1-1V��(��w�J�n�4�H.:6�
���}�l+�i��3X"��!�QV\�����Fן&2�@z��rs+�2��)���,n���q����n*�\������[�V�u��bFN3�Y�=Q4��2�� �P,Bͣ��8L��i�e���{�.FCG
(iB>��L謁��' �O�u�
��=!���� ��<�W(:'Y,�0�p~u��E�V�!t��d��mN8�|d� =DJL�ǟ��;E�*9�L��zeT,Q�l�SCS��������
4QS�Ɍ�Ac�L�Oc(wsţ��7(x1/q^�*���o��#b*4I+@�u�F]�Ep��gt1`�%	�Sp9iZ�²�i�2�o�<t#8-�;����U����������������"E�Ei�$a�ᾞ����l�Bb\}�ŗ��`[�)M�U���B�7���8�2�W�QG���`wҎ��W���tM���G2$�����H���
S�@ҽ蝡��g}8�B�j�R+���dr4vI�}��}Õ��
�F�V�D6���`��J��OC��ύūv�X!2���{-l���F��B��h#�{�2}�_)��n��No�5'���m�+h&�����W�lv;�;i�V����=t�9|�������VL�l�`�+ڐaÿ��rN^���΢�uTd�M���iCG�����w�����Ȉ�g3���ځ��ؼAJ��P�7\ ,Ri7�O��$��!R���E��C�0��c�FD�"��^�ʇ>1�"�	����k�y��Brmx�n�&��k���!�Z�-���H@���$�e��W�F|8d��(��`h,v�헦���u%t�E܌Rk���3��]���g��K���}2E��X*T:)=g�Av�U���Knl�r�u��a�1`=����_���"�Ww�>��Pl$�f�yBy1�ۖ��D��V���_�K	g ��O<c�t�XMA�&䯟q�ޟ\�Vi�$�v��c�gA�޸���j�z��T}H^�%��r��Z���iC�ԏtA���aW�1��e�n		����[�7
9�EZ!hOߚO�h�/5*�����2�Aܞf���d���>�����K���`���m�1��h`���`4 ��I���]�]k��$h"�8�P��>��C����6�ґ�ᬨ���9���.����_]��L��l�2x��
=.� ef��R}^A
��/������w,�v�R���U��úP�)�ڴi�H;#�@'�NI��cB���Q����m=*������tJ����(C�F@T��; )$�;Qg®��NA�"�����{7ĸ���=Q�=�䍛�-h�DY����%�g��.i{h��a�u����	�@nG5N�0��,�+`]Y�\R�+�r �S�=S	V�a� 
�<�rl�j���/�<��,\� �v���8m�� nH�3��"4���J	���W��v��dO/� e��]�#*�-�)C���RQ�N��|b/z�cFL��%����Y�ެMS��y�'���E�a�b����lR���D���'��yek):G��X}{���k�)�O~v����H&C)XH[�����kq�ೖQESu��͉&$��t+)K(���DZ���f�fU-����e�JgHg�a���	:�ە��S����?�uJg�`���
$8�� ������~�׮�\CFk�k,BF�["W��w�>�#p4l�Bιp%��4z��e��H�j���B�\��kᲣ[��}/r3�����^ă��-�Q�lZ[E��5�*:����53-���nJ��e8�VA3S�+n�*,{}	�a�"��x���ښR�46R�H-�)�"]w`�>��T�if9a�p�KI���<(A�:@�g��t�ԟ	!k�gR�J;H�|�hJ�ȼ h�o�;�o�k*HT	�M�0�M�5p�8�Q?;謀�g�|��CcA��F�}Q(�l��*aJ�`�la�U�KF��_�/�����҉���UN��{r��~���(qԈ��"�����^�_MT&i�NB-.Ț�|�&�k�I_+P�P��{# ����^�)==f^����o��P���>R�l���[G��x��w/A{48bG�V���&�|��?�98�TV��s�=�YSꞷ�RЖ����LT��!8jU�X�_E9����f���Ʒ.� U!G+��9�}���3�&�>�d��jԤd��]���<'��X�A��9�&8�i�#҈�R%(r��3J���̯ 1���Ͱ$�j�]/v�Hj�)wl*㑳騀��ى�[�ᨋ]��d<�1)����VՇ�WBe�O����1�T	B��XXp�h��bH��*��l�q�~A5l�߉������rd]�I��eT�"D��-_?!{qc�����׼����v6��!r��!��I�㡨FY�:5�'�>	q��X���7��~�������.L�*A�����>uX�S4;pku�L����g��Օ��)�;b���5�@U4����� z^��}���`�'�����Ӹm��Ǻ��A����w�:�mpA	��'�����y���s��Cf0"�%˼�6�J6�j�Kg�<�3D��x!g�y��vA�`j��*i��X�p�����ɯ=6=�{�C�4���J�y�%КsM�?�C��RU�����y~�`n��`C�cn�5��W|ϥ���3�q9�d�_�W�_ym����ݴ�$���p���Z�����Qā��CtV۫<���A�FPo�Rj�oz0�כq,�_�Y��{W���H�� E�G�B����*{�����L&(�TiUao��y��)�Fu�14 �?�9��C�n��CDg����`�6�5������km���{���"����g� Z���#������;W7i䶉,��c�CB��v&���שzt�(N�c.1./�A����������(���UΟ�� ���|LS��~���^���DT�|�y������sc? ON,�S͞�蔣�Y���$_�$+�����)�bS��b*����e#�X5�B+GD��0�
�ឞ��ۻ�8uّ��V+&�>�k"�Ujv$}�w�QO��,+��J�1����dS�d�!+���5V66Խ�N�j���
��o�i!E�W���8�����He��(�ϒδ;sn�gb�!��q@��R@�(a��ش�����Cp�ٸ��� BЎ
��p�Z���Ŀ�|�ٍ���W�`*��^���v�*���g���wҩen�a�TL�����f�"��Ix���b�/�Y�����S��
�[9d]���_���q��Q��{;���EnT5�����-��1í]�@�u]�~M^v���(�O1ݔR`��u�b�U#��X<c~���9G��
NP��r��RІ�.F��;aҹ� �[C:�n�!�eh�z����T\t����*$�b�$���5��Ǿw��]~��J}QR��J�C�u
u�f8z⊓|�{�ꖈ�Y�5ɵq��Rt��	]a�D0�U�xw �h�\�O�K�vT�v�Š�J�.���y�(���(5��	�r�:����l����ΰ��l���d~�
틈|��7��]��hq���	<ZJ�=yf�']�Yg"���V�K*HHV,.t���C_�Ͳ�'�y��ՀX�#��'�ϼ{�b'ݶC�[���1u���%,�v~�W�,x-���6�H�/sܸ�����1C����QE�J���-'S�������tC�D��Ӕ��9&®w��ҍ��]�ޛ��bt)����h�_�D�+4d��װ��RY��.(F�����$r���l�d�sχ��D�R)T!�7M��-#�H�)��sS�Y Y"�W�"��v3Kn���6�{��"J���P�jt�,0.Q$�j�3mK�\��,���eܖ��9hʃ�C]�P-���:�Id�5MȦ�2�gfT4�#�!D�<��:)����ݲ��l�fA��6g:v/Blv^��ƚwv!���j���-&3�SQ�<hw�m5� K]�:(��S4��4��,�M��Dڀ�j��p+��0׊^`\���zEH���\JQ#<ۉG�E鵢k��v��"�,����.�I���׽�ӼX��(��@=ĠYX�F8�ҡw�X��4��{g'�SϿ��C�m*��`]Ae����S�������T��/@�($��T�Cg٬�����⾾�?�!Ѫ^�D@̸9b��]����5%Ȫ�s���TЂ(>�X9�m����Z���#�������䙎?s-$h�'��lkI��}�2�2�?oX�xq��mFh9��:;�JX��
��.B��ڕ��n[@3��f�מ��Q>cX��,pI4�[*L�9�,[m}>�8u~�Z8rw���Ui|HL�yQ%��$6~zGSPxa-��w/.�=G�W�ի�2���r���?�-Zc�� �]��ܧzN������gWx<~�̣�D�&�4��e<�'��$-���?Ȼ3�sn�`�o�%��}U���k�Wl|,]
�)cCT��(
*Q��,����Nv¡
��~>��D��4c{��h����]��E7*��k�2Ï�Z��z�H��#��G62Եi�����>�;���N��WΡowEi��^A��p��U����H4�'f]����`9����#���a*��	�+q���M4)Wr���w�l�h)��\Y'5f|��/Ix�(���!$l�|�,���\�t*ȅܦ����G+��z����]�歨�N�����y!�E'J����O|$W�ć5��W��M�F���= �$ޡ��g��q��*�1n.�0�q���A�b�����r���d������rɘu�������}�=]�`���Cl��-�Q~-�ٯ)�;�NU-�2�\"�{^�(B��N�JQF����� i��Jc�P�Tط���d �`��{�z�my�V�Z-^���V�雧������¡S(�.�ǆ�_�QE��]r(��6��lQ���?&[��s�����ܫtO� �0z�lÂ����rQ��Q���R�
�Z�nӢ����X��k<�,	��%�ŕ���Fm�X�|���1N�Q�����V��ӏG����ꑒ0��p~�ʘ����D�P�I�N:�(ն��}�����A�!t=����'�"�� R�����h��%�*HĩR��ݲ���IO�x����@���ߎb�} 撊q`e򠲇L�#��\ު�X���j[d�K��(�Z��lQ\��8?��_N��KĝX%�V}bK�M[��m*��B������)#)�\J��m�ca�+|�-VҤV����q�d����q�:�]���"ӂDd�"�r+�y�Eцۭ0T@�<�Xk��DA"���GPu��%Т��<��-����m���H����p��@�w�;&�B0�n�� �d�`Y�7�~/�H�J�\����d�F:�����r7W<�e�*�˘-��	��G�"����?�У�Z�ۉ1$��%<����g*���q��i�\qt��_~�_�J�����:�u�n	/�حcPqw�60����cԬW0�^����TJ�ly���~�]�oȖÿ(=�28�t���6��PЖ�SA���c� W�����_�h�����SGB�t�2��8Җ�h�D��.��g��"�v&�y���J��D�y4'��NI���Α�-�N��+*H��`���H�����\ok�E̷�i"�i���� �
�\�X�Y� �����M��Bt��@��I��	w��y'�^f���D�{(?��T���e[�fUe�Q�>4�^9�F��g��9����4�������N�k�
�±*
su��v�a	g��c�}Ŕ�kl�ê��6`	3-�dA$[`���#�_���iZ|��-E۪���z��Rh}��tGV�@��!h�jڅ���uRX���畞>���c�Zo��K��d��[�D�%�ބ�lH6��"A�*a��8C�k�,㭳��.y��=�2�~�oE��tZ���S�=S��3Z�.7�ݣ�(M�?>��
Ru-.���&��W�X*�Rj����M��{�kž|�#)O�3@5�d�Y�
���x������n�kl��Xj��挲����r���OB�ڣ_�c⊞�ϵb�xR�R�Q+)���u��ų�ϊ�<�/�,�ݨ	tX�g䖖8A�_;��Qƕ��/ �|��i�=h�?�����g9s�c�]�7�FK_��/����#&o�����ܭ�7a ���_�[P���������[��C�d�.Ƃ��Sp=��-���2��Њj��H06�B8��<Orx�. R���N瓀5�y����ھu�(�zd�#�t0�:'��_,t<ƕ���-�k>��u+B�'���]�9%Ƀ��^�|$� ����a����ŕ ��6;�M�"jP��*�)�8%>h��9�E�Q%���ׂ�I�����5!�b��-�ZQ)�VA���(���;��l��2(��jJ݆դ���?�S~���>h���K��W�r��N�Sq9kD��%iUX�j�9�tE���p���1Ǖ�E�@fΤ�m��A�T�Y�{�\��Ӵ�0s�U=uxǁ��nOX��Ξ Z��2�5��T���/�En}(�����:���|N����(e<�ٕ������2
-�I�4�6�T���k��[i�'�o����3l� �:�
���,\YGEi\���1fK�-��ү�H���Vq��tѷjm���hk�_5���nx(H?���i�O�?�`���)6hi�h���e˼�Fi���ߩ#T���V�N��o��_��Gk �B�M���hjmY�S�H{�Vdo�؞M�G�\NAZܬ~��Je(�\�솕�`�~J����X�V=Qɑ��Uy9xG"�ӓ(�.x��|��w��� 듉�ȇ�fa
�>ݾ�F0�C���� B�쪮&�@T�C��1]p���%ܫRHK���~�E<�h?���V��Ͻ�����@
�ˠO���$�@N�1�3���%�x|ty��X#�e���d�)�ԱelE��V�_��9Ydd���VӣnT�����(g�
�5��PZFv�?�w��wH�����N5|�9ó�	�Hy5���I�[*�:�x�1��%����}�;����;�J��қs^P�o��y�k�k�ߛh'��Qjb莵��J�s���R��fZ"bN����:}�y|o[�5�������|C��;�X�_W܁h��E���(�"���ڃ�,Z`����\W��5�K-·~_,C���.vh�܋l6�(Aw� 3?~���U-�n"#�Ŵ������z ��&�h]S�L����5�E�����3}.� -����̵Hd2�Z ��B��	��K, ����`x����D�}|}!���<��!������΋a��y�@���yJ*��;
��I_x)v(	|Җ�3�����:��K��3�)��'�`<���Z���;)�F�9���XCX��U��TA��*��狿�E@�nGfie-��V ÿX�L��.�7�RG�Kh\Sۢ6���.ƫ�1 Qz�p�V\�(S9�͇̔y����E�XXu\��b5Q#�u�24�\]�h�#4W6��B(.R���9��_���2Ue�vjZ����,!zXH��(��oĽޢ�w���0dݑwP�����(G��J2��ֽXFsp�gp'C�
���ϣ%�n����a)2�Se�ciW�)� sѓ͊��B; �8oS�a��p9i���Ȃ�����?��I�7P���B�
�"��^��s ��0�k�P�ұ���\�R7p.�=l�˙�,�r$�.E�9�T�FgͰ�d�'ױ� y��g-º���g��ƫ�v��[�Em��J�"���(���=Uɢ� $l�5ޥ�@�m[6d]�����_]�1�4J<V�L�u�����g����]}����h[5>����&i�ʧ���^Aϵ�!�4ͤX��w~�G��+�����bJ�Qʴ�Qǯ�X/Z�c�~P��<g!fح�.���xͷG����bE�j��\(HIZv��Xҩ��Y��3���N#X���d�H4�;e'��2|(`�	����}�n:��oK�lF����m�Hp�|.� �Ն����P~�H��3�Yc�����Dyǁ"�r�3�݂T�"[�z5��IC��6��h�,>w^����'<cQ �w�ԃ�
#Em��ȳm���-�{0�0��&E�i}���J0̺8�u�[֣��FO��|X��vN�&��+6�Ƣ�Z���T���(��������wCn��&���9�)�zGH�n��LV�v����z�nȐkk���G�����yFr�����}%e�����	Q�H�b50�o�|�\EA/T��c����"b��F0��JE�W�*���]������4ߕGxj��OO?T<�lx�s@�L^�n�Wb��Nl�`��e�ʇ��,"O�]�f
�?��I��ع�� 3��(�W�.��}Ԋ��r�ڃ�e\�z{_���(�$FPpݛ��>*�V��ոD	�&�.�!gL��J�3X	4ʡ���$]HP��NWcwog�����߾xzL�;�|�8������74H��%@/�Jj��/.v��se^�,�Z9��1f��'���?PaS��%�SY�nih`�=��Z�N�/�Ok*���Ec��n������Y��C-��f�$$��o�H���4�-v��̲�L����h?j*����Sz-�"��*t���P:�8��Ӑ.� a�M�����x����0��'�J��� I����S����k�����hd���n6I�Fi� ��4�2�q7�i�ɱ�tbA�|>M7(�|xX[t�9�N��l�VgtYe�m�F�VR0�i&�Jp��B��r���(E����bm�t��4����t�?u��.�Zūԭ��$��䙚�T��m.OT�ƮcꖳZ&5e.���(GI�\���A����)(gs�@%�y �i��
yрR^�>��ag=��tƿ���VY/�1b��I�r �F8�y(��
NuSfb��)�fey��\RA����S�O��n�S'�~#��. >�RZ+�w�nM5�#��IH۝Ŋ�5�ֲ���@�Z�0�~5�Z�y�����3�7��{-T��Zbޭ�&��,�O��s���P;����d�L�[��/0q���?�����>-�)Z�,%V��>����ޥH+�(���*�x\C�H�t?�v��ȯi��B�5���^Z'�A f�՜�5F$;�3�tP���F�`-��R�mm��K�����hJ�����U �a��!N�\�6v:�����޻hK���b�s���g�Hz$���IN��{��JHB\|�*�����e�;BH�Qr/����B"�(�#�z�YV�j��hi����U�l�3�Fe�
 ����r_{����igA8�4�9C��x�h�\7�ԡ_�j���B��Γ�:2��tb=��qJ�{����O�Ѯ�Z���䂭l�������&�|yfz��j��P�� �\�얥����SzXL���m�2���U�M�Q�R�ۏyCTv�i(ՔW���z��<Hz�o��C�nև�#���j���Q�Oj���d��??K�h:�0?�Dو>ܑЩ�
7�Jg3|�%n��u��ߏ&���ll	LF��N����Ƣ1���y@:��Ĩv�,��ҾhБE4y��2�Y��fĤO֌���n ��gۜ��%y0��)��U��I�-J��N@�ztr�U�l��*��ˏ�o�+`��7�^�� �o�KFDotn�e���e��:_��˝[p�ϕƢ�-��k����[E��+ԅ���I�N�I�7���֧�~	���Y	��6r�Oe����{:ȅ$Vf��*��ƴ���1[-��ᆼ4��j9�H���z��1Vƺ�(/��)���g��joݫIi��05M���a>�I�+�hǧ|�X8�{a��x~CʷJd�̾x5����,[��uଵ��n�j��o�@��<K��H|�I���,Y���3qR)2T�޷Aף�3bQٮ��&.4�z��#���ه.{���g���t�B��x�:��`��T�c���.�(��,Sr-W�ڙ�zͦ��tn魹���Z�ҷi*3�1��d2l�Ju�h�?��\�����(l����Y
��YHnS lGӧ�F	f��Sk|��e�Z��|j���.��Wf9~�l��;��1&T���C��ρ{�ܡ|�1�|�\�:��͛҄{7�|Am]���{������f��;��NIB�o�f�<#*��{qJ�w�r@�ٰ+QEZ����&Z�{hEi�ݩck[��p[�8�Ð�+�##�X%)|�1W9�e�yo<�\�j9y-Ę&�įJf��Py�i>��ؓ�L���Y<S���֜���V���ֳVxjڕ�6��R��y��nEmK-%�>��dN��e6�:{�<	S*I�n$���mk�S�[�D��VQW�ܢ�"]>���4ƴ*M�� ���J�N��E������p� �'�fAX��/�tά�}�^�J&V�Ơ]5Zh	}U��⟨>�*g��B�5ain곳�t������s���K����e�!��D�L����Ȳ�W9�:ϫZ�D���vY&�����v�d�8�R��}�S�]4�E�l�{m���2�#�c�v�w�	Z/�G�8���H�S)��4�8�rL@�\�QM]����ֲs��&<X�V�{E�E P��rYJ�rr=rd��%%��)��壱���,�NT�z5.�� ��_�O�͈��GVB�ķ��r{���i�B��`�&b)�~Pʼ�"_���V0?�vΧ" T*[Ҍ���xdU�;����K��*
���3�-:j�CC�(2 5��`,����,��6�Q��|���±�R!+�:R�7f�]%�f/�^M3~����m'�$�mNg��Zu�:u�� E(tr��;.�թT0Q�5�s���
�ѡK��J�|_A�hM�&R1~��|�t�c^���9��_���x��`��4��@IF�l�JM��q�I�{U��
�'�d���,��P����p�p�AH
Q��-�d�Pv#'4)����(dM�¬��#k�R�M�?*��Na�O��q�@͛���5��\ LJEx��h�[F	���K�kE�+e$�e�\�rw����*��E�r/��ј�Yw�VPGa�c{�D]&f�ø��b��3E�v�����aΟ���s��X�#��[b1'�ij�mm��*�IU�x�^I����z�ʂJ�=�+)�3���ļO�l V~չ'y����TR�Ebk��dNQ��u�5�c?T����"�X[Ξ�2���Q�wWG�k��*y��xP3�ܕ@�\��9!��d{h���5��r��rEo��o��������@e���8a Q2��_��ì�?~�"]4�\���#b��qѣt�j���ד2����ִY���6��5�)$-�3N���Ho�m��h��=n���߄z9�<��">�T:!E��A"&�3r��t� ҈"���N��/��������i��:�Wt�5!�W�r��/�da�f�$<0��hPy�)R���V��$[t����nneX���wd�d��}Hy�cR"��]9ޞq��Ls�P���w���Ć��sA�`�D�l(0�>\��;��0�{�ی��L�^���Ѵ���keޅS*HL��ЍH�Q-C0�lK�C�I�t�Šs��zO��:Ɔ��B#�(H�6�u�Ǒ�x��4�"��6z%�E^�{M֌U�]G�Kz}��9K[(sJ�Q�33=�([2�[ٖ�iqn54�ns�J��G���A-�&Lի-β��o�8�dW���P��x�v'�*�QH��iT���vju�%��&��[��|G�ᐅ���nF�M�����r�P	�o_��]I�]�c�w��x.?�3�5%XY��w��BY��y>vB᭄�F���Q���A��Ǔ|7MbŴ�T��r�dzOMs<Dd��Y��S*H^x�XQ-8��E�VZ:]I_8面\f����\�R\6L�L����;8HV}'��Y ��%�_���sm��"�M&b�g�Ε��:�F��V�N�|%�g)�|����8[�6���ߡ�^+�w��{.�g��4�\�F�u�UE$�n�	`�m-9�䵌��>����ȧ>���b��넷Bʛ�W�vs��'l�O�����CBj��;d�[2���_̃���~�*@YI��m^�`�[[�����*i�|�6V��UY{�z^��8V[���F��M�����!�}e��P�<��?��f�c���I�/��5�UPK�<��� 0�s
�d����R�*�o�	$L*HI$b�o>?QJ�5�?Q�bg��`mIo{7m�۬��w���⿩��l#�3�D�� 9��v~E)IP5),	k����|#uKYcMэ���˾ԯ|�����RT�.����&I�`v�vY��k����z[z�տ���,
Z�:�4���W�j��yX�96�2�
�Fk%VxaӅOs�L���Nj6	`��]��*��:�i��.��%䅧.y*��1x��ô����l�m\�����i�7?ia3��(�i�����4u��qθ��n�O� ��v��P}9F���u8�=�v�p酛��װ��m3�1pM�Zq'���3k�<�e$uL�da@���ʕ�{)�E/�o�"�ń��>�I	c�0���5���v��1�7���l �za_��ve}���]'c��W�Hɟ
NB��X�j��H3�\ځ(���d�xy���>Tز�cX���:�in����G�n�~�R�J KKjc3�`B$=�b�YT�Ltڍ�~����U�K���X��<��GB�!�{/:���K��s\z�]�o���i/��@zc�sk�kz�JSŹ@+�h�����ݟr���(/�|���7|�-�-��V���j�� �-�9��7�Ŵ�4OVD�['�<Z����� �Z)�U����{ ��硹���0MՔ�+@T�����iH'T���U�B<1��x�%=�)K���#˘�F��6��Ù�f���+��Ѱ��b����V��Fhj+�`q ����i��v:%{��7VaK�G�@Cb�pMEv�JVE;�qS:Qe2��{��_�S:f�{K"Gi����x���
R�c������bl�Ԑ��NAN�`���x;�l6gt��CE�J�ncF#�UHQ��F��I��	�y�n���Ak�s���oS:�E�4��cZ�N|�R�{h��Gk�e���h��>;����Vt��ck���<�yt߷�}=�]eNg!�%5{q��}�	G F��!�~w��=*��̺���̋b˼�|���#��rs�7�r[�KQS�E��ޏK(H�`����_9T=d=���hx+	%��.W��O:>�!6^����}H}7��ëi� ��)��~�ʜ�y��[�,���aΉ����g	f-z�L��������5�"H��^Ar���z�T�z��A������je_p�2��Ag	����5��b�Vۚe�S�Yg����Qe��9���DW�/V֧�Xc�$��gє�2g߲[ECX�f�{iʲ?]IRV�oտՇ�u��5'�������N4���N����f~����wG7����|�����^�PA
,G�p�K %�e�)ۚ�u)�`�5��Ve%0?��WoT0`�=s36�Ys`7,�~�H)Ӕ�w�H�Y?c,P������'�߻����E�,�o�n8#�W�Zqo��w�]���Z�y�2����~���AQ��.�wO� -�˺�A�CV���rD9�����?)
1Ce�����v!*��G.G,�y�3I�L�y��(R�X%LZ�A^g�ɕ�&hX�ԷV=m��̓,ψ��*��*Cou����T�I�3����P���5�9��>O}
�iS���Rʳ��H���y�,��F��PQΏ��S�]=~��k��+��y7P4��i{ήUO+��+���ŤǓ-�RA
m��/�u��5�	&�z�\4AHy� ��ݳ}�z�ZP�#R�4�	�$�������I<��OJN��ҙ�Ty���H��9*Px�{Cj�	��Ӷ�����x�n�YYfӪ��R��� x��6�!�񪹈�r�M�P��\i�I�<���T��
�@��Q�7�_��+燑~��wC��)��g����k��v_��o �Ɛ�}N�x,���=V���اT��b��vfB��p�##�u��0��W�?j\]e�xL�4nQ�_dg�)&X箭��}��B8��dVc3M� �&g��![ñ���_�|j-6��X)��w��S�5��C�;"xE��hy�^�9�"�Z���g��P��<�Ek���.(y�Pj��n����'V�,A`������VeU���d�A8G��q��E��M/^i�y�TvB�=���<Y���=���I��(��^��Z���5�~���wt֋��B�%h������8l�W}��ߧ�ZY�.�<����B['��E�S�T��؉�0�5���
D�L?�w,���X�'M4]�:ߓ�6�塼�r�&�!Kk-?ce��t
�.��[��F�p�*� elMo%���]�[��C	�û�!Zۓ8KW���n��{IZ��oP��\V��F�ͪ���䣭+K-���X{1Ϲ��y��OOm�/�Ưw��
��1�8mr�Z�d#�Q����/v������/P����CiD%Ʒa��ҙ��*<"X����gmO\LV���6����eK/��W��q�p?0�[s�4�M2��)�D�����K�1�jO�U��0��\����k5Efr!%�a�z�VW���1��8c�Pzb� �쒋\^nn��)v�s����»����>��tn��L�ߛ,ӱ��i6dv���W�1���&,�����>:���	���V!X�xow왧[���T�9
nS|��n�$7�s���'��UZt�)N+V�j@ՇͰn�������z�։�X�{�e?��d���*,�w���!���j()�ϟ�	�� Ki�����*��7B{}Z�g���{{[iɿa��l��x���|N�1��K�Okɹ>��#��]��6hW�OB)gf��~ް�ǘ�8��Z h�Ý
R��4��t#�$�oP�n|v�-G�i�s�������q�����m|���g���^�J˨Z*��e5ޮ<�ފq�F_�%Ⱥu5�A���ɯ�����K�7�B9����{b>Em�Cg}
�� ��%����}'!��V�߁3�B�ۘi�h^_�ƃ����c�|��d�� �U��M�_�j�ڌ�g�V��pڍ5]ȋ�H��Wn�L�~��֬u%�#/I���O��;o��(H��yP��;t����Hn�	{i��w����(i�<{��GWL}"��4^�4�1�v�H�Xy|"��bt+���0����7�6���y� Vc�|�A�C�FG���ŭ5W�t�5��·*Uath�<�:I�\TA��@����F*M�^qC'��������a�	{[��Mk�j+��`�'���HB�����W;oEFwoqz3j<؜Mtcv�����C#�<g-A6�9'AY|w��������U9?L��$�� �DN���[��$]=��3c�+�W�!py��%ӽ���d�W���r�]Ic�1����|�}Ÿ��t�9+a��\�n�_����j%y��p#bT�}V���$�V����2���@�;�A�oE�����撼ǐ�,Q������G#1:�ǅ?�7�L)Iv�<7 Nx�\�m���d�__j��J�`K��Oo�Å�
���v=u@����p�:z���A8��)�Eۣ��K
�ߊ/�S���C�vˍ9\�N>oƵ'�'ߎF������B
R���Ԥ��$�1�pKQO?��N-��p��ѥ����B0W6�sW����P�Z�-h�#m��!��b��z�UT���+IE87n���8�hIPc��f�M���876Ŋw�(OGK�o���ݥ�Z\HAZ0 :����T7Bګ����h��T� ��!�:�x;Qc���Ӎ�aՙ���%�'\�x�uH�y���F_
�n`0`M{~�s2�)IW��p1��ޞ]�,8������'��B�v��g���"ѻa܇�����WM+�%t6�'8vXsg��t�{�u�ﵭ��wbH_��%	{�E�ֽc�����6|�2��)e�'��l����{��Y�_����&�?i�8P�y�����|%�F��0.l�;��w�F�h� �m��L?C4�Kp�qKWڣ���� ��6�z
�b�����pވ������Om{!]N����c��	�s|,�r�yĮ6JS��y�LO[����s��V"씧V�j\Y�����)�G�U�!��Q�=�k�9Fi_GkԱu^Ol9�v���m��P&z4�FЮ���gƐf�&��Җ��.���$����E� FJ��o�}9���T�o�1�Aa���{�.��� yP����eX�����R�v� x7Ř�5�M2���!+E76㛚���7�����;%��=o���FB�Q�-���E$�����y���^d-��YO!����qO<�{���5>1�P�竛����]��?k��V.��O����v���Z��@���+�wӚc�#�m�aJ
z��8	�y�k�j�_+��h�>�|s�|��$j�� ��츐<͕4���3���]'�i����� �=Nv�޼�V�£]�Bř��*a�^v����gR�eKo�Ӻ�(��nV��3�Zz�Y_+���˟gaʛAғ[*�O�����P�k��F���FI�lu��Ҫ���1+�UPV��Bm�y�z=]��<�
o�Q7Ƨ±�P5߫����(w�#faX?�]�zi�x�zv�y/P��������F��P���������k�wk2l�gJK���x�3Y�P���k'�?�sT��`��%��R�zJp��pGk�XjT�,�����V5�w�鈗$����`��Іk�)4Zd�k���A�M1�g�L~!����&��-���<�-&�EϘ�/�S*H�q�$��Go��Q���"yRxF�:��oV��il?�	��-�J��I�pti�M�k菶���$���{譨P�˯n.�PbY;�+.G���S�+FYI�(�/��7:�7z�=�#ށs*H+�� Ɇ�{x�'�.0Z���x��͔�Z�b<l��[3��P��(m�jPlK�-+��1o$w_�A���a�-A���"����ÈD��F��ŢP�]�����lъI	�7Bk^�����Y-����)���-|�AA���ஃa#�|�vj�rd\T_�r3�Y ^;d��-Ͻ��O�m�\,\��/
�UUY����pBi�ݓ��*G1/������ �܉Ѥ+%��a�,�Hs#��!���8�Ϥ�ϩ)/4_#d���X��J�N:9�?��t�pzUh$�	�����CV�b��5��*�'(G��v
ԧTZ]����yxC^
MX��A�ӓ��S�7K̟��%;�v�PA� ���"�+�#P�7n��SGO���Y��^`n�'3W�+�~��m��l;h�nC��y>=b��Q�g<I�l��b���������P�fuZ~�ĕU!��1l��g,���uq�Uɴʁ�w�>v^���:rKH�A��_�mTU��ӝ��z.-�:��r�񸈂tBv������:�}Bx�����~�jp��Ԍ�Ɍ��F~o]b�~|y��lx�ᬬ�V�-Z����}�2�v���Lv�`3]�2;4UK�Eu�:��q?��DM�a�ݘ<~\��%�>D��=ϡZ%��(�W�����I�7���(H7n\�{�u���䊥ta-�[�����ʽ[Ż�}4�P��������ʳ4�4�c�������ǭU^W`7Ɇh�W��Gxje�H��3�>�W׭��(ڡ�8��:�*�uYV U:_U�7^�s*HZ�녽q�(,p��9۷�kE�G�Z���ߛo�y>��/�S,Z�R�"����E��U�(� M"��C�]{�tnE���|,�o���ݯT�x��9$?���
7�^5�ά0�7K�7�P[KG#@k���:/��g���"G빒�/�:��]n�I8������y�婶�F�!����r�&�g���/|zk&����W$�b!R7@���J���g�9s��H�Zc��`y�="�#9ðV���х��}�C�	�o.����:�X�V�=嬧yh��ִ{ߪ*L�j���Z����n(j��O�t����1������@}n�x=N� -�0X��u�b�Y�S}����H����9׀���tפ?��N��-E3|#���X�PzV7���rd���ۋR����y=�}�x��dǝ�|�=6_{��P���~�E�������&�A)�Ż��n�'V�V��3н9��A�(FZCw�T�
u���s-�[S'�gĭl���f{����`O?���*J]�V�6�ݼP��| ��(Y����آ>kޭ�����]Qê����B��p%����!�Y+GŞ�7N��P�nܸ:P	q�%	dR0���^J�zk�茼��oS�L�h+��F���m�1�ٯ�XqK\���Q���W`3ݍi?���:�?��� ���r�����CaN����N32����6���ʍ�»OC#>D�� �du�<Դu��,o�k�Z=�Pw�����N�p!i���ƍ��b�'�`VIGLl|Ԕ��ȤT+]!uK(�-���B�)H�U ?�ee��b�9�lW@�DS�e̷RK����?��k�շC��Z�?�(4�&����iM�VT����d -1b�!G�w�p�V��O�Nޖ���ԡc��z�V�z��*oց:���ƽ�g��
Z/�<�X��=����q$H6�B~8\��$�ŗ� �m�%�be�����rD�L#_=�.���&Z_)�0L�E�7%�K呵�*�pe:��+'1�����Mo�7_����*[�Z5m�mVɷp�>g�!<ϡ���y|'�9eu��~��K��0�Xȋ1�¥�Ƕ,]i�]�⃞fi$�w�>b���r%����w�^�qaGPU��0�+oN<�X��c�����--I��<� �5ȿY��h����RT��X�w��ʻ5��S+H�p�aYk۞S�{L�x1 �M�'Fe�g~��#Q$)�Wrx�-#n��"�� Y6\p��i.�sO�����t�6+��-�z��tF�� ���M��r5����R��q1�Ad��ض*�g8�&�f���F�P�Hu*�A
k[r�A��j�0�.eh�!Z�4Z�n"��������դW©�`v.��},Ch��o�X��l�ڴ�@��	��=�$Q�%�N�db]��Y���H��O�ؕ���OH�l�fO����m��>���_G��3hr���ɛ@��҆>؁��[?컅�E�YP��.����w֤\���EI
���M�[����E�<OW%�y��<.C1�F�\Az=��Ŵq�	XKOZ譥��f\K��	h�1y>SP��kw.�<_c�κ����G;�ZbÅ��Eʗ��"H�Ў �b�b�Z����<Zw࿢/��0���H\�
5�瘱_��|��3`Ȑ+$��ַ�����/q��Z9�m��7��dj���3�UNӅvJ���u��+��������V��(l�7n� ��o	I��"����
][�����L�|cB�
%��c�B%�R��v����ۑ���ΌvK*����bk~:/.L�\x��u�>,c� ��a��y �/���[�ӂ}�VGW5k�X�H�^�S��fj�
������3���{��
�a��ݸ�U����Z���VX�sT&zʥJ�k�d��S#9�(���%Tp!ʯ�[����G�PbX��`]�%�f�:�Eق�%��*�E�/���`
��D_�V4m��V�ƄK�<f�@)�N�ÌX�#�M��C�Av��ש����h�s$�_���R����h�VI�U�$�%�O΃")�W9R�`�d(����"�Zu�V@a��Vֿ���<���Y|�]P{M�����o�S+HP�7_����Yo�XK�Rʁ��ǁ���ڇ�3Uoe��^���H�k�e�����G�cR;����(�,�m.«��V`>��5$W���Y�w�h$�ʄ����BN��x���+Ŭ��R_^�`mg��dGۄ�e��B1'��*���Ǹ��K��f�{jϐ�_넜�J�	��Q�a�o�=�[����量�ѣy�	h�ڃx��8���z�+ڹƔQ�:N�� A1`d�\0��.������2H�p���zڜQ|n��{�bɞ���
AQ��Ip��m¿ǩ�V缧���~F���2����0L�Y��c��e�d�NM���A��<1�� ��"�I��*�C��ʪ�%xy�3�u�v7�#�%I�J�j�<�<���`+Q���1y�'��$!?N�Y���ܬo.���/�r��U��-d�ʞ���_���CQ+�z��`
�eĪ���Y.�G��UUm�o���1�E 3��F,�D������)��@����0�� ]t�#�)��FXɣ%͗Ϯ������;�Q��4���7J'�,�`o�z3W6d>D,�,,�8��T�����@Y_�����h{����I��c�IW�4����|wA>����Q���?A�ReV�Jrzr�w�^��o���H����V�[s�ڢ_z{�ޢV���ґs�u��� z��8�iH*��Q���x�X0{H�H�¹���-gF�#s�-�]D�
��+�ǶR���ɧ�ʍ�A,#풤G'e=����K�V����֌��ʗ�U�oS)�t���Tt #B��qɓ�dn�a+�Ci��+hr���EW/gV ��].�6T~�%dg����V2w�fA��+Kz�@�����)�Z7��T%zE�ȨF���!�@o��B������R1���j�[��r,����ܒ�W<����Ȑ����y�Ċ5<���B
R��Zg��7����qc=<ml��N���[���O��� ������,�1p`�n���cuH҅+߹ָ1��26��9�a�ҭ�O��p���N��h�N�5�#H�r����J��t3]л�ݎ�V�e�.��9�$���1Xq����؊e����b���_�<��&��t�p�ۼ�?�6
9��M�\yU�}hC��+�������ފoں�XPiC�2<�e#��<&yW��֒ 0�c*/���8��㝌����{�fH���<�.����xԛe�+HQHۼ�f$���O�w7Ns)����w.h��!�U�c�-Д��|���y����qZ���G�F��ϕ�A�ޅԒkaz��C�Ө`��5�Pj/.-�Lg��J�}ɒa�������N�D����(}#,9a����J�hk-��I9b�]q�-I���v
�e�B�k�L��ߵ��4��N<K�g{��U�)�#�C�T2=��mkfב-�.̊���LJ�\^R*��Oi�;9�Z-�gn�ѝ3J�LUvx�(�[�k�l<����V�>G�Ȋ޿o&�*H����1����封�hrZ����x��O�?���͉>������!�d6&��0� Z%�j�dJzI�g�{)ˌet�� �{{Y*���0����U���U;4'��Q���I�bM�
SN�>��C�����<{�'%oA�޷JUfB��\��U�ԥ�FZL�� �g� ���>�^ϨKoA��(�S�b_�n!���B���g�!P&���?N���nVg��c�(�kR���`y!�#P����k�Ii�T�yl!ȒP$1��#�S>ir�Loa b�&�_�����:JY����g���~UبN�~�J� �dT�w��q=IX@鏴��K�2Yq!/2/�
�����/%��D���VT���x����� 	�^��� ^#��3��cK������[��YB.�O�4n�G�I���0JB~ڑ�N1�9Ņ"�,��:>v��r)����j̳�ݍ���̷�������n#�m��'�?�Y��>��]���EL�=��M�V��D��RB-˔�����x _OLIr�R�|'��4�ɼt�VqY�������]�֨���dE2�׷ �rI���8}�a�x��Q�'~�(5o��*մLO��J~'�1��G������4�"�8�D㉌b�����Ϗ�Ӳ*��S\����^���U;6�X�[YG�
��
� �d9R�5<-vyho!B��+p�y���q�1�N�K������vs
�X�)L���_�d�P����-�|�\&����H�s��]��gq.ǀ�׾­|�yJ�M{�ؑ���Ng����� )�୪$`O�� `��qQ_r��.����BZ���Bj��J'$A��)A�I-{T�]V�\�����=�[t���L�RT20l5���M1l2`��F?A�s�a�Z��"���Q�:61O�{�:�:��<��X����|p�����w�Bj��O����stnh�r�.�J������]���i� ɲ�T�Y�?{����g�ЮA�{���w�����onv�J�%�.�b	��{�O��($�3�Xz�[���}t�P*_?��+9	��]O$��鲠ZZ�~z�e&���Y\�3�O|�7�{�Gh�</+n�H*TġZ�{6�H���[��D��Q*��4����N\OA�s+��4�q��g�7� �[�i����f/���~��ě�g�w�9{Ac��M"��")&1>	ʉ��.�kꗢ�0��JB�����S ;�8y�g]ī?n�5��:%+d�Q�Y�Y۪�ҭ��J���J%I�������=��-:��~|��w_&G�eOK�֤⛔���9f��5�ۅ���/�՛����8��,�K�=FE�H�H�Lg[�����I�$mzQ�~�EQ�p��}ƶ�E�!��bm��t_����sq)p$�kE.1\��hZ{��<���2�����zp������[fs?[� �]`[y��{`q3��h'9^v�!�GE_��'v9��J��m�!E�F���������������7ަ]
��	��Q_��$ܒFed��3'����4�k��~@�9>�s�+p-�h���X��(�LF�y.�|�S�'��3�Q�A�X؆N�)�������?��a'j�����f�(|f+0�?Y�8%����D�	�aE��u�����ݸs'�S�VS��~�X@�Q>�����JQ�cu~B+L���Cxu���s�򷃿�r�����+J��|�&b�,j�;��$�,���ϣ��l�svӼ��?��ά�����\��y�</]�GJr�0�0N�?KhVh����g�6WF�^E��e%~�b�T�_�r?��?���~�)������0>旎�3���`�]:��(֜VN��I�?�8�ǯ�߸q�g�H1�i-49���v�LǍ9��]b�(N�F�#�K��<�P#���ۂ�[��:��B����ˊ��������/�/��q3�3_�)�B�E�H:�]��	2]��S]��嫽]~֍�"fM�A'y�,��ɔ��R�x����gSd���[�`��hh���=]�y(
������r�F r�Œ7yƔ��wedɌ��0�u���<��n��*�����:D���y	K�H[��1�	�E��'���<R�y<���t?�����{V�@��К����:?�抬��'Q���pzH���_7�?������p���\\A
�g�x��x��ODhҹ&9k�����р��œ�
�O���q�u?�sT���6�������{��E�R��s\5��0z�G����/�N};�?���������ߎ�5~���f%4�?v���z�0c�bb��$���0�3��s���&2,�v�w�E�(nU�gN!�F����T-�`����m���O7-����Z�|���!�h�<d�$@;��	�ԩ��-VE5P�㽗��\��$=7ʆ6�w��
��y�;;�u�#�NL ����d�u4
��uhK�e� �����q����b��=�"�����N[���Z��+619#NUJە@�qy�&A�L'�*SOJa�
O'��NP���P.o�Z$�Gi��߼��=�����mt!��!Y�$F�F 9fz4������ ��>�A���g5�4�BV����!+iY���G����8��-^�^�}X5��K:7�4�_�kD�ɲ���ǯ����o�}�r��.��k� �ԙ����!���*�`�q��+n��w�����?���ү*�|���H��w�m8�+E� 	ZԕNƥF�3�₿U6_o��`�m��gؖ�G{��|���x�j���v~& eBXv�,��.*�k��`"i��̦�N�uh�c�}{Uf��g�<�箱�D� "�p�F�Sf2<��Մҡ�����E�),�?Zb�;qK9�8�<� &�5����&�d�S�{�U5oΘR ?��aK���SͿA�]��LD3��0)%�e���:я���
l��!��QN'6YS�Oj�>]ۚE�	��
A5�8�{�}&I��3\��<�š�3�63�5Zj�N��(I�p���R�[o���u�	�0u��CJ׽�!��"e�w�%�(�L�� ��y�J�sV~���}`�JV���<�����!�1��>��2��807�$��~�29�GƋ�  �6K�i���9��"���(�il,�����\T�sQTբ+��$-�a5��TCwLN�щwpb�?��ܜ_��	���?��?����=.�9�_�����j$���+�0�h�h�kq������3�i9i�+E~�0�T��x.+��/[����?����~�?ހ��]l@�����ho옉�Fg/�/��|�!r:�"2���͑N�at�71_<��aH��.��\6����Eo�{�(���>7��6~��4��6�?��?O�o�%$	��Suέ�bW3��%.�ѣ���hh��:��Ń�X�nN�[���$[Y���&�%D�D*����x�i������B�\��}3�f[1�3�_ �����j�|�+��\���(�M�6�ؗ�&��TDH��ٖ^�А��]��/~�8��9{pC򽉶���Å,����~>�̕�hj=0�K���Ŕ�.}�W}6�R�g��l��:�8	V� @�a�TJ�Q�"���1k�U;"}&����w$�@w��R�y�f���Z�|�.�I	�m���R���ijI��͈�@���V�?$e)��:��˒�v��,V<
�s�b�
]^���n6�Q�qS�́���dB�PxX��ͱ��v&Ld��Ù<P�mI�u'/��znu���N�+���q�iC�B� %�A�kY�ڌ��\9�*.�F�Nawۏ*Hu�n�^��qD6��G�A�P��Y��W�u�y8��O+�!���Ο�ɑV���!V�D5��#%Ge�b~"n�b��� ƦT����`|yo��JPP�0�s�H�/�%%���K�}���k'|�v7�6����u��S�q^��F|v΋�4[���Z�=��#ч�3W��/��S:�		5�Vy]8p<��9"V���G�@��!bl*���%5:�^yP�Ȍ�gƍŞ��,��v���s��������&'"/T�tQ�LWq��2''ڌ^���C�?���d_�r�����+l�w�ٔ� d(��ˤ�F+�Ѱue������P���w������veĺ��f�ʤp���'�=��M0�>@��r`e:l��}���Z��@����t���`C�i�J��t���٦C���߱���ʚ;��x���ɻ�8�"�m�`��W�$ʾ���T-�ȅj>&*�8mBS��"���#��b+��3�!��Ĵ����@�D
�J�k�F��^>��E9R�	zF������,*�\�$�EzF�l:g�eM�nc�0ok�Q�#���E"�\8U	}�'=sT2.�e�l2�� (��~�U$�խZY��zY�TD9^�j6t��Xߙ4�u����6niP�M(�߫�(�d�&S�:L�����>��Ga�� ��(�Δ9ξ|N�]-RJ%�X.��T��,�+�+�Mz]9���Ԭ5H�����R&Ĳi<�u7���̀ݩ�����P%I	�ݰ+2�G"�3Et�i:7��{JA�8Ut�o�U,$��z�� ��6M� �c�!��HJ
_���Шt�t̂\�K}�>�7I���IY��-2�ƕ���ڜU�O�ʷ�w%!�Ŷ����,�hb��v���1ѹ�8��S�aX�ފ��_�Gւ2�ɐ\_cR���)\�h��[����^�Rc_���@浱��8��Ԑ�4�� 2�`f��4}��6�SA��C�������ڧ��畐��z��BH��.�,n�q�CoE+4Yߖ�K��mFJH�>P�J�\�:fZ�Syb�ǁ�	Iܴ#k!L��W�]=���|��
�JJ��9��;¿���l@*�4aI���`���$Wz�Q��\O�\c�mb>̜+��ߨ�V�δ.��\I�T�)ӭ!���hN�I9��å�P���&x�C��1�QX���K۬b}A��C`��X�]�ӛSxc8F�v�|k;��	s�*������s��p����XX��8qĲU�j����9�� ^?�����Ў>e~6�|�w�'���x�W�%A0�J����rL�q�`E�S�
*����4���5fv��S��b.�4��J�L
<������ϩ �?�na�t�pׇE�ݚ���&��!��.mGb����1��$l�q�W �\��-?��3�,[�%?[?�N,R�h,�ɉ��N�!:c��1�e�?/�&]�-�U��`T�hѫ��# �x��B�BQ�w��on������=ի�w��d���� �t����E۞��9֑��K-)�x���S�<��h��K;�Sp:�~�v�^�\R0���ч�ٺpR
E�1q��\!J�5�#��]��FJ� �W�H�ʆ��.��w%?�gG��$�f��L8�όC�i�)�lW���4�vC��o�d��rg�b�����|/<8���JN��"��s�uC����@}��&��^S\A�h���
MK���
"=1*�yQL%K(َ|j�+s�H��bI�z3�KU18��T�d�6���?�4��0!+���x?�A>�4�ͮ8V��F��DP/h�����`�@v��F����^�E�FJ.R��R��۔\%�ud0�zTm41hi7�K�%��䏦�Z���/����pҠKV+_�\·�<y���ºJ���L������]/,�n�)�]������ �?�E�a��׬��o�4��$���z�+mC�R�V�F�G���8�V0��d�ͱ��8�Gr�б6�3��.�t�n��$.�
-Y$"V���.nW����{�fd�n���S�`ShY��J.��y���9�gq�Z�+�r]Z�ɰ!��ƷM�qE+CtGO���m�,� ��Oך��3��:�@�Z�7�G��X���vV9�� �/���b�+=��ׇ�!E�e�l������x�[�Sȅ�S*H���@��?����vc=�-s�B�Y�}<R1jtn��_�����?U�I�n��M���	[�@1xI���4���]�2xP�e3ĕ=:CS���<Y+zo��DTF+?R ��*O��I�#)uP+�ç�����KEs�|�@a���9�c�?���ʷ��a�y�"Y/��d@�2F#��}���߭Q0(�8.�$�a��*�R���!�LJ��������%�|~L��wJ1rz7n��
�fl���4��������ݫ�E��5�Fk5W��\.��g)��-g+��5�Ry�	
������ ��#�mKn��ϔH��"�Y�����s��R�إ���VY�Ӂ�"��T;舯M͚jL�|��%{�J[�+��9�V�_��F-���nd��6���>��Dm�������*Fp&�ݤ$��{4��΢y#�m�y�6N��,Ad��X�p|��ͷ$O�_��Ha��}�o���]�f�ٛ)�33���H�������C�z��D������I���ȹ���p�(�SAٻaq�#������!�͍�ᙗ�	�%p+��;&M"���I)�I�bQ�,b�P�I�eq �˙�H�{_�B9�ɴE�RH7ӧ�#�DM*9L�q�b�/�%�,+WÎ�����=�Z"�W�l� &�t_��nԎڼ���i���g-}�w3}$��m9���P@�̨�� yCE�K�\L欀��n��g6����ݬ[�OR���'�z#EP��0g�qDn��5j
��ǎ�*-0�U�=F����\.�{��餠�R���i�o4�Q4�dg4�����ib���^_)�Nm�n+��ޘ�!y<T�d�H���8CU������pBi[�����Q�\��d5��$Mu%�2ה�Fd��^F.�g�H�B�,�9���E@[,��ǝ5,��ջf���1V�E�e�U�M��)
By%-m�L�󥞑�h5-�$FB�W��ۥF��z�~G�R}tN�Gc��k��Գ�L���+��^��j���0��B�Vc�){���>z�I�\����q#,�0GN��ډO��o�uǤ��P`*�C���b��|%ƍ�pB�|���A����ʞ�i�8�]/������0EX�<N���5ߌ��H
F�}���(g�͹V���m�y)pdOv�?SY���ӒoYw)�-vnL>!+���P��U�mg��^~&�۟�e镡O��k����hZ��z�6W�lIs[��v��3�ց5�-q�����h�F�/F�=�ؠ�9�E� �Q�*J����%�9��+Vl�_�[A* �+1qܸ,z������,�%:a\��a�b�g�5��l�"k��m�,�
0��/���p�"(�lV����v�[�kY5��V�u��թ��{�>�n)_a�h9���&��Z���c�������0;�z�,NH��=��blB.��&,C��af�iҙR�B}Fs:v���]���d�����֊q�1:v儊�Y�(�x�V}�d5VY����
���d+L-�jh	c#��{���݆;$NEA�-M�V����l�њÏą���e�1:�ߍV�4	$�� ������9��|le���b���e����ϻ�f~�p>7�iie��7���&�O{uE��D���c�`�:�x�ϲ���;�т��wK�=����K>�E/� -X���u�W�R��+Wy�*Wʻ�����F�m���J��ت�����zҙ�Z�g�cD�b�[��[�����4�v�ʒE!���kf���x�+k����l���mH��Pw����V�ԍY_]�Ϸ�4��V�r�XA�>ݻ�=��l��Mn| 
k?8��.B��=��Hb$d���du,�a�$�=k�-�d_9�N��@�2���;O��/�3���-a:�I�>���[�
+t�NbAR=��'�7��כ����9F{�n�J��R�9�к��I@C���|�y���Gô�d�Dg�,��%��>AX��ۨp�t��5��QY���6�U�[.�GH�-h��b{�r�q�%�	r:�K�JDfQrZy�'�es�4ɋ��5��ґ�|H��8�HC���R{ �v|>u*0���(}S���t�PAb�bk�1�h|x�d��wby�T�o���6�U������&�A��&Lkk�єh����#kh	&t/�w4��-�k��_��Ap�앥솙O�6�X�z�{�q��,�1��ؔ��s��<����쎂>?������eWJCR�ׂw��S���P�����>"�(�GJr|��v�^����������	CGI���e�<d%&4�`��|8�U�̰�?���B��� �6�@R�e��4HE��L������CW��ӥ�*H�p��ς�0vrH���ޟ�m�ƥ�6�a�ǻ���պl�n�ZI�:�˧���m�+]�[c�;}{����M">��G�9�=:$�K��U����ĝ���Z��-	��x�6�V���8���_~i��Ḯ����
)�����Q`��fx=��j��&��-�#a�w�h��L�DwF-�JR�٢�Sg�ϟr�֒��$�hL�%x�w��B�}na+�OO�Zs��+�zm�b�s���vlK3nt����[r$A����ڶe���m��=x1�SNg[
��'���빸����/G�!��`�-A�m����e�yl�[}jđ��^�NF���*J����]�E9�4����t�&�Wu�8~��$ w]<Iq���.�n?�%�b�?`<�ĞO0q�Y�Ù�iO�y�>>�O���j��c3epO�+�Z��<Ҩ�4^�rkߍ�DC.����{>BA�B"��������/���GM.��i��^��RĿ��~Oq��d�d�����R��bg��9%���h����	�#+��D"�#�������r4�V'�>!�����o���P"�^ڤ;w���y3쳷���z�8·���N%��g���%�+���zj��0�k����s��\PA���c�|�X��7��w�`"���  
՟�?��~���,�[޿�e�h�Ԃ	�@�(?Xy��V�:�*i��W0{@��(6�q�K8|�8�!*��'B����@dPٱ�JV5�����ߥ��pI��U�.#V�v�2�;��8a��J@+kY(����+b�(4,���K-�T�Dc�6��3VV�V��ޝ7^p_繎�
�d���8%�CV���;洔���O�O��-G$~��v1&Q�Z�`��(��l�ީ��w���mM��l��Q#����������z�%����^3���a�'���\N@�'R\@"F̮�)�/k*��[}W�=�^����C ����Ë�8�x�!�
�s�;���@%j���W��4��?0�#���	������h��N�,�wI>��x�Vb��A�����dop����p�5)2R�pNӠ�`[b�"�yA3�VA�A	��Ք�"����_���2-�2X���/��(}��k�@p=QNU1���*��΋pA���&�=^�OG-�F�7,��*���ëy�v^���ZI������%�􎬫�¾~䊱��+Jb)��.1�^���mg)*����C�k����Pf�p��+��;$�sk0��k6���Y�%-���Q���,��𛞳���jzcJ:W���R`��xIV���0�x9��$����f0�o�
#�}�u�;fm>���]6N�ZI��n��u�'0�7v��dv^��,�W3ƼR ,��bOa}��w4�R�^7����J��=��F�t��|��gc�J.1~��3��^iA��x�w9��]K ���̋o�]	�S�o2ec|��|~K�{e��_���ݸ1�*HzIu����p��Q+��Ls��p��/��Hnf/G%���G;F=?Y8Zذ���1q\��M���)$_c�����r��9Ц4_yp{s>��)#�l\���ڒ3v=�^f���|�T���Z��*qǸp����u)��ܓ�neTG��~�����؏���2��I�~Ox7�~�y����L���{m>� ?/6�y,W�X��'s�#
�>kzk�	��Ǘ���B�E:7T���or{J:�s��]ԥ��W��Æ:nT���%�v��ߍ#�	�"0fW�@�1�4��<�����2����1t���	ƈD�1����T�#��m[����fw�@�����
�������cxa�|I��[�6��p�z#�J����%,H�;�kd�/�+��}9����ڤ]�>�L�,��H�L�e^��%.*2�^��gF?�����F�h�����Wd|9Ϙ��SP�hX�l*rUU�%aX;�<[B�J%X��̕�M��t�������w�Gm$���B�te{����;��˩������¶8��e���ĕ���$Y�uXW��}���M��삇否�����#���j˙;���'�sx��q=�E_�l�����Y(�x�PA���W~NNwvB3	۬\ZX�rĭ�J��bm�{a��FS�V�J���"��.����V��C������ˍ��>,0ϑ$A�忕�� ^�g�� q� ��]���::sSP�lzI_Y�L�>OK���b��,�~���Z�����~\�̍1Z�<�l;s�Z��3����$i����� I/4n��.���H_���`l=�Mo��UJVk��8e?�%�HH�$�vK���w�]I-WAiJ��ԇ���vn�	�1�7t�	�����t���F�H�E+i��)��s��������t!�3T����-B=�d�La�ʣ��eD�R�`����&�:|E:��} ����(���vM�տ��ߪ��u��$$��=@�/��B���{��R-B����{JPo��ϱն��?W��#��J�4X�� ��'_m��e���˖�N� /Q����C�G�ǜ��:Z!�Y��Aнt�]#1��Y��O5�A�a��ۑ��G
<-�[[[S���1���z�g���[�����)�hcTȭ~�H5Z;�0ң�u�joN:M�96�ح��ޞ��J������^}B��U|sL{�����Yid�aZ�ەÍgᛶB�RA��$h���ߠ���O�6�la}S�F�:vg �
Kem�8����k����I>���zy"\�w�q�'B,UR�r���� ��գV�#�A���varIۄ>~V8��q7G������@���/ԑV�#�}�c�0�K�8��.��I��'|�!���|_5��Mug�V�hՁV�FYoR��!����f��[�Ӂ��X8[��=���k+�Q�C���So� ε��hH�on�/�pH&���bXCke�������r޽,y['�o,��xU�e	���]���v���$���x�b������+�~��_Lq�E�e�-]�Oܸ$nI�ې/������4�������P(1�
Yt��r=3%J��$��s��I������8�S��ژ�2�r��Zf����;e$�V�(�[+�ړg]`ȫ�4���BVp�2�u����2B�o*�)ɏ�9?�9=��n�2�W�i��ׯ�A��J[�'?2n,���ߤHV���hU�
�Y�kI�@F+���A�B6.��_�'(l^�ɩ e��slU"�D�~@PmbQ��b%8O�>(BV��F��i?��卌,���O�[AZ����EuvDέ�s �����B��Qk�Q�t�V�
OJ�	�:��i��W$��5k}p���L��S��.s��	5˽
�rdrg����/k�߽\g+>��S����h@r��ғ@� )(l6xߊ�JR�,^��G,f,w��LwV�*��%:��V��݊��H�7V��|�O��V$:�tn�[�;��b�I��V���;��'�[��	Eݼ����ʇ$���]F?]�c���@�����z�*�O��GE+�E~�9��wx�����V�?���E��0.����U4�|�Z�]���(�bd��[�]�娈1#���Ug�n�'⹊D��3�x�[�_�+�b4���z� b���a߄o��=&�qY����!��S��'��
R�e̖r�E�o#��`-�=�A��B�4�����~�,i�%�33`����pN`��������VF��o=����xXc"���R��Q"�L�Iy��)LgQx/�KL"��(x<Z�i{t�[A�q�����ނ�J�~$�o�$���`V�����-�4�xy����úv�M=g�Mq�cG+��s\5�%��V����H%mE�g��*��n<'T� ���Gv���Vy�d�y��Uz����2WHl�Ź��L�+T�1W�D����	)��,R��I�*��ap�oi5ˈJ��~�.���΃�+�Z&���=��.j@��A]J��� ��'��(�B�a �w�sPV�~�d�(j��A�A��B���xi`l7��JiE¢�=��n@q���F�\1{&L�\&�������Zy���:���dY(z��e����r8�_����3H_��'T��O��r�����\�;�x��0��:�[L
�������!���DZP܊X��P�P��/y��1�$��l�?U�R�&�L�(�W�8��p]�uQ���� �zQ���E���������h�6���|��~a��5+S��滍�c�L�[�-z)<��x�Td=��tE���Jې|w���w�1�^zP��2��|�o�n@�ϕUY�Tn�o�^7~�!f��_!L�K���V����5�6���M)�)��t�Wy�(����S^�&}Jә}�i�VO�����{�
�&��X�v-�q�7���+HA0�/]i�J� �<�8
��j\��ڻ(��5�𕃑���޼~�w�ߞP
gk �ݲ��Umhᚮ5��������u4[ :�j���2�/�5[��d�3�V`�?b�����N������Y�T#	*���Nl�K�d��]�<�5#&'�[�؎Cd�/���'�vM�O����1"�,`<{�[+�^����o��[��y���'��N��^B<���OI�9���,z�y%�~�籽��u�{�v�H^���%U>
�h��}��t��p}㥹�*u�[Iڃ�o��⚽}�7n\�0�����9�� �?ѩ��[7�Z{F�H:�������*ﾡ������?���e�b��ƍ�
R:���5@�R�~k��	ê脅�=�2<��k�8���aw�4��o�z�=q�<��~��XM��w����'�x7<�޻�Y��<%A�Y]�Y�Bw4����&K[�W�Rsڜ��g\����72�
����N"�`��h��Qh�1)Ga��؞9dn��sq)]~K|B3:�y_	vK�P�Ll��U��3��:��?�&�4����}������N����`(�������:�^J��{��a`M>3=�Sx�Q8����=4Ԝ���c�{1��	(�e�翹p@b�R ӓ��B�<�]ݙ��n����0nk�����W�x~e���ʢ򎶮�ն�$=-KE�{ )�|Ҥ�� �:Bs���,�Jτ���1����#�'���sa�;�4X���Q4���v٤��6B����|�Gt�I�s@��/���n|'�0�l-v���y�tлJf��U����h4V޽E�:��>筞�[�N��,�<�����WL�}(���3�T�����:�`��Ab�&7��n�|��*��.+��^=�Rǳ�e���F^C4�4���8�r��2橔U:��dD�uTG���b�8'�'g�O,W��ę��[A���F���G��-5��A��H��mV��A�h�;]N��>@���K���6R�����m�ɕ�B z[�X8�.]"^�lFkY�^'P�=ܓi �Su�����-1�
%�9}�4���6��7��Y7n<T����rږ�em{�7�SZJ��c���Qڅ���4����1����r�ga�x�F?B���/ވ������ؠ�3,C|�v�����R��(h���ls��C�E���i��a,7/"k��vI8��Cpk�ρҙ�/9�*H��&6Bf����iA�$(0�ĝy�]�=�%���x�1��z��~�粽.M��ֱ�t�M�vސ������ �)E}�d?��eh��r��@+k�wz��^m�:��GͬzN��j����h��n�Q�!�O�+���̔h��B��
^�h0�۽�<c�J[��>��o�
m�9��LO.��z�D+��)�#�+���O��{��\�j�}��^��F�Dt�㗼b���+E�!}�m���T�`�p-%=Oq ���M0�hL����7킒��Z�*Zdy���Q�r�m�S��Q,�aq�>R ̍�_�
�gc��={#8v:z�z��fi�44������k�X�V�ҪI�3�[�{��=ߍ�e�/�9�h~J��T�WI������k3�{п_�5��2و�+
?��eԸ2:T��N��km�)�2�nW*r[��$6�qC%���,=d�}�[���m���\})9W���)&��>�$y�����9���W���,���������CeR" o�ҵ<��.��9��'%@��� �]������(����jqbh��^��XL��{�8��F�ƿAj=���ܥ]�+���Goc��1��d�w჻��9���
��y��pri�W���-]#�Q�F��f�7T���E��S��.���2!H���-���7�����c(��',���x���P/w����V��:�7�(\�8� �(d>\Εtrwm�c"��7��}�VϖA�#��ι{�̐��[f��-*���n ֓^T.��o�-v.�w����1�غ�
��_0\O� YC��6}���W�4݃��Q��7tx��H,Zx϶�c�Iȑ�H/��d�u���i���: y/�h" �v㞨.~�V�e6Uj$0"�q�\�sfrن�2I7��|B�b����`.8��R}�q6�;�;�{A#އ�
����0�v��ُH�_Dm'�v�w4" \f0{���;o���r���"�jM�%LZ��Ѝ������Z#���Nb�:<Y:n��h�b���;Ff3��%��l�-VC�m��m�c�^��W���֡�pH��-mi?!��x[rNX[�Ҹ2o�TyN|�W�>��N� -�6�o���'Y*#A�����o�4��V"�L��u�Np	�"-�m��Y�W4�
?쎮V">F�މ�+X�U7�"|�͓-�>I�kn'��yaKbaD}w����-���ChMG遍/�����#4��$@�S�Q\
�d��;��)�(D>�K]ȧD�~���E�����t��p��J��"����6/=�Uڔ��VΦ���V�G]�?j2J���on	�c�s2��kM��]-_)H��t�a�憂T8o���0�|78�ѴC瑸����uN�����ڽ�3��� qA�����G���B��g��J���>p�ķvGf��2�9
�d���-i'aa6�i�-�}���)�.<׼����sa0��J-������i�9�����G2�Y.�&��9&����W�hP$b2�BS���ot���A�V��<��%}Պ�94P
����~Z[� 4��o�BĴҶ��E7�4G�g:���%�����E����.��[ȑ��B'�J���K:�4&&��,�Br�|�|���{��+����ļR��0-������y~yoyV�;�_��qL���'� �"�P�8�:[Hr���.^B�=�_�������e�L��WGs�f�wK�e��I.�ӷi����z7�n�$#$���>��Ω q|zܸa!�7�kn3@rg�s	�ɳ�2+�Yh�B���_���Jv[r�D���F�(��W�^�����*:�My�2�L�����Ch#�$�U�9}�Uz�k|�h �cb� Z.�g�R�p��G��EXA���?W�
�)���;��DX3������D�{�(4B>L��p��ք�N��[��*@��=(���FQ������)�o��<��ʆ�o�����ѹ�98 ˲�X��oLW���.@������ܥcXVD| �j;T(�0�,��S����ů��J�8��!��h.+�~�H�!>v��H8�!cHWY�7d߱�`*�JA�"ҍs�
R���*A� [���I��B��Oˈ�e�.	�Q�G�@
`�0��&�d´�#j`-���|r?�{�γ�@IT��K7�^���1��2���iiMjB�oy�^�R�Ū��xOi�cXZ^�0�ᎩO�3`L��-�ߐ��V����0��q�����@_�X����-ɕ)(�ǽ vvց���2P�Z�,2&���n��T������M��`1�C˄���/\�E�����$W���uC4��`K��}@L�C�)�Mw4��K$s9�W���-���A� ��I)��iU�]/>�sZ�����*�q�~�>�^�Ԥ}��sc��4o���
��F�����CE��[�Պ������z�-�"��$]hKE��
�F_���>F��gN䶛Qw���Z��.NR��&I�9g�2�<��+yrl�mIaB�����+�gR�byRI��}7n�� %󅶓B_ekĳ�{,���6�5%��I�Uګ��.�ª�':?��,B+��BC����@�I9�0Fu��P��CL��ñ��#MfRT�@��9y�G�z�P�,�!]%	�Tyrq9�mG�mP��\����tg�7X�y�虤^���Of��M���]j��D[[�ψV9'/�^9n�YP�e(1��b�?AQ��5o�V����+}x���e9n�"�.W�F,���7�'V���<9'3�c����q��5�V�>D�.,`J}���K�"5��!D�˘�
��q֙�R��$�\�����g�0I�<��BE{��r�ޣ]�Ɔ�9�.y��c�33wbN5�hL��Z��f���3p�uJ{G��c�d�uf�N�J[���~]A�a{���{<4(`��-�nq�>�)�9��=S�#o7BQ*S��o+�"Ѧz���,i ~T-R%�yFc��yp"��*�X�G�ۓ!c��{䋴dV$r�,U� �Lz���>O�y#�N��E���;\4 �O�J	����8v�Y�][�V����WK��so��7,�WArG�!������jtx�����k�èd�\�ʓ	�j�
6��0�VP�%\+�=���J^�Pt��V�K��S3pn`;�ȩ[���*��:WH[���� ��QxRJS;�����oOz��(�by���kZ"r�ʏ"�$���ʲ�l���Ӗ�HM���Ԯ�á�-b����'���>�W�qef0V�JzA
o�����.����b{�3G�xy[�:d%�ݸq	�XA��Gpk���IL�&ݸ�ո�ɚ	Zʾ�d��jE���ǠT�ه���3B�k76���_=fi���E޾�-͆Y����b�fEK�$!:�be����Z}��i�i)��>� ���9�Y������L-�\N�����޶��8��`ucB�n-��Uݟ�<08oX�5�u����ӵ�v}���&�zf����	H��+�u��+|^SP2��*}�hY��LE�
M�i�����H��|��o򱰒F�r�i'�_�ykN7΅+H��$&C5>�;��#y\ݖ�Hނ���Sn�D���d��l����]\X��[.�����( %�ar�M�͕��M�Bbc�>���X����E�N>�]��F�*$���DQ���z��d��v�BA.v~U1ی�M�$�'�,�&!k?���f�ȳ�7�F;�����uq�� �E�X5��Y?��t�5c��*n_hū|�4+I��1cQ�\� Τ	�k"�w1�̷lF�y)��b�v��h��$�
����E��4£�իX2��|hg^�F���9G ��L��k�n�x.� E�Kf��N�?�Iw�ֻC�K�q7N��.��kx
䳕V��6����f��z��&^���sOq0Swr8ĥ7&�[UN�w��2�p�2�!�� ha�.�\;Ԫ��8\k�	�}��0�O����e��o��P�]X8����D7�L����(�i��g�Rml�~)�� �@:�M�宑���)ޔR�}�Eݥ��Y�#C�%����Y�)�SLIr�tB�b�(�;��J"��J&�/ѹz�
�߱�#���|�:~�qM�q>*��iC���.��|��V���-ݸ�� J�����c��Z���P����'vda�X���{�r&m��&��)Z)5��I�]V����T�<�&u�����Z���ќgca0�I�$Eq�.cv��-עZ@n�>��km�kG�H�MT�g�D/��1�͓���>&�lWRZ���5K���E�9U8yN,�?>��6��?#"o�`��LCԊ�6�H3a��8���A�;&`ϳ*��|�k��8���q���
��%�R���h�;��^57ǥ]��d����V��n���ZAJ��Ƥ����Jh�Ra�ܓy��2�H�󭭝	b.�E�6��2\3�
Ȫ��!
|���f�h���3��p��Z[)��d�5Q�,%�$�0K,U�Б�{] C�ꂹZJ���(��Q5.��,xMx
�iQ����=5Ԧ�SSSDq���T��Ja����RC�2�	״U��������%�"`�I	��+m��䦔}�[���09�2�T$ږ3�+��J����S�u�$zCj�(�������������B��\I�o���Zf�"�l^^y�����5s�8�1�K�+Y�j�}�ȭ��C%?�)�����"O������"�^*g��r���9YΘ�D��Z:�D�IYS8Gƪ\w`��x��k�p��9p^i��l��ƍ��V���kD1�/���.���C���(�5�ʄ)
I�(L�F1Y��a�i�ZWe��H��)��G-�\��M�3��x�'��o�Qx)��kt3씦���x~[�b��з���4�ZE&|)���W�Y�)Ui,~�U�n���^�?����7��CZ?p")��| S��g����쬶k'T�a�M�Xș̜9�\�HK�ax�o��Rn����f����Q;}�t��pW)�2��{Ƣh�fRBl�q����:�·������߷�s��8�����b��'�d�qi�H�X�T4�VM<yKDVq|:)])�͎��ǉiJ��e�]"@r�*�S�I��*���	�
\Me�#քG
��O~�pE��"��y���K�>�n���)�v�z��l�-���v�q�E*��v��a0$m��rL6͏�X\z/+s�;�6�45O~���J���9Pwn+�XX��xh������mNws��c���Iw�y�qN��Y4$�ǁК)��MAHl%��C�f���D_�ɹ|�n���w�ۂ��9����F���(������V9�2V^���"Xɿ�mQH|Ә�a��v�_� (�I�4���U�5�T����%ˋ	�
#�"�2Ӎ+�
R�ݧC��y��%+�����ٵ�&�*s	��׉�{�d���^��.��Q�5d��◬��=�F���g��K�����P �y+_�i
+o��J��/:٨�=(v���0���i�
��aE8��"���))��5M.�<��H��YC����VK�q`X�|�,*�}O��(6_wT ��}���\�͠��K!P̋���80L��)��2���
��U�sP�L���f�E��okc�RS��^��?Fڤ��i]��mw�A�'�AÀTja���z�n�Q��9/��ü�7n�83.� ��q�9��:p����'�B��k�����W������w�����q����.��a���01y��5��{�T3ݺ^~�*��8��C1�ƾD��VE�B[���q�X�[\E�n�9��T�(If���꓈�Ng�:>�yQ~~�M�C�pg���:�UZ� �m�97�*�%�sn��*6�=���.}��5qY�c��Ӆ�(������I�����٠���e=�Q;>~�HOs�L����rT%���w��n�4��p��|�C�@�d�
+m��k���s���V֟h:Eq�+^��c�h�ͦ�c�Ft��ƍw�B
҂� �g����wkK��o+8�_y�z��~� ����H�������??1Aݳ���W۰,�xGy�j�C�c�j^e��渝����$rȂ��3��,m�<��$=��w�q�`˶�vp8�b��F"N~K؏o��AG���G���_
��Q��g{Xv��1B1���ʗ����hA�_�����JI�i{�/���[.\x����k`=5a��IC	���~���\�W�'R,����7�7}D��N�B=�t����.ɷ�2�v���j�Viw�rf��A�^�� �4���J-��L�am�&SK�[�}�W���&7�
�U���i��QUR�2���K9b�f�]���V��?��C��FZ�����96aD:��ւB��x�;����ܿ>��z|],���A��%F-*HT���>����-��[��Z�02k2�g���{e�qM����ꚪ�ݍ؈}����鮪����H� �dɒ}�e�ǶD�
�F�*t��g"?6<KQP��%h�]�Q�>������׿8x��lLSTn��\c��O�
{H�خ���2�`'ܯ2�O�~����"q���Iɜ����Ln�����~�yY����]Za����ˢ1Ĭ�h~;4���A{yһ�x��W��^�p�E��\4n���+ko��g*'|Nk�~��a���/fփnV-w��E^��Wp���%i�
E�P��B'�e������ǼZlǿ�����w���������_��:�N<<��˶Ay.��*퐩��}���
&���5���J_S
F:��l����m	+�û���<��G��/�{}vv������v���c��Y[���ۇ����E)�;%���o�8�5��ɾ�k�L��j�d*�IW��%W nh-���޴�)�J"%tv_�G��/���_���?����@�c|~����@��7��R3
�]j�L�MF�ե�v�1qM�k�&�*@I��QO�!?�6��-+G���J�w��3PS��B7B0P�]ͧІ�5H���+�����������o��0��\C:'5�0��[њ̴����
�����8�tOс0�W'�hw�zl�1��83� ��$����ڏˊ�w쏰¤iv'��v�����;3Fȑa ǀ�J�_��(�J��on�������~=4��ۑQ��/�y�Ȳ0���U3y�$_���,�</�8Fh>�*�uۚ#������(�ňZB������#,�ͼ:��%�=�٘�]��SVd����J��tc;٘Me��H�qI\�@����<�)��*��$��޳�
������>M,�T�p�b��7�ʽ��A~�Z�X�i���>N�Pc>�g�2V�i�&e�]Jٛ+HQ�PO<���M]O���2����3bH'0AW���jiU����*����"Ҡ����6{O��>`�۴������uE$[3��(����"�E������L�c+HC�V����\N�*�4�D���l�����p�T��_1~�b���:�i-ko�4i8�H������//��x�y���� x�H#��YC�H�A��f����~��]ߪ0�"����Q�d�d���`��� ���qe�^Q�f
��&�o���D�q�RBÈ�mb��76U	v�9��ʷ�
��t�x{��hI(+��+A�?���Xd�{	�ֽ4����)|�W�q�\�\���('�`����'�s��.{�ԇ���a����:�Y�Mk�z��*��c^#O����_i���� �+#{qp�`�XU2��a����m�/�/-IR��|֮�g��#��ⶲW��@�!����|ǀ���f�Fa{���I'/72�S[��2Ӳ�r�W���l��qn���2�yQ���x����W��O*׮�T {4o�A�?-׾����%�w��9��� ��%t��6������,�ǭ'ݸnI��y�_���슻�9x�hr��P�F��P�x�%{
  ��IDATzh�w3�+{��ʂ^����M�ޒ�T��]^v�в�8�:���U0�k�n5�IP����yD4�VvzR9F��5�m�k�R�\FG��H2�YU���葵�_q+18^�z[J��F[��>Q?^HT�V�)*�Q1+k���蠇�k��O�5�#m.�P�����󿌺�Kb������Fhy(]�����<�ֵ�\Ͼ�8�b+���;����l�}X��GVM�4���8!��*�B�0���8!��iq����7�m =��8�4��Ms�Ǩ2��-I���V���{�$,�������㵂c�%c*e�{��]� �R�[f��2�wnh u�|bXF��H,}��v�s�g+iM'�,�
�������H�a�Q��+*�KX"�;��2\}�<� T1\m���	�hMR@�a.� ��{r�en�Wa�B�Tjc;�Y��F�k%Ƣ��-z�hp�?[%��{b�{>�v��c��ؕ��Y�zd�b�#�9(�I���M@f�Z��V���������5)=�a>�L,��g���~@XU��g3R�?��~���e.�
�k�tA7�	�5�<T�߁�:��/����'�k]����d�B!x��(��/��KX
�C��zE'^�㿃a���� ��b~F}�ƨv����{�~~A��D����X<!8�-K��B}x6ym���\4E+<L�l�hg���6�D��>?�L�'�+����`����s���u�q95i�A_h����B�S=�
ߢA���,���qA���7��!�t�q')Z���z�������Ui�Z��DHlh�z�\�m(�bL���.ļ@�/4G�E;(�D��.�׈��d�VH��3�Bߦ>Ou8\(���V+#��u����I�U{ٺg����
��������Ƥ<
�~��ݸ�R\�@ډ[ݸq�}I�+�%���LA��Ջ��]���O�O�X�F��f!�F��9���O�){�g�&;�ވGx���4����� '����	~O ��o�ɑ��J��$hRX�B�1�v30��dō�F���؃��)��_�Ė�q|Dz���A<� �-�82t�ƣZ�2����an�d����'K{�>����\\�@�/�f���a!щe�Ha��չ��V��������'�e�d���/Ϫ���r��/`姍"�Mž9����E�i(��Ӧ�M���j���������g_�uz�-:A�ݴ@���½���әu��v�¡i��� -�hE&c`�Nz�t�����̀�&�t}I>�����o�+�
�ˍ��`h2nR�H@�e�U��<�#��n'ٰ�PM��=<	�vtZ �a���	�au7�5��o�����!|�iJ䍵�6�I�l�=6���.���V��@�eV�A�������\R��uE[/��P:�
	�)��~V]���S�����qc��� R\9�ɽ�,�Z�܎�AQ��:���Vc%�Y�M)�k�C	x�Y��q��(�(�Ehw��l5�A�Qe�8ڢ(E�J�b;E�,�.`�8K��}^l�Z��o=x��g�6����Sk[7#�	(�5N	���/	x�6ŧg���L��9
�RH��m�Yz�s
��y�A��Y�S;���<?z�����)W�z5����9�ET�P�M�Ѿ;*�[]�Wۮ�3"}�|=�4`�AL�V�ţx/QP�Q���W0N��l�H-����͈lé��.�
M�s8IH�~⍅���𭐯
'�Qd}R98_z�aع@�=5���
M��Vų�xx��e��A%�l/������k3�Y���[w��>x	귎�n��ӳ������W�I�e$>˕�g�ˊ����axg���LbV�%��{\`��DY:3�Dj��gB�*�*��e����иF5�B�2=�4Ñh��S^2^K���:x���Ҥ����=��>���^���i�a���'ŷb�P5vJ�ξ�������&E�+I�A��x����-_����'�c�I�&dV��qB�c��g}t\p��Ŕ��d�����=c��rM]����'���6��
?T��vta����/�����Z�Z����������1��i=��Ё��ȰI,��)�t��-G3���&U�f���	x,�����Q�2`�m��}��k9_!X�d�Py%�;zQ��/uFR�,e�z��u}���v�f��4��{����+��×�]�_IQ�u����MNX�W�S]� P����a�#��S<��T`f��y�WM]�槓9W����� l�����gR3E6付��Ώ���}�Jb^0�C���
��P/*�Y_������\
-��oX&��H��}Y~v_Ỻ&g׋�0'�gapY�Q�h���ӥ��	e�8��ٹ�3�P�8�`E��5�o�1�X�xr�)�Xx�/]��4�z��ܿq�=(֍���Tad�|�r��[��f�s+A(�����������tɧ[T����k"{9�Q�ھ���4*��$�!�+�Y����wp��3kxh,�ʎ�~��W��Bq�$#X�z:�M�\�c�}鲺�2}U���=����dD���\��8�:��)�ƍsp9Iz+N4OҞ�����Os�V�EA?���(�SoeK?�,�,A����ɻ��x�Ȇ]�볓��y�x�g{����_v3�ǂ1F�ZI�üe)O!?'���P3���"��)����J�5�H{��)�v�6�>?~\v�<�l���-���J��J���(���û���e��Tv得?�����.w��}L�M�C1M��;�s�S�o'��9O�6���_i�-�,�Z�MG|��ɾ�E�Ǿ��û��ˈ��kx?�3��0��Ű�PY�������Z�
��s����Y�q�&�P8M����ԻH;��.��0^�s�ڃ��\�b*6�S\k���[���I���SI� k����u����}�X�=���8�
���r��Oz�3��/�4�D��2m���՘�k�]s��*���^�Ǒ��R���k��1��������˄Կ@
sy�q����2�.�^p#d4��2o|�,�jE���&agvY���V��D}Z{k9�}�y�Ϻ���W���h�p�)��r�6��!6ΎA��X<^�	6*Fe����	yee��"_�v��������pM��L�r���$��f�?�K�j�R�TT!9M�
����9	�PW/��al�~��٢{L�FRMa�^����/+���9��ħ[}6Χ�	�B�c�P��y]C��G OA����"��yܩqP]GsdJ !Ӽb=��P��� ��`keiU��pO��x˂3Z�T��e:�b&H��r�(0��6b)m�ܫk�W�EW��6�%�-�9�!�>�F7�T?Yr��}��\�2�b�vω�s���,-�{��Zhk5�c�Hk3.�ɇGv�Q�w �3~��=�z	��R6�Y�����g=&˧���Z_ߺ�Ua��>\�4��ט�4>7.n$�W��
��D�_��]������%��am��Q/3=�$|���Of��������	G�V��%�Xʨ�ޗ
��@�٬����q?@�k:FC���9�|�TG�J����T�vv{�W��M��ʃ1O��A�/2�G !��g�TA}����i|�k����ѕ������-��}|�43�&0������(�ǅ$�ב-�Vʸ��F���Ђ�%�/K�t��ۅ����:� [��Y*Yu��_���ޗ)
e��^�P����X�n�o��K�b�OK�lU����c����s�WO糾�#�q�y����s��o�2�"E���-eM�2W���	g���_Q.��]1�Z�F�!�ɔ�)�H=
x�{����kP�4_���aC�F34�@'Ƕa����<,����r%�0c	ǸIln�Y��V�Z�:���Zq�h���G�ya�iJt�O�?�U
�)ww�z(�����Ҙ��ƍ��N�-�ѪLBqh���g�Ρ��J'���kI�c��?P.]���Օ��A�O�,��)�5��j��j�&\d�
��y��p��!������[۱[΄"��r)�ƍO�$�r�0U�nC�,�9��r�)��=^�d�G��ߥ�j��ۤ�޼�Z�K�C�i��}�2K������Ki�ګ���ڌ�U�����С���!{ܵz��mꚹg�C{Xb��SʰHk�׋޹�kX��<�c��Vǌ$�3�ڄ�
���/|�ĸQ���mh]��e���\�@"D!�����|ܸ�)��n�B���{�:���ӏ�o��	D�U�ɡ��*���[ǈ=����
���'�̞tғW�嵽鋯�{f< 2Z[CF�GL��#Ow��@�&҂�bT����H�����jRY�Yyv�&����wO���ۺ�g��ڥ�\@������(�����V��J����4K�d�[e��ګT���B�F��3���i�݀��F#׶��@�=T�*�U�F�8�O��[���	�<�H�c5��qm���2���v��5Q�� ~�|K���Z���q	Z�J=�P���70�VqVk^^��΄���E������p���H����eyG���<Of<��holG��l9S�XQ�3^���eyl��0�a/=����1���^|��ثu{�.П�^��J�H|zƢّ�[���p�|��[닽�ڳ���k�?�?>C���h�R�{�X���Pџ���ԚZ��sWF���n=��u��W��b'��\N���;�^(W9�e���B>|�o�K�B%�i�;���E�%�I�۩�fƳ����%;����P���b����ȩ��&q偺Y
�����Ьo�-q�%��&�U�K�E�7�<B��:Y��j�1cbn��ZnA�y#��3�T�֤y�_���{���8��k����^�7�5$�C�/|�qc Ch���|�s�cu���T�fC����,�V<T����v$�3b����}W�ṋ�V7����`�:�J.��o���#=����ws���:�T��ynEbĨ�Qt7DÔϏk�>L�4��7�n��A�m�����֛�[��C���( <O?5:D}����hZ��4^ï`����]㿣y��<�Y�Q��;�n$�o^�z\�@jP�M87>sϨzf��OE���Bz?��ؐ��?���"#�8���Z9��� ���]t*��j�5��
 �5Ɨ�i�ie�1^�ƍ�ϒ>�\��a�sv���:to+�u�_w��l��nh����K�����7~�&���?X��FͿj
�����Ϯ��������囖/���x�x��R%��^�9Tg����V y�SrW�=�4`K�������ո��nr�:��@ӌwn��Ƨ��hd�:W~�<���|�{s�i�� 1�6;X޽Oi�V���ӻ
S��=�1��O��K�=�����K������#��X��^���W�J/��_]7o��xU1��Fz�"������3�������U��1��iw{Y$��ȏ~G�-.~Z����~	G��(�*��ڍ��H��v�a ���$��@��h�X}�lݻ����O�?���A��`���=�p�k���s��G2<ɿ��H�jc�I�,��F�;�6�vb�_ǩr.YNs��:��#��wW�H7n�<��J��V����A��*`g/|o?w��F�Oƃ���.��a^e���K}:��P�KE��U7�A����{����;��<|��Tsd옿(��7�4.3�{��贶��P�JGO�'@���~���o��n��L�V >e5�Jh��ʤrU����ɺ�HH�v�>+#��I�J����WSJӑ����Ċ4;�"��0�I�{�����[�B:$n�~���Cf,G���L�_Y���[�;qų�[1}:���>��
�тN�Ox~C���OAO�~����KC�@~B�>~���y?��w��9�{{gxT?�&n� �nT����1��ǭ�У�~oT�s������t0���F���^�x9��U��NFd��l.�>!N{�a(�wV�'�{8fv}Bf���W�j�_f$�"�>ۗڻ��!x?I�ҍ7n��!�֞o����b�|�\-Y�̹qq.�~�`hύ�����qK���%àq�^~$F��WtZk����-�'�"z#��au/]=�����t�ƛ�+���(�7�@�f�Z����[+���e1��w1��4<J�{͕w��	��� n ic���>od A��Jrq��y��g��5��~�1<��G����=���VZ�\�1���α-mӨ�v������[��{�p��Ko�c�:���y}�U�?od �.Z��7n�0l9[�ƍO�=�7�/P=��ù3��$u�Ꞝ�LCO8x|�[}-��_������.`qs�)~�3�bҁ���<	j[úy`^W~z�Bu�����Q#(���*z���?ё����Iw�ڍ�(��o�d�
n���Mw� �8of �Q���27>���A�O�т��$?A��Q@ox��?��+�p�ƍ7�GH�ѐ>Ʋ�7z�*R�Qqot�q$�^�v�3^!���#��w��~���Z�E�����W�ϤU�SïX���%n���"q�
ݸ:��@,�2:^ӈe�q�(l�Ћ�E�_����
M��(��f\�~�𦙅�A�S▱�N-"o:h}��Ą2��8��qmb�qI�#�rA�}�@|�����W�Ɗ�2�@�&��ݸqqX(:�k �� ߳G�u*^I�ݯg�����	"���`�<��EQ��{��yx���C��i;�#�YKx�G7.��ᖵW5�0N�35[8ҡ7n\��Ҳ�~-�I,l�ΰ$��tzw���x�턿q��pI	�$ZL�Ms�T/�O�[��x[��jh����-h���>��{�j�r.����i���p��0*�9Q�q�Q��J>D���9P�;䔽/D!S�[*��4��
��<!,C��<鴝7߸q��@'�*�8�ߙ��0�H�ݛ������ݸ�s��h�c�P1�U�Z��)�Y�JJʇ3���R�sYX]�����T�u6��<Hr��%ъ�[p�i*�#1�r��!3�������|���b2CZ��7*��J����(�vڽ�&�pG�ƨAA��D�F��5o�,�,��I�ZQWM�v����3��ޮq�P��odx��8ѥ�I���y���n�_�(㈹rV�-
��>�k��4�#`�s���B�|B����Fh�C���|(M�Zr��t�]qj�*���%�?�>���Lַ����׻��-ÏԱF �G঩�1���}Vǀ�r�����=%�b�M?G�"7�J(pvop�ƍ���A0����N��7����=��ᨮ��ײ�F�=�O'�qe ��f"�^�&�|タi�������:����ٸ�����k�����ס䵽=�}�':���_�x��^�]�$ɣ���f����c0Jk֦�#V���׸��ն{�8�!��z_ܫd���{���!��!+A�m����U܋H�U�+H����B7���@������^M&]�7M�^Z{���1�0~���6ΠG�����ݸ���jw-\�@���i�{1n\;xzJ���!hJ���^	:=�~�6��n��x���Q�FԄ�^0�ȧ\�P�7.�'��.m A��ɧ��⭏��x��uB���^���A��7�R��:��Eƅ�g~a��[K��-d��K��z%t��x�%[�?ٙ�g�!�`��|�]I�D�g^F;����A�=&�k������c�^�ׯ5s/m ـ�{�?�O��uy�o�W�v����g*P���cUl�_�2|��d|/���M;��/-�Û)���^l�{�V6���&�1dO�.k^�5���j�z�ɹ���Ui����i�5
������m$���J_�.g -$2�2��a}��rI;ܚ�r�A��򅬟1-G�uC�ġ%��(�w�^�]Ưc��70j����۬��(p_�*�Iv��}PC��h
�
������r�[�R�2��1�N�D���q8nOѫ��ϋ���oNS����\�·��;M��������.W�၆�Sd6mT���β��[�^>�XAc�^Az�1�4�~3�:�f������	!$O'Hy�g^��UZ?d޾|cO�Í�p牪�p�#��Z}z�.A]�K-'6(�7k��h�6��ċ�3ԟ�
�~L�����^h�ݶ�k 
�-�Ag�.7�>V�gA�D(������jN��KR)[@�EX��:3�>G1�²�QY
���|utc6۞��Y��
��}�XMI�۲�r��@�,�|�]�so���BJ�	2m��	�/�}�λaa��Aߺb������qt��� \�⿠��<ы�#�(]y|,��gak���h|�00@��&�\��r�����Zy?/�c3@}~4+C|�-�W��h���u�YY�7�Q���25Z}\��'c��i]����I��#2�5��9W���(�ArAO�y�H�Hn[�5�>�(b�H�c���L1���p�_cpn��i��a�}!7v�V�þ�z`�5���Osa0]�KzI!�?	|� �D^�4�l?�QY柷��3���j��rRYv�-�:?��'��<˲l��v�S�@��ܳ��Vx�d���P��V�`����x��/taO�Z��{dt5P �+C�{c�����,S֥_L�,�����L��j!c��ӳՐ9�!u��ɽ��|�_����bpf�a��]�����gW��#��|F��� ���r]��w��~���)yH�U���Vz�{��X�<l���q>�4��g�.2�ۅe(�#l����;4�,cH�@�rꯣ�|�'�3�D�so����o=:D��������D��r���c�*jJ�y���4������Mɴ�m���d�s_uJ3�J��잵�u��~OZ�,`a�#��P؂�L��$�}�d�TƮ�4�޻�KW���qž���|�*.�t䘅\�&@#HC�p��ΓWJ��#"�tqI��;]�^�@���k����G<�L3���O'Y�+�~]��h-%Wt��s9��?��M��ǉ����p|�5�oJ�<e��D��w�y�͒�<2�a��09��_ ��B=�����v ���qW�6��Y�,<3״�w��Z�N�YYQ�|HC�]�_Y/A�+Y��2�f^�����p�3�Y�(9�U]X���YN#�b\���S-ٴc�,�WG�V��=ɕ�X@�0W��@�˕|����1b>8B>f�)�L�<_�SAN$j��k�Q������e|v����S˽�xd���̯7��\
c#���}K|y��Rgy��<O��P(�D�z9I��M����B��Q�.�E�<�ɲeD�a*���j�5�	̩�I�=}=��|�e����#���5<�Y�C�������H�)hs�2������ͤi#C�K�0��d�`�����H�=q�r�����?yt.n t��?���q9��a������Լ;�g���!�#�����0������5��骯=-k��H("�����֔�n�+i��O�c���!թ+4g�j��_�)��Z�=k��+����F/4T�=y�e�Vgo��7z��)s㽸� �,K��#�8��������s��}�<�	����9�o׵�5v
��t���CMF��x��ޗg^��h*�bF�r�3qۘ���&h�E�f�����]U���������o�7�Fg�嵤7%��䢽�DN{��x݅1��*�*�*ș�E rDE��;�)^&�s���UC�)_%�[r�F���� n��ǀ�_��C���sYE�fc_i�*���I���Ѵ7�r>���	4R��o�+��N$-�XB���ʛ�E�tp�p�����ֆ��IcE�7k�܃�������CW����8���>��7у��l��P�@����w^�K��ۺz�V���U�N9�Wd�yOe�4�2�c��-��aZc���ATQ"���ۀ<G~/}��/�KI�X��+3h��98[�^�@�zR#J,[(�JY��Ν*���N8%���F!���Q�a���'_O��A����������� 곖������[ُ�*u��4fh �j���8�NRHj��k��̭щ�-l�Y��k� 4,$ɣ���;W�E`S�gl==��9��(����*)w=6Z��X��@�r�.�;٘�&7AS��0l�t���=�,�U�|Eє��5P�m�N�{�Ko�8f}\�[m-�e�4���$�]�~m�`�GM��~v��7���	W��e��(��
��~�ز�4]��[@lҒ��?�2]Z�����ಊ��+M�ˣ��A�۟��Z��5��K~�7@�D��tl=��3"�Jdz��>w22�r�/{%Q��O*��LCi�O�R��U�G�l�Lbsɑt&.i i�n�-�1房��s��Q�GBz�9#d��w�Jސ��[�bJ*� |�	plBz��]��H��˅teov���f
/_�ѹ-��V�����Ԣ�B��ި�rw�ӣ��++S��9�f�7��Td���~ �LI+2�ν�����!9�-w�n4T/�!scW�)न&)7��g�JI�E��+E�������v6=�i��d�s�0�i<�,�åJ'�ѷ�l����:�t�d5�M���*L�ʰ垠����_���p��
�終��<G.�%�͟��=;�΁A�32U窔���ʃ}�Ɯ��`�=2�Q�
�(_UR�E��ŀ,������ɂWE��|?�4�p#s����k�O���Gܧu��g>�y����s��<`�9
5���Zg���=��������M� �׭+�E��k����k�LOi��d �:�)Z.1�$m<k�=�)Yn�)��"RZSI���|�N�V�}�w~`��ʣo� E��а��Ji3A��ָ"]C�D��C�m:�b��$?n\�&0vr�e��%��a)�$���<;�<R�+��Y�B�;�"�s���+I���-_��W���w���0�����\�+!3�&=m+�`11��#̣�;rK 5����g���I1��O)���H��P����Ώq>Y��ݥ��
Hm��h/�$Nf���Ӿ6nd�i3]�@�j ����qM@E10`j�Qѵś+�G��M��9�C�R�\�X�M���z���e�lcjG�N��+��ޥ&�t��<�ln�Z�Ԟm��B�B�)�M���R�h�gnЄAj¸`���S��=Te�M ��4�yZk��1�l���*Χ��I�u���Jwӡ����r;�'+�ymG@��v��2���!��HC��p{�w�F�:��8���'V��N�Z�dE�Tk��^V�*S�R����J��fG���L���*���2�i����\e��Q@)� ��d1�T��c9m�a>�����>u&~�A>:m�q���y�riX��R�R��NaY�;y:g��9Z���FJ��Qà�����B���[Ɇ���$qR�$-�T��imh=�������
�q�w��t���\|�ÕT�i�Ѳs�*@�-� �#�A�=���r�O�;4�f��ȣڃ�6��5�b��� �KGy7�/u���l�/'�Z�m)�� }��$=�����-)��&"�:ut~0g�j,<�� �jo����ɿJF�Cv0�&"����S.y���ɞ�c�2�c�zGz�̛�r���W��$��5�MC/�ٝf�;�3��)�e�ㇺ~!L�����dϕ�u��Vd��K��{�� @q����C��y��A����g�`�c�7\�d�{��V0��W�$�|����R`c������l1�M�۸���
~�����2�f�x���#imL�����G���6�=�j�Ȟ�!�2J"Ů�r�z'�6�B8ձ數�6�u�9����R�8vc���j��L'+HL@�$��� �Q꬛��z5��?=���J��F�8kz{}j�*�'To�\=O�^�@��$��*˛�'�(�o�
�V�������2�cUtk�RI9�����]�H�TcPX�F�m�̘{c�\E���PS�7װ2U<�*�^]½�d��w�gY�9���g̴��R�0�|�G*�E�?[sЮ����_�t�D���7�h��G�s�>��((���Ʊ�����Jf^W�B�J))��	��`�����hLp��֣o�|�y#���x����g #��/���9��g*{����22g��͋��^������~����c������t4Q�XM�I&��� �|o�D&��\A>i���z������n%��S�	�ᶟ%�£�'u�9�&�(�\$�0m���λ���
�~z#1>�?��7nx���>��O� ��V��>�B8ӦuY�� �N�J�f� �Hֺ��6l�� �+
aH)f߫@��9!#���e���)<HðΓ�)]���4U��5��3{a��HG����� 0��NQFښW�q:=,�^�K���(���{����1y��B����EV!�O�a��K�&���{��Z	��S}�o�S`���]�GG ��g|3Փ�i�c�W���:�7�d�ה���a�HH_3m!�&Oy��5Y�k~��/�^n�˩����ur�f�|V!�y�'�����y6,��gބi��ʛ=W���YBP�61YM՛�}=��p����������<m�%PSC=��'�BB<�m/��ů��D�4���I��ZҿS�=��r�$/$�������LN�,���$4ͺ��^�޲^X'E�����e�OǔS��qFR�Qx.��[&��W�������G�x=����j�@�D=�7 ��j��h魏�o�SG�m��_��$BvK��[e��x�P:�s�w$��QР�wA��I�]��)�:�� ����Fo�SZ���FB�oZU �pWzf�Z��k�Iz�s�͋{��+�����i�@Mu��;l�lm��QG�� Q��@!]=?�8	�u�T�hT����Ns�,t.��_i?�w�$:Z�&'�;�X^�9={�`�	JAV�c����<�����)�{�Z�q�g8�ю>-FK�P2<!�S��;Q�_Γd":�J9B�.W�o6�U�qMɹua��;�Sw��z�q��|�� 2b��Tʒ4�_���t�H��~����A��j��g8U���-ۥ���Fkj��P������{�w���js9�rE��l��M���X�����S�FM��P�����M��J�t4t�/^�
> �F�<f����c9��/�6�q�
��/ԅf�<�B:����ւ,X��1e��r�櫓t0rlb���W�R��:�0@����q�63dn&���Mt���Z:��$�*d�3��͠�x��N����Y,�:��7�nYb�y�H|�����|�k+t����y����	�9���M=q�%F��\�XU�rUͭ�,��ٔGT��R(��~J����٦S�?�����Ql�|��QϣY��cZ-�I�@"l�5ѻ�/"�_)������J!]��f������PY��0�Wz�AI_��M�)'��W$���yv���� 7J�B�bF��9|'�I次n���zh��=��mU�F����t{��Y�]�<��1�&��^��u==���A��UaA�ޫ5��)����lY����-���7�����H+�}>�6D�:�%�B���;)tj]��2��g�������kxBPX:N�J�	}S36I)	ŕ�~Z�v����c�p��ʍ$�Jn$e�5�<�y�4��gy%�@t����}oAkc)�
-��h�<%ANv��L��!-5B,�./�����x��HnU}`~-�zfLD2����#O�tl ��`��i��g�'Q��7�5������ˆ}韙�m&Z�Α�͊�H�U��@���Ov�k�E�������������\�TG�Л�@��;�|�3��B+�j�r�̪�خ�5�3V���_A�F'�l�Me_T��ɨ���1�>���^N��`�cdDz����[R�k܃��u��A��ȡ|���h��0Vj�pm� �Ģ����4���)���uTd��dr:_�5�d?�S=�=�օ�/j -��ۭ�S!m�w�Y� 1>>*�b$�b��	'w��J�sB�(Ns7������T�B�<4�7� ��z�åK'��S���^Z�gR<�%ƍ�^�@�B�ϵ�Ig�#�ݐb�SEi��@F��	�1ۿ�,E0�N����ی9�k��Svy�B=��Iȣ� 6uQ��P�o\a�&kW���g q��a��o0�����0!w�+�s��k�9x�)t�[^f�Ҋ����PȧȥĐc��:���e��>M�U-��̘��F����9�T4ρ9�X-ټf�D����`�c�(x�ot�:��ķ׎�*��m��<�"Fe��� yp�h��1��AAz7�w<9�$^�#m.M\V��$�)���Y�/'>��hd*NsxĶ*K<�"F#w�V���� �)􈨫͎����P��/��)�5�[͜����IB/����I���S���8��#?���*5��E���ww0kSL8��5z�4}������	%b��Ѳ'Cy��0��T�vſP��t
\&���;�M����U�S̥�rR
ۼ�d(�Te$�}ƪk�q��L�i�M�˵�;���z�P�.���~_l,9�.���q;�dx&�+��d�ؽZ�1��[���/�����V��VbZ7킟IأQ�~L�2�j��s�iG�6���2�a2P��a��T�� �v��Nߡ߿��N"IL�٪�a��
�dbr�Q�h�].*L��:�i-�S�cgM�K�?�I�sH^9���>;\S�<�+�c/4��	~�A!��{���N�3���"��/g�,��}{�R�`�<̓.Gʻ�4f��~�b��A��%?�.�D�킌��y����6R|$;6�;�P�+A�ҟf<(R��yPv�?|��^U��g�,[��-�ۨ��ƨDm%��CIǛ̫uj5�Sb��s����.9���vZ���'u���^s�q��r�z����q�t�����	N�(���Q���������%1'(Ģ+�ݨ�9���������Tb(�s���4i�����N�ʒ	�a������P��U�*���e@n�y[���'lj[����i�֕����_X�X@����N4N�a(i'�.!	(^W��b6�=������(I�R�����?�]W@KJVm �N��N�^�P��{u�0F�h��[���S���ј^YE:����Q�Nl�<ܫqUh�5��]u��jO.B�,����|,�6��ceC�J�\��4�<[Z��3�EN�Z���#���L��k��j2�~#)�)#B�W+��Y�R֜� �~��bU.��AP�1�����H�q��1�9W6=q�Y"�R��J遥��#��̛���B1tJQr����5䳆?�'&����inRąs� _V�4b��&>)�q��>S�;G�\�NM�2P׃Xϕ�|QP�҇��	>�V3���J�V�qk���
��n�ye����^a�
�����������'����Z�F��i9k��̙-:F#v���E���#�����ܜ\zO�c��y Y�ݣ���gh.5�Q$���j�̗�s��ѫ�q����a,iR8��9O��b��$˘#�[��L����7�M�o���&� �^��!+���D{UV�<�J?\ ӧ�"s^�G+G��w
+��S�%ˍ�5>��hj��jJy`x��=]\�g�zޭȅ���~�AC�^=t�;@���V�t�_X)�o�kzZ��;�
�|$�����ވȣ[�w=�&YV��*�^�6ߏ9�����`�c�Њ�,�r|��#�3��I�\��}�� �	l���h(򽮓��}�0�<j��q�����#G�j�h:����7T�2Z��:���GT o\��PK{%����Jc��e�r	���"NN��h$"/����*�+������E$�����J5W��e�K�}N��,���V��CK�<��,�l�0�%�Z:s��#�� ��uX{V�Z2����I]�	#L=���e���D�a��z?�*_��8��.	���BgL�I͹��=��W��x�za��*V�Z�*��)&�:����;��1tH��]���Ow�g -���G ?���0�!i��;;�~��.��b /��Y�l)��,��˯`�bf6�!�V_
��
\\y�YDᾒl��Ə�	&���Er�����c��|D����s��u��1��-O���:n��})�ӮҾ�� G��S��_��b��1�+A��1� >��/d/J��d���)��g
S��Ջ�J,�꫐Dc�������r�`BP���]�����}��/������.��z�c�I0��F�I�������_�~���t�Ac�P�)�0�r���D��� ^fT�p}��PWGs���A���nC�T���<�hLy�9�)�
���+�M��W�>8z2]�ь�>�2�W���JJ9�B���*���3z���O������_n�\��^�����aI'����2*�G�� i2Y}N��e���N���z�G�Q�����U�Y[���'y�@�7��Ͽ:�����m͓k��2��;}'�K�W���C���������_�r�P���^˝S��&5u��4MQ~��.�"k�4˕w�Β	3�������J�|� �p�bz��c��
�<R���j����Jׂ���{���Y����=���?��C�<�����cbq��ĝ�F~�����fGT�0�䍴	��I�U�%k��1�O�;L����;�LR����4�EeC�d������>�F,^��ܯ�1��cl����_��W6���r�N����������BbUج��b��C�嵏�-�G�~��O7���v���wP�"�X=�������<p���SZA�V��;�Y�F�Vz�o�9�%�J���u^�>/��^�j~��߿����_���nD
e^����!���������%O��֬E���v�(th�Ɗ-���G_���@z�[���)�B�`3*��B�Vn_g%&^�D[�$o|k���_�	{֒W9�{@?Y8=�~UP���YxكoM�RҗP�kr��E�)�K|B�y��6Ґ�ܴ1����,˹�`�/����v_��/����Y��}�r$a��W#`������6���>���u��,�Pv�L�����/~�7CtP�U�E����͋s���~{��o���q��Y��.�3E�M�YGb�X�g�q�3A����1EVDy�1���X;��!/>6�4/M�1��Ҡ���U�v�I`�u ��ܽ���<;�Ut9���)f�!#z�+�=���F�E��e>-2�۝��H���1��q�rnUz�ئ�6Z2u)�>�X 's)�|凴|�dٞ̽<�d��&������x�O�^$��$o� ��#KB��@���.�GzKA0�V�V0�Ǐ_���{��,
����=-a
�G��P[/zG�G��O���������J�C�֭�2��_n��o�cuZ�֜h'�ڡ_[�"�Jك�^�� G����,�虫�8X_H4.�RU��W��D
q)������2���|=f���pA�$����_2K�d�5M1=���S�Fk}E	��O�MJ=���m��/�t��TW�q�}�ûZ�̛��8�G�S8MOY�&����v��S�q�w�  Փ>!(�A�O+/[V5�����śk��O�O��E!����ke�L$]����K�37ot�?)��͝�oH)�b1*ʾ_V)��NO|0�0������$fH&;����Ru�^)�#�2 _���,���C-�*��.��43u�
��"#��C��b�-���]�+�d���Z���;IZ�N|�u��<�GZ������鈈:фH�ZơC���p�.���� ��&�	�m\����䊩��b��N�W�%�t�W��"�fA3~�	���FJeP�S��Զ����yW��T,�c���l�g�GW4�|���c+'�F�(�D�e�y:����8�yH1Q��|��L@)��T-�E#�	����K� z�ٲ��E9.!2��y��?ۺ�w�j�k��w�j�p��8Ǖw�ⱟ�˚����u}Ʊ^�~��W�M�k٘�By�Ea�.[�������in])��@	�F�vh5е\�FZ��Nd���Ô< ?����/��H�l��Z����n�/��k~�g�닾��Q���A]���ml(6K%ZJ� �{��1@i�y��j��G{�����SZU){��^g��Z�vo�k��iXF��Oti� �˺_r
�u��b�)�L^�
.{���G��~��K�<O��*iw�����(�ӳ!�^sV*L^�e�8+W�xr_�j���g~=ha]-Y�q��U:t�+��E�@�i�d�\�U�b�a�2�)U6�����b������+�i.�a�S��5����/�Q�\��ҹ����Z��q.���4�:9�X&�S�E�/��Q=y:��2������0�e?������*/�'�������R����Ǽ6�7���,�"m��@�X�&�^�r�S�k�u}?}z1~ēWzhșq=ɹV'�Ni*�ٿ#�خ <O.B�= {�q��k��S��>&�+��
L�P0�������^!��b�:5C}�`T@�>���XH �������,���*���<�G^�Cz2����ړ�>���T4V����Jn��T��U�/}�(�?�@��Ӟ,	�l"R��68��T%JH+��x�d�W_��>�$�\�ƍN��z���!F�Xi~0Ê	���y�*�S4x�y��$�l����2�����/&��[Ɍ�L�`K���'?���֟�~��"�軖5�C�M���J��9�q-�EVH�%��?�v֐�i����¢�T}R�0T[5��d�ύ�5c����b��?
��ZL^\�S'�o�e��5�eS����}��l�.J�	irD6R�z.h ��&�OroW�t�R�z���(I�(�2T�`�M�8�o.������q�Ǘ��R�+Xz���!���@��@ֈ�J�VƖ�$�xHd���:�]����9�B���"�pHt�ѵ�E���)UQ�	;f+A�wă
+U�>w0��� '��֥'qs7�&�R<��9ǂ�K�ə��UV�J��cb�-
h��Eۖ�H�p�sq����&M������/�S`WǸQI�e��=�p'O�\ç�A�/��(�bJ!������������(>DF6���!��+LU�ʦ.	�K��.�LL6H�v}�h�j=9`e�:f����C&|���O��G��\�GV�����{�4�\�3%�B����N��q�^����̾�d�ֆ���-<yK^�v='�%b0n3[e��j@�.1}������@QJ���d�r�8�^P{mX�&��˷g�GT�:Ivi�zR"1Fz�G�HP�GO*"����#�)́��:D�E��!�-��T�K|@��H�vx�d��O"3V�{0���"��MgBw/Y�uj	E��V~
��H���n`(�SH��l��Po�P�}j��� �}:�I��!wD��V:������_�0Scm<�xv���:���CKs!
��}5��L}C9@�.�KH�Xjʩ����%ﳩj�#��h d�&��5]i��±�S���~Ń;�(d����ϓ����AD�.�xzZ�e9l�u�|��7y���{_����.:x}�
���ZZ�*b�����9{v]���� �WG���hNx����8���Cݐ�=g*S4z���$H�S� *��
��I��r�P���!}D_�\�Y��8V#1�W8�>�R\�sf;I>prEE�
]���m\�j>��,ҕ�6BZI��І5>�sc�)���3'���$f�S���Ǯ�i�-'~L.�����8F�������]x������C��R@!K ���b�ʳ�����j?�`F��~�}��/%E㡖01�V.���`��!}|�L�^WX��aW��,5��-nP#+"�tP������Y�58Q��V��ƱN�s�����p���j>�'�F��;�e�(>6�G��X����[�t�^]��W�G����S->z�����L��6��t�'��H�0:cM�1<y
�yj��[y���iݾ�Qa��H3$	��
��5d Dۮf$q����U�OV�9��=^bu]��}�v0�Dt��v�B��\H[R3�?�T$%$���Nau�C���H��G�f��t\�J>�ϕ�k��; c"����'vP��Z�@~'��㊈!=)���Ç�_���^9Jt�_�Ly��P�'�d�)�%�θ=&�П�{h�X'�{����+t Ox@��J@����u[�ؘ�2��U��1��Y���J�(4.�\�Q�ʨ'LNu��/�U�H���%����r���ҴO��Ϝ��4���"d�1��JL6i �(叝��&�p���<��En���Mz��)���t����p��ǈb��Zv(��@�<	D�c�N�n^z���K�/��9���T[�y�� ���;"��ʞƜ�(����9�F"���@<��b�,Vj�3ՎAg�0
���,��8���ّ���6�d(k��[��O���T�oOBAg-W	x�5-�������P�xiN��4X�5~j{���S� �����Uf���ң�#�@>��>�_q�Dr�$"�/��:Q:�L=�H�_�N5�/^
�k����.'��';-����C�%pfZP$�e���#o�4R�U2��4��Qi�>ͷ�ʶn\N3��x���e?:�����ך�l[��b���JF��x��l\�@B�ww�Oqɤ#����7T_&c�]��f��d��ZD�q���4z)�t�=�3�!�}j��cD	�W�2(�bC�o�R:A;"��i���r��oQ�<�lԕ �,Y�z�u�	�:�g�dn%#��_�3��M�s�eS��i��˥zK/{4�2	(Y��K�ϓ�c��9=�`��K�|Ճ�zlA�i��js"�va����Aq�����x�ʷ��P����g�R���3�Rv�����PN҇�T�r,7(�y��v��'F������s��tI��Ͼ3����V=�t�#o�L�6�	�W�x(.d0NT@R?��{ҖK�����+��H�Y2�y+r�0^/Г|�T�o�V�트� H�
,�M���g+��y}2)U)o�YӸ*p��������P���F��W@u��;�!H��̜Ee�t_���rt�|'�XFP�>&T͛���n(���z�\)cn����AϿt�c,U�1p�"��[<�6�F)N��RK���s���S����Bj�����36��v��r&�y���no�.Wf�+��y����\k�?E���0�7���%$�_)��"W�T|�����19p��6䡰L�tW��U��EVwf�i��"Y���%��^.j{)���jISi�Bk�K�s��4��C��� ���G҉~�ƄJ�{��r?��N�hO�]rB��Ž�;�g�	4�&���mfɋ���C���]T�}%�O���R_�;�j��t]���N��|�p�4J���ʻ����u���b���~��}�n���S߲�����yg9�[��^T��u��,��gI����g�4�t,��hX���ʐʅ�;�yv�����s�z��i ����?	Q�I�]��J���8����yn
�}�Ʒʒ:ޗ�^���#)�
��7{��1X��@E@*�i����O>�T�8Љ�,���������<��������A�6�yՋ�����V#Y���Kv޺�Od����J��"����P^L��!�eL�X�Τ�sƹ�+�Cj g�� o��(;mC�1�?4���s�?{�C(|w���J 8�ձFt�/��n*�m�"o�Mx{�+�U�׋p=�d}���H��"!�z����jp�j���P8�b`}Q �Wz�w�EX�����:���͹��~��+��@���G��ˮ�6�O�u����>ݔPT��&A��x�z�t�`�=O�Pӱ�VA����
 �n�����g�މ0혲��4�A=Γ�eDH�SWCY>�6��Sz�w�n2Y̗�8L�b���'��VHKJ�䑺�,����'�br���rj��{\��	�t��u�s�Е�P���SF���S�,/f(O��i#ǔ9�M�!{W��bk�bx��չ�s9i�)�o��N�,�O%���W�J��}��G
ŤX���/�X3]^�$��i����w9���)kуm�d~��9y�AR]
;/�{�h�ԚU"YnFY����S��w�*T�Ӟ��������Q��Z��O�>FST��O���r�����ط�c��G?�B݆��p�7���4�|��,��g����tb�i%
t(����3n&V$~\������!�������4T��^0����p�G}�&i�Ľb�1J��th��([c�#��Y؁�R9�C��M.�d�}3k�̴6�sob��ֆ���SiQ��0�����yf�J�i�7��]kZy�*��A�b�<1�M�/�ks� ��)�&�r���R��Ð��GiJ�2v[d"�/�cE��O�=������=��ǵ	قd?��&�N@�(��ŲX��;�/�q������G8n@��(�=���x>�.Z�$��Zihr��r҂�JdC+�Ս~/�{7X���W��D0�h ���z��"$��*�x���˹_(�����=z��!�W�j4��'�:o*�c��Fa�
g`��?Ԗw2��2[��!�R���gJ�*��/W���4��%=�G�4)�v�q�̥��5��/�c�@��ԗ�"g���V��wdz��u�^_w�S�3��~���k�]5����0�*?���t�9�>%C,��E{�{��2��$�&A�z�����zuٮ�cl�Ϻ#�2��+A��w8 o���M��/M�p9I��N�_ٸ�,t?KF��{)��q�㍾����R�����fxF�Rw�����EbӞ�[����԰�anSl
-�U�N��V�.��pb�����n�y�>�-g�1�����H1�q�ː�"���j�=��ƌ,ԅ�M��8���GT���t�۹�(���RM�K���4ԒC����V�HJp5�n����0VX)���tF��Z���(>և�H+ 8�F����窖��g�*�o�U?k9>Ȯ��2���M^d��Lȉ���rV�Чɋ��^��%O�+V�i�(W��jҳuĐ�ґ���@��Q@���Vs)�Lw�kM'&n�m�>�;�zh�ot&A�ۓ�@��pXxR^1���6�I��G6XdM4��Oi��!�"��|��_M��2���ff��J���udBin�9�����<Y]�@��n�S'�d�c�Cn̼�^�����V��3��\�k}8�T�>���
�|��0�E �^�,@JD���F��g`�]�z��iQ�,�a����k�0'~��<�����e��ϧQ�赴���$�ɻ���O	T���B~�>^z\�������C����謔�5:�>���d��O�4�!�k��\��)��:?��:ړg�:Vr���$A{������o63=ù|��P%ZN�#0"+MW�|-|=ps��l\�@�1�Y��3��,+	`G�#y8�_��;lDwgK(��ֳ4���a1����;ZLZ�LƄb�w_1�\`�v�V�d$�h^)5ܯʹ1�A�ޤ��`{l��@<d3)"LH``3S���'��`��$�^�w5��������%�.�4$:,����g�~�X��L2�Ž{�έ��AD�%�e MY�����̊k��']y�םk�,�U)��J��[��QTyX�t��)2X��S�9_�=NS`�-�^E�_��#���/^�k���$��Gj��>U���t��I�	y5��y��/�Y �zH�˿p���"95�U�/_�[��V����#.i -X��ķGOˁT����ğ�pj�:Q�۩'V�y`�s�o�A��:�_n9�i�8�0�+t^�3y�YLd:@�AQk����f;|���pBQ��ș}�����3LtTEE���pW� #��p�w�`^d���0�o|B��%60�t.X���ޡr>��Ҝ�K+�Ҧ�X2,��R8��*^wD_�P��̔y��,��v|6?�R�;���9��79px�X{�Z���$�(�F��G�*r��5��y��a�?�-h;�L`=��]+ϊ���9�j�f��鳟�"Þ:���\���m����S�y�hjp�������2ҧݕ\6��q�@�4�7��;C�G2�6���&���?��9�������s#����+;��l$�����5��ɖ�ǝ+�Ի�<����nC`r�{	����{��tx'��������Y�V-�t�E?��n��e����z�|�X
��W{6�Y` .���E�ʀ��dc�5�
ML$��EZ�0�z���Qɇ-�(̷����P��\��W��L�d�~�E+u��D
Jw�/�y��2��E�q9GV�R�#|M�Ц�m:L�(�;���>�<�+�B�3XG��h�r/,�}g�-�t*-�j2�v�b���픭�S�y1.k eh룍�-�G]!"���#��)b�ۖ�XN�-�0�M�do�0�aCxe�%`�l��<�ICҝ�Bn�(��8�	���^qi��y���Q��\��%*-/)]u��-��������E�>��ƺZ�P�]��ս>#��;+�q�F�hG�4��L�(�\��Qz֛WFJ�&6�ǲ��q,�=��;�z��4�8����7m�}��g����+OBm��Ű\����* O��S_^Vm|��s(pҫ�h�g�ͭڳ�C>F+��`��×��u��#^jQ���d��0��h��|����B�zl_��%��Ȩ�x'�w���Ψ�����O�[�ʕ�ˮrq�;_����-�f;���^��}-��(B����}M��i���}d�U�k�$ Fy�8���a�Q6���C�h^	b<^�@���1T�V��XM��(�#no�!7x�+N��z��0��]��j����[鮁��xIيF�{�r�N)��G�z��.7��7��H�+���⯁J��� ���Ĝ97z��
m1J�WD����V��j�aI�Ut:b����4���2#�.���>��6����h�#+k��[�fU�E�U�FM��u��#��Ɍp��zx�*���2����[Z���r�.������gPt 8�]�;mwi�҂p���d�lx�=@��+Gg�_�Կ����L�?�s<V(51�,|��K
r���EYK)֜>h�`A%i/�����Q�e+�\�Ah��2�m���SH�e���]�À�\�����L�(����K'��x�g�Rh�䭖#k�xo�Sn�g�*�<$XN����؃�7���e���M��,����e�sr���W^@Hm�C<R?�ϔV8 �a��[X]�jaŧ{���q�J�ǰ����L�d����'�+��m)�i��t����g��Q�J�4�<'�����8��̜�9���j����9��:Ǟ1� �����̽_(��D=έ��ũx���V�F'ሢ`��YE��j@����(H]��[Kh�L��7���¨U�[>��=>����gi�wv��z67[y��0�}l��2����*hcs0{ f�X֯�I[)�+����ʞ��B�m�Y���%v���p���^+K���\"�9v��o_1�唱x�$����.��ٔ՞�ι�>5vy��x<8n��ey�����Q��b�_�՚}�����^M��p���A�[t���|�ׁ'-�������v�8#�U��g���U+ ����Q�ǳf~�<\�@2�
p��g�w�պ���q���Q>�	�̰��]��G׊�A:��z��3�L��#��К$S�44Kj�.d��f��W���������-����J{��~~�.C:C�ȒԳ6�&v����a�F�sn����T�����ս�����@���ls��ڏxumW?u��`^i�ʁly�����q���X�ɯ7�����U�>҅�q�0�ݬ�,�7�>��8ɠ�}��)�=�Go䬕�ϑ�s3,�c˖>g�/ːz��1���5������YsZ��vz+�x��m�Ci�R�1�v��cq�+~+�)/'�;L�v�8d4ųq{�RU:>���8JZ��C����&U��@Z;�w���5�+;����4���{����q�Z(z�R�My��^�����;4��ӳ~�sb,|��c��Z��`G"/�pl9Z��㦐�d	C):گV���K{)J�m{�1����=��_t�^F�vRfi~C�>�d{���Q�x�X�m�U�Qޥ��v�RHwZ�wg��oa i���L<��-���n��8�ܟ��H�Ñ	�'�̫hN����Y�3頋�H��;�݃�Wh@�{�W�ud9㥙�b���j{	���Lq����$v��Lzt�-І�Q�d�q��r�\-,�r_�sC������@�dm��r+|����2~�#�	W��J�ª5.�� �)�
�wu�t�B��{:��Sb�|3���~�⁧[�?�!PxR�)���5/���ţ�ҁEz�K+m���({�H��<ܽ���m\t䠍wA���p(l+����Ġ�.o'���E�3�\���e��]�H�����K�����a��kW��1�QzK��\��.�9i�醧��N_�V�G�V2���6]D�ʓ,�5��� �����%ݱ�u���O�k`u&������goU�}�K���!��@�����A�XO�y%�噳n�@��q�Le �4`+���\\����}��E�I�{b�u
��D���?�J`���P�%�u6��X�yWcLhwW��A�ZH�=2�e���򹚳�LƩ�'�4�ˑ�D4�`�ޛbA���A����P����}�����R�}"O��ϓ�u���G����zR����1Fs�kY> �bX�:�<Ke����H�)밢#Q�rqT��m�� Q�B���@����`����>Ih�]�O��+�o�?`��Bo����y�;ןEg���άH��t{���֫����|(7c�5�=%�+5�f���}ytJ��'u�����/*��Ծ3���H�����!�2/e(��|N"�#�c��^xqX�`g:/y��Kqx-�5����Qʮ��-<���ފ!�n�k�P{����ˠ�#l���ƻ��^8۪���~�������@��}%�ge	 �<��"�7���a����aQ<;�����CUN�
�����O���j�k����^�~�Q��4���yTυPVJ���#ڱܒ�Tzf7��C�F�c�̗#�vS�}�M��v9�%/|�7/��#D�Z���2;���i-�Wj\�6�w|#�s0OS�TgM���Oȴ��`�t���oe q���q�����H>���������i���7��'9mDI!�8�[�s#�l��iê�O௞�D��,��nO94���������Z6��Bt�<[���Z�8D��k��C� �P��;�F�Q�b^ƹ�nw��Ґp����)�R;;�C��Ŀ#�k�u�@<��ra~\�*2v�*�Sβr-<>p<R�qkx���A�-ꁟ�4&#�G�6�von��r,�S��3͹/���?�>�ц���N���`��r�f4�+igJ��*G�+30z���W���Z#>����	�8}�5=CM\���sE�o�L��e ��Z�݃��_WD.��#�H\	䱑@�~Dp�q��[��I��O0'5=�a��5#����3�B�x�U�੝�w��K��MN?V.�ĆYgz�|jh�7k���C��2���;*9y�����{Vp��C�C:��Y8?�%�T-�%p���'э��+4�xqԵx.>m��u�[�nK�g�����R�'@�[�("S6�V��@��rГqP�h����	�o��c�*��q��1����A�t�~4��w~u���#_�Cm�;q�_�@j�&�����	�����R��p>n�/Pc���+ͬ� �բ���g�� =J{��IL������=W*{���+�ۗ��ݞ.,=k~k��m*��k�@F�"����o2�@��������X�4Ȝ��{�3~�l|7�;&oj �G��$x�)A�F�+E�Vu�p��j�œ��?^�|Fy
?Y���1��vso�i�z�[h��`+����c,)�G�
|�aE-��`��H^{�Y�~S��x����R��K���I������1~�T�ժ���`��کn�>G���������+8��m-�",wJ^�3��w߆@�%3d�.�*R�v��؊�1��������Q���D*>��96t��-תz�+6�6�8:���tm���D��tkA��~������X�Q���Y�b�����3��t�|n���aHI��Q;����ϛ�n�KH&���P�6[�|'��a�u'|��e�� n=s6=��C8`�ڶ+���/	�g{��`�B?���f:˳��)z�sc���N�ἏS��c� �ְ!>P��m����[�)����7
�8��$���s_s�΂�p��e,/k	7-}��^����2`��EpzWjo�����y-P@�8�; l�-cCB��[�;�l�>���.l�؈�2��&v����3�Y|-h�G��]@��҃tz]�0�{��@�9����O{�+`X�T�C��b-��G0Su��{�H��ƞ8�ia�=�R��YX�l� �Z1�}��̔�!{�'oz\U��e���<����}��ڍ������e8eN\I2���B9"7up���+�S:� ��u����)W]Ŧ�x3�� ;��"|��R��g�8۩�/i�V����������-z������5Johu������w0~_���8�*4���'���n�ǵ~R����.�����.Ԥ�9�@9%/����ƫ��ob ��gbo���s�IIg�[��.ͼi%��?E���G^�&������Ap��[�@�k���А��� �=ZJ�,�O�}Q^=»>�RΜ����+��\���{��5�w�宀�2�n��L���L�l��PW�_o�e4�i�}��[���#�{ ��֊K���Ûy��CB�J$��U�`g.`������°w���<����I��&E۵� �W���p�ܸ��� �M�+T_��0����k����a;�g��[AWg}u���_�m�w���>��[/%^��O(��q��5)}����8b��R���ӽ�֧����~7���I�82�o^ג�C�Jy�O�%�� g%y�r��/��IwO��}��*��I��;���#^l4V��p�
R���]!�I��d�|�6��(/��JO�KH���w�9_�Y�����LC�$]�t�K*>�H�j� ��<��q���
�>K�b�5	��n<Ң�����ħ ۸����l�G>��?��;.��X���"7�!0sC�JcL��|j^qV��;}DM��m��
W\9ӫm�-���$�>���W�@��Ԡh��e#��}���Y^�i�h�^Fg�X]X��b8��'o�ǣ���[Kj?��E��O�<�}g"S���<U�W�'>� y�
D�>+��n�9c"{<���BT_��~���b%��+��qg�v�pg��?��·t��$�gw.i �b|�=���_�UKLT|��/=ш�$��/N�㫳�z��:��~+�A�+KpO���F5I��+��Z��,���S��yd�V�C�@�PKs��lz\?�HB�q&E:}���c�R���EX� �����Zq:<��H�uP�En��΄�{+����O&?1�e��]//��Սף%Gb�{i�����;��Z��I��X�:�]V;��#�>J� Q��]������|��R{�eivv0�����s�trА]}z��į�ܽI�y���������C�Gzd�����ęΡ75��D�^N�'�u�[7���j�Ua
�R�Hw3���Wa��  gx�y��n��O�G/�H�q��CV��k����n�}�����]9_���� ; �(F�C�:��춾���/��w��-:���(�}�k�ŷ0��dK�V=
���}�g��q����'�]iO]/]g�x��s˗�_�Yw�B��":h�PX�����7eQb��?�}@z��-�#�)]g-ۚ��b���E���zo$M���QحiP���=
��0;+��X:_dcf�SƳK)�@�k��+��l��
�S*����'ZJ:��^�ҡ";��U���T�~�^��8�6���$��;����:TB-FVVdL�� �0��Iv�y ��f\4x���%!n��o�v���@CU0�)�-K�� ���
�gV�bá���_��5@%�pE�ɥ�k���C*W�Ϭ��ě�Dlr�W�1{����q:�\#�:+k0�*�s��L=�th�NSӳ�O<y5�R:��A�SZ��.�,�hwI��k�\�`�"��o�X�R��?��tԲ�l/��7H>����8��#H�V3j��7�k�1#�$X�_+3��?CY���L��ܹ�֫x-��)��?~��hlαm~m�z|/���)�{�0{�0�kpe9ׂ���s��KJ�X�s1ɧ�<�1���{����c�t���v�t��g�}~�Y���̺�u��ϸg�m��X�� ��@���;Ă�b��l�d`���X�B� �kcy[43̌ml�=�ޭ�VfFdDd䏪S�:���}頻�̬���������S��X��I���J�D|��+{3H���ok�%�~u�)$�l�4�i-�Cc��9!�_�yy�a��0����#YN��E+�j���1Q[,Ԁ�����,��ky�������ц�D��Rm�����87i�ؚc��L�st�p�R��꥿����%�:�##�����f���Ez H� ��X�~��f�5��@��M���(m�pE�g�B��FV/�p���+*���%)�Q!Y�[�{��=?�u�$D6�\�#nĄ8�S���j�M�6ۢ�Fw��G���9ܳ���e(��ZgB8v���Õ�3o��p��m{nO�(�69�9�C`���qg<�[�w&��<��.����לA�qt=?O�'ҥ��=�4�6�X�q/ST�`�8g�s �se��Q�5��đj�^�Y�ڵ�*]H'�^%��й���к�ui�20�[iv�g�ȸ��k��-�q`{�%W0^���t���y��k덕��䮱i8E@]�{�K�D�(d�����1�FX^��%�GӁ���0�Z8�zx�z�㮠��j�F���]/୽���� #�4tBW$�@�/f�&�ka��{����{��Q�z����8:Z��!����Nmޚױ�W|{V���V���j�޶���0w���T^4F�(K~>T=���5���2����樶2���˰�k���W��V�ca���q?K�Q�z����^�Z�/��f���.^��-2T��H���#��Yy/�T1�kd|:� ]vjD���z��w(4�I/B�Ӭ9P!�)��L��^;��݆]����������B/H����<g*�}���^H��b%f�>w��5Hq��vi����{���<0C��}�*����{�3�t�+I�g`7E~a2�1S���b�Oӽ��i�=��ȻJ��fU�j����ج�+C��!����F�1�
2g�p^��P��
E3e`v?I`յ��f�Pk=n�,#�|��i�k.g 	�R�ٴ4=��=��4��g'�O�=��
&$<wrV��q"'c��y�T��C�10���w%�1��p#�
a��2��E��cǋ���H����%{�'���cp� ����d�ܣs��Y4{�ω72r�-W�@댻��m�"Ֆ\��/g EO�Gc.�ñ�@N7���`y�_M\��I�~�Q;�������!�\4��$F!Ofw�����48\QG��3��c!h��988Ϳ,\[y��PzC��.nj���{�[�yl;\�;�N\iT ѭ��ЮZkڪ"x����SX��%m
s��dm��b�W�\a��o�ݦ�.�q3���귤�|��h���{j�.F�і��z�:ҳ�ʐzr��96C�Lj�9z^ @`�p#�K���h%���,�$�����=���\�Y���ص�9{���	6�FJ��F��T&9�B�D~,̂N_ |Ss@{gR^A��\du�D�p'�2���,��:{d�XF��=����%�����q�F��1���!�| �Q���Bhx��( ��5(���e��z�m{ץ2U~�ᰇaL����O���H3��P�F��EP׾������R���	R
*��t��5���JFsP�!ӈ�:�E�~#�NRR�QpJ�љr��-t�p�u<x4��>��n?ϫ�A�PB+ĈO�%���Z.c �v����(�`�1��H���f�P`��9-�\K^fI �b�<q��^�f�]�躤��୍��������&*��9�t	h�U��œ��+�zA��>)u�{�x��ӳ~s�\yt٭<X2��m��c�جSmg��0�`ȭ�|����₀�r �w�;Y�:�`���L��ƿ8�!ϲ�hhP�Y�1�$���f����%?K��\��F"�Q<��7Y_j��`~RSN�h�Q|��M��@��o,�r�/�x����e���H�G�V3��ᲈ����
�ܩj�$�s��Sτ��bt]R�Z���_@���&������V���O<	���u��ʟ��Uϫs��cK_�U�1à��6��3�$�nJ@T3|AP��Dv�EK�}��C,�nx� k|؉���<h	�6��*��o`P�Fl�j�&��p����*��6ڤB5P�'���H!�|��$9Q�W�?�m��y@AyٸL,i��h��w#��"�!WEky8.g y��(F���i$��^��[v$�Gn���L���1��>�i��`K�h"��&�4lc��1&����
!�Y��2��b�~C��.|<���2\̣�+s�;���-����|�F3m�������|}��I�eޟ=Rv��䬋�i�tI�`C�Y����>�C�OG�#�����m�,.���I�Q7��|�iFR����{� ��1}o��pYL!�����b��B0����(�f�=�}�����v��-����0�_L��p��� ��;	�-j%��ճL��eV�4Jf��ݟ���j��T����J���@E�ǌ�'r�!HT
��.ͩ��<^-��/.���h�Y뎀�6� &�ض��|&��4�p�߰�}q��EZM�C��Fk��ߵ4�J�-�!��/��E��M���tnx[Ͱ�~�깪Y��$d-GXJx�,z���{�唂��8����Sy��$��@0O˫�ͫ�e:V9�?E/�C���5�6XX�FZo)����}�/"�EV�>�����5�_�ɷ�>����n0V�JRG�^��ƪj]�g�|��I�B��)�#�v!ے��7���'�w��cu�Q������l��tg%M���;3��߫�2���F+-*J�@S>9a<������Îb[s��h��Z�+!y�s�7'!�u[3�����M�)q�ӂ���S��d��|S��@S��xI������B��M}.|�JW@��1dy7�|T�������Zc�r2숸�����Y��D�| 7�rtp��J�3h��O��H�HZ�uv�0q:T�;�}���A�e�e}	)�]Ԏj֬�ݫ�%�΄�f:'Dg�p��9�@��ƞ6��sSE�+Oa+�\l�_Ī<�I�?�<��QH|�	� ��:Ɍ�uJ;�i��bp� k[���:�Ӈ��ئ �]Wn;▸ۿq�#�Ix�w)7��m�<�is�+�5���b�L�������q
Yec�BQ��^\p?�m��h��f5
$}.n��5�'���X|�Çp��9��l�v�i{����hե]��#�0��i�m+z���	���z�82�>hP�	��9�5��$�maY*���8En���+�b��+c�W���!TI*s��z��A�`fu{$�ދ���;��B��{"�EfRYo�UqlW+�Khs��J?�q��H�Ϳ�¶a\�@�웍NC��h0�{���ۚ��^jvA'u�d��y�a;@L��a.N����b�4�=}2��e�FV��G�=���Wt�"�VUR0\^�?�&3e�+S��/�D�@�v�4H�-}�Q,^���p���0�:FΓ�k9�+�Ws~"�"�;�6E�f�o����r��_4e�VyY`��l��2y#�L�:5�A���.�携3�)�|*���m�,|k���Ѩ�F�W�׸�g'�T8 Ȉ���ɋ/�Ϝ��-D�P.��T�PT���0�}̂v�ӻ{.i �<�]R]Ni!;t�hƖ�p��U3"j5����%k��j��7�pE�oݦ̑g�f��/ܧ<�TP��#Wf����=.i�ܺ�N��(��|R���glw:�5||?9XY!tƻ�޳��YF����o����o��9���+�͕�Zgkk#��3UE~& S�U8%WT��S��+��1?֧���5��;u���v0�3�OkVn6 ������q�q
9tS��6���4ꄼq�gT�)�V�C��Ё�ܖ�}z��l��4%e"XI�x��j���~(!'�����$�2F���W5�i[��Lۉ��X�華W���$��q�0���A�U��>Ÿs�bo?���w`q�EO����Q`9N�e�0�x��,ܧ�/͋ε�n��լ�|(m2��w��)�T�P��m����TcX����v�����;��V>;@v5)HkI��W��Պ�N�6y�u[���PO�-c��;��{�p ����ĻFxKV�(<̍︵������ �=����U�am�z􂌙�<�=��������!�"5�<��7�ƙ�q9صO�ƹѱ�r1���t"6_�����?��Z݂hQ\2N���}<b]}�H���b33᐀t́�P,h�k؟�KH����(2�AɁgT�4����xv"
t�2:�O��߫17�y`��IϢ 1pij	4#��Ng*x���Y0�V�^xw	�7�X���{6�PL"�G%;)�>�ߑ-�i��;�aٺNJ�GmZ4�C��S$Q�7S�4#*�S�5lB>:�G(�۪��q-2��ۂε�E���u�e��/R�V�X�����9R��݊Ǟ1�J�F�����,/�lO�}C�W*��S����,�N�h�>������W+@�r�b"�q��`ż&&�V��V�r�b,�
P����g�x��E|n�,��L�v���0{DO%]�0`�ި�t?���s������N��e�2�Hy�,�!�{��sQ���'�[�ty}uM-���3�!]�@�4��|\{A�kj1$��H ��ם�⺄ƯL���gj�E^�ي0��<�Ӽo����c�ͽ�[`\>�r�.ox��[�t����P���>��U:��J��t�l��++��]^6�������S&�ϰ9Z�o&d��|��������63�ļ�o�s؊DV��u܄�&����t�ޖʹ��[vo����&[��aV$��������;
J�f%i��h`
E�A2�g��T%=fU��G ��g���T��^�_פ<�>�:b������vd�OK
�8p6=�<�:�:l`��ꓶ�k�_ޠͭ�ki [���/�h��+�٦��[n��b���xs>)�Ʉĝ(C"g��Ρ�t m5^Wɸ�*��O�m���:�c�D���<��6���9f(�TH�k��A	@彳�s,-��"�d��-S��E:��x�̀a�n�)�j����<�F��M�k�<�ĽРE��R/�$h����?3�cQ�!��3Hhؙ�D{A���C�!~�[�m|A���3����
aR��|j�Y�JI�[D���#)�$��w���(�L^�}ʚh#��лc�=A��b��"�#|�>�����pI�)���оl�L4�.l�;��r=��m�3�n2�� ��O�+t���8
h!*PX���1v�Pk�+T¨���}�dAڇ!�� �pO�����E�*��ľv�Z�B0TW���睞��<e�N�E��px���҄(1XH�aX�G�I+����V�.�"ˆ9���t�Yqg�ud��NP��6�n�}�y'Hl�M��iN7�SQl�s_P��4��xG�"��`'6;��Q�� �f��7�D�1�Ɔ��\7wO�M �9�~s��N�	��m��p����1�ˤ�=Ǫ�JlI�Z�ҰS�)�X�g�q�DCy�Fi9��6��+�q��c/����!��Z}�'�xΙ�n�����(�]�m+�]�=2���-�2&*�����]�@R@a��l'����V�8�QГ
�m]�;�= �Do�u�k��x�CW�{UJ%O'.�S�s �"�1���fI�ר�m��C �c"e������ҍ����.� H-��A,"SIm���6��y,����U�r/��/��:�-��>*\2m�����m�C�5x�x�VhST��7�sb�)72������W�|4�R���X�iMgh���I��}i���fH�F+�@wj�k��~c��*�$p2�d���36��qWCZ���a�i���i}�x�7�����-b��\�9��۬/)i���/��\�i���'�5�S:A�u�o��#���Y�a�k�J|D��d4�-B�.�sP.f���2�m�_NutrІ��O@��G=t�k�I'��;�o�$#�u�]�0���,>n��NZ���kjeM�f�nݾ�`�T���G���X���uSr@�ȇ'���7�a".�;r[�j�0ي���:�����`�ȃ+�Ҡ<���v���(ّ�j��77@�!�?I��J�Y.��G��|�m��
���C�X1��R4W×M���l������+��L	K�+�j���5�}lm�����l��.�c�j�@�G$	��Y����i&��������l���Ljj�{����n+	�WB2ė`(mҦ�-.� :��|S>�{N�o�2�g��QgT����l��O�5:]�=͌����$KvOEf�7o~!���qm��5�b�/�ã�Υ ��I�_��ӶW�!�یђ���7^}�Jlmv+�u9c�������c|*4e֊�a>�.�K�{�{�C��۩�I����J��3��S����pmY�����o�[(�d�x:�:�1��V�]�H\�̋�R�1��|Pt�C2Zc�g0�	ٝ����"��k�v8��	>�s�-A��g �,�5���2S���?RFa�bkAe�Z4o-"s����{�Y� ���ni�έv��e��)�م���Ҡ�( ����Zm&�6f��y݄d(\	t$����z�'㬄���t�a�Ѧ=[���8��=>]6��-���V0Lå��}��j���=wc@��ee�Y%��N�N�eE�o��׸���7�㼅5$��s��2�5xZisN8�Q����F[�&�Ц���:�&�y�� �T]H3)P6��l��~�&z�0���Ѱ�9��y�X�/��a��OPx�k��]ѮD�^0�uEE��X�7�=}�v̊3Gi�Ҷ0�-�*��)^�Q��o���{���9�9*K���Z;��h����l�G������_����5[Eb׽W���2�gg9O���;;�Y�z����
Tf��Y\��f��dG!d���pC#�; Y���&�\��W�����#r&ޘ~o�j���l��ry����Ӻܐ'��Q1g�c~ ��� �7���U��ϡ_�ͅU�k~��C�J�鸞��1�oc�|����k�^�p/^�Nax�̓%p}��+�I�g`�>��X���/=ߊT�gjW�p��8},��.��}��-����7�ͷ?�`voaBX���t?���ޏ	Tr�?X��V�ޥM����͇���o?H�s�\�!b;|�q�������v�E���_c|We�$�`���O���hG��Rߐn�
ɢ����}k2Xb��?8�-|��훰�*���ֈ���� ^�eҥa;Yi[��{y�l|;�iJV�Tʹ[@���~�3�1�����	��qN-l���M��*4���k4egT�իm��y�����&�&^��M��Q)I�?h~�����R��i�_��\Om�C�,��ș�X�n�$i�Tt��r�9!b����dh��ϖ�%��d��/��4��{�j꭛��  ��e�d��[.ė�?����E�fw�xS,á�A@~��6��N��x����|a4[�͝���J�Ş�?.��Kxߜ]�E�0E�����2gb��a��ϗ���w�&�;�����W��:�����}�ڞ����$H�!��3L������z�7������fAӦ��J7���>��Kx!%�!F�L_[�v�v&�Aj�SQ�t3u�)|��̟Z�;��^ 4k=eO��G�������C����wܦ��A�2�3αj�r/��(�*�'���{\�e`��'��}�'�䯹�(�ZS�B�����7C4����!�qIP
�F����o����G�׭<��_�Em�Ř� ��F�������~�=Q<sҰ��IaQ�f�4�U�>�A�.��=@%m{���Y� _KPҕ�#*a�s?����'���7q>�q�n�W,�)��\�X���M�0���'����l4o����_̩�=[�r_���
�������)L���}fn����UGf�-��σ�kM�4��y��ƹ��h[��� �S���_~�kmY��e����vV�w����K�!���flY#=�Q��-��Ŀq�ʀ�H7�h�������-�fs�}��f����H chu�8��c>�l�r}ޣ����v��ݒx��O_~�'�ۯ�ع��,n2��ݒې��_����w	)#���T��X2�_�<����(��������_D�/��@�΢,9����=�3��CQ���oݼ�K�\�R���
x4��J�}J�;�(M�pǚ^O�ȧ?�B��V�`Gz�4��mXaЀg��;ܹ�3�P��~�4�=*���ýy�`R��������GE��Uf���Ἴ�I�l?����[6!�wk܄�;$��mW����0X��s;G��Cj��(k�l�Қ|V�[�z2�q�Y�܁��w����)����[��ے�����	�7�����@[A�v��JLa<��a���������	��(�C��Ū��H�|�*3��J�����}�0`Z�^(��Dvw������� ���7�w%6�Ю���<�����`D�)�ɼ��mv�'�:��خ?�3e���Jqu��8�g�#���u�U�xO:�����6""Uo�lkp��L��n1�6����o�	�J��d3tEm>�+�u*�ы akxs�w~��s���6C;l~0Ю��>3��_�h��M�&Ib���-d@�YfEgϙ+o�K���$���Un(A�r��.EX]j�ͩB>���t����M���O�p�-<ƣ�\��F�ڊW�ާ{a�ds Y\&�A�1�M��굫��e�=�=m�7�������pPZw$�o,�����o�:��m�Kڌ ��>���>�Hb���6]����h��Hj��1�o�צ���f\��k!ީ<�+�2�v���kN�U�/3[�ɕcO�am��5��Mq^ ���$bVH�&Ic<�����[r{��^Rm}�7���j�F7�*�]��b2F�1��P|��5�~�O��d�Up<2dx�y�[�e��W�ei�����<����B���p�1��TL� ��9��Jh0e S"$�4�v�~c������4�3���aK�6�� ö��+�	���_����0�5�Ժ�[7�8��^�����8s�(s� ��4�\C	X\��e�K]+쪍����6�66�C2����$���#'
� Ƀ7Q.5��(��z`Y��k_�A�_/ׯv@�;pF�*�: ���
�1�d&T�N���8Ho#��oOۦ�z�۔ü. �xb8}���[���̟�YcRxzӻ1!K���l4�����Z�V���w���.W���<׬���-x��hܘ`Rd�%�6�����F_�Z�^�����X��s���ؾ�=�����C�Ŀ4[Ǐ�BV�������*8���ɨ_C�,�g�22�\��k߉���8h������=�:��B��B��.�9�������k'���(
i|dFȆ���A�iJ;��_F�����zO����c(Tҁ���h��j?�iŚ����|P���I���Ĉ�M��6�Bܧ�	�A�a�2t&��f�I����}N:���J#�`������F�Z|	�$�v���:�iu)��nѺBo>�n���s���=^��1��ñʞ'yZ-L0��52pF��	��z�wZ����o�3���н3Q����s����<���޾��6����3I��5� �T��|v�`Q%��IS���,�^G�:p��u�	����6�i>���KN�w�Z�x��t{tj9�ܗ&[���6�[c#a{5hf���Ĵޝ�B=V&xSZ̝�|��בY�:�"OD�2�J� VD���MpAe�r�wC\D��/w�vp��
rSķ��) yjy��P��X���&�g@^��$�!����f]9�� (w9$cI/�;���Π5Ft�es5c�H�a
l2��C���R�("���@�z�M��k�`�bP,h�oEI���4�ؽv�x��7+}��>ˤ(ˡ�>��wh2����i��jt����8-�pL�y(�a�R[#��0�$�x�	���87��&#�fK0u�J��YUf�֠wiſ8n��5�ux_�HS�}G_ҙ|ɡ󆡶�G��k\g��<X߱��9�b=���d1��%b�RZ�l�eSŞ2���/V���37�M��3ͧY��Wv�*D$���<%��ҩ�ͳ*G����5��6�F�i��w?%Irdn��sR�ل�I�W�D�&�iY�����3E�Ɉ���7��d�ѥ��n 
�~y�:���H[S�/Q���4�B]�'��x"ƚ�:pBʫ�y�v�A�S$�(N�[�*
��-�6���}��g���Ly�����f�Fڗ����.���	���-@�ΰ)�g�R�<F��ƾ�-D|
� :��iP���+O��;g�;��4$�wB-��9�@�'8���1���Q�!Y	%C�s����٤t��؞�i�p�Mnl���-*�f׷�/ME��;���F6x�n>Й��V�r�����K�4�	�l��5V�ݜ�rZ��������=���!�����:���Ί�A�$Y�&����_��q_���`{���MQe��G�5��`Qb�S�v-|�F�������e���u+����J/�G� s�v����|C+qV!&A�*�IrWcD��T*��e>� ��*�?ب��y�O����x4�YD��i-7�y�v���K/{� �����뀡�(�=<�P����ޟ�j���є�>6<_D��,)�dL�z�IU��AP�1b�;g_�~�+"����P�-�!�E��")�*������p�[�'e�O�#0����^7���H:�83���Jf�%{� 	
3���S�-�~ϴO�U����"^�#[�Y�v'�Ћ�Y��N�ۭg|F�M������܍���g���,A�*E�p�.�!ߵEw	���*i�hVT�n��`�l�Z0�Y\�E#A�{"�رv���W�>�3	^D4������'��h}T0��u���]��a���օfo�I�|���0E���|�x(������$r�:~�2H�4[��ٖ&���tw�� �~�L�(�=_�f����a��Do�����h�i��:�$��+6��9e��B���q@0��Ya'Y)��NK��F\��J_��Y���8�9&r�3�:>��gi���X���M�c\�瞆�H��!h~����"�h[u�������r�_��1ԣF�0������rA)f����}�.�T�Q�� J����}2|��Q
�v�Gu��
�c�ԿH�)�IG�� �T��
ꊏ��bLwF\�� �(SP�gD�Gւ;=z���o�^>)�-���cxv-4�x�0?��ޫ)r��P�h�`�H�S�o�r�Q�"[_虡m���]ۗ Ґ�3�!@㌜�~5E���r�k��	�g��f4�����3mg��� �ƫ
"��?�q�\yq])@�뢩V��[ �5rb4��%��V5�-Rc�	��u643���B���HE�TmKL"�x�?���3͊I��:4��	�W*u���a/������*/�	�i7�[&��.aB��yiohv�N��E;78{\B�	���Y�w���Lʨ��y����_���S�)�&d��C]\��6uӒ��Z�o�Ep�v���U}�M��
<K�^{���N����V��)�����~��ָ����;x�0�X(�.?>9JA�aش�{�����|��v�<qW��Q6M��^�`�
���*���ږ�\~���Q�!G�4�#�D������f�T�.m q~���0��
�U��Ȼ:�/�p"1��pahZ�=#����+�uR�*�v�՞��/L�Z��4��^��O�:���KdX��v˷\�_>�-�J�"��M��n�C�-�o ����,��1㟤�YJ�ksz�cH���ˬ��r�vp�2o�cS=/n��L�zF��xա�1-I�6�O���s�
GJT�/Y�f�r(=�m��r��oz:��{�|�IsEz�F��!�k8p�wU��d(��8m����6BVU�#g���޵ֶ��k㽣<����҆1�
�{��A���+��+���e/�?�{������_Hڌ�3&i�
Z��UP�mh�� \�-�����2K�7=����i����,L�@��BI��@�k��mhy��{]eL_C,#li���`�����&��yV�f����j7*�s��u!5��W(�١�Lw��p�T�X@�hmɷ/���hV���ߣ�ÝW��^>'Bo~�4�c$J4����n����P'Tٳ����v�����׏i}��{y��C!.ucr?�.����l��>�ې`���qD��[EĢ���1�h�_��д���Q�&��v�Վ�����N����зZg.]���3�-�r�m[�	7H#��00���]�=�x]�!.���E�>��<�p���%��Q��æK�&&�*h�m nߏ���-�L���H},w8�GQ������C���'��6�4-�va��%$��!���01'�q-]�qǻ"g�6t/g��=�Ŗe�J�����'��S������#�ғ�g�m�l�ْ����0õhyp��Ad�J=�/�� �7�҇�z�Q���wfN�pT�;��;��ۦ�kP(�\%In�Q�V`�:�!S	F���r��W� ac?�1�����¤~`_,�7���Il�cZk-�jT��t9{�W1@kG�߶�5��?���ԎԽ@�E���/�;ܨ �sצI5���^��/�m���z�t�qN碠����ta<��zC����m�_.�S�뚯a߻2�a�<�' �_b�����n�.x�����q>�u��V�C�5<��
X��Kb���%l�,v-�8ؖ��x�x`)�r��gq�o����ZU�Na[�K(��sU�~�����sj�>]s�Ef���ȄWg�j�z~3c�ă�^�%
��J����$|v4��5KΉ˫j��Y�E� v����^��A������+��:�ʻw�O�o����L[�r�]�9��-��l��u{&i�u'����` L�Pz�����w��@�p� ^y��]�6�rlS���:��J͟L�x�LA;]52�gUXu�����Nz��.�8�r��k�<t������sc_e;�(�j.꜑��|k,��EJ��a�}n����R�S<_JV:���u�@*���9ҁT/_<�G�;�'�ez��i=dڧbc��#־#do�"W}������d����8�(|��#�Q���*N\w���~>�	�/�4;����~r'T]��Իg�5�jxX^'�ee�o����)���"��[�\u-�e���=�a��:׫˟y-ό�Z+ ������^<���TW����_�;Q;R*k���z��P��!Θj� qG�����LŘ8h%x`�K�g�0��~���V=��qV㇒5�-�Z(Ş��p�����7;�O�A�s� ��}�!��'vQ7�o�<>���)��C�	�g�'W�e�eZ��yYFJW��x�ȳY����|��S�Ow�Ģ���%=>�]�E�C�k���p��|عp�(�w����u�/E#,u���Y�=z�^�xeN5Ӵe,��a��?/j m���`�ڙ#'t�IK�?��s��ء��,⮱��܁�;���ք�6󒡣�B��3�9k�}���ݯæ�K��v���U��CUMc�B��yV6���_G�Ta9'vi�\��0�|g���\�p�����K������R�˙��਽x=��)*�����Ō�Õ�~s%�9�yG���i��1��O�͙u]~���V����S��n��n�������g��N1��5z{}��"-��������"��G�����րBu"���ְ������4�)�{.^�@ڀJI����i�̾��8#%wW��q���{��۲�3�֨��Ze��p�p��l��˺�8���Tu(=2<���w�kyŪt\��@8\�F�+�k��=Ҧum�I`Ve0��� uQ��X��+�sT}����������B3w��!HF2�y {q�p^fl4�U�1���Wu�}*F�5)���gK�V��'���j��bX��/@�Ն��Rߨa��KaЖq���lVmm#�\7���a`EdKE��j9B�h���=���N�V��܂-��$�������(C�����F��-�S9�c6f��2�l5�3uJ��c��}0a%X��
ٗ~ͭd�Y�BUg�+�ɸ�w3�h\��xc@��`h����O��z��ȳc�Z0�7&q��y&`0^?Bvo{�gI�-�������p�p@c�%���"HO$��'�q�n�oF����ʥz�TZ}4�	�M*�U���u2��ZrÞ!�َg�׻�M5�ⷷ(>���U�IXc�cHѐ%'4p��C�������]���I��^����`�\Y�j�n�J�~��Η�e�Vs��X�Z=)�X]B6���<�ư8R�Pha|<�I@�����lC{j$��0�0TC6lCeh�:S�r�h�ݑ�s�.h(����閻*��_��2�M]�4�p���ƵD����Oy�dA��rEx��<d-�wBXI� �6}������_���C��ې���۽���/�N.���w�}NL!rYu��:n��"+<[�6�\�J��I����Bh���1]6	��.֓ys5�^�.V��������p�@����NkY��*�}䷖��;����!@Y��m����I�e������<����ٕ��c�ã7�XW\?��*�%��z�v��}0��v5�H¬�yQ>n<µT���ې�|Y�n�K��E����}���[��F�O0j���v�~��K?S��6@� �=��^�SMD�!�'�'�%�\�O�"e#vdd6x�0�xH8�Q�y�.�{H[�3C��
����)�V�e�rA���:_֝�]n|�����󞸤���&!���������ʺ�Ӡ�=��Ee��5q�q�F���l�	�tw2u��(^��u�A�7{����Y�&�q����^�'�3<�Y>�ψ�=b5��s��+5X~_�kZ;d����`������LYryzI�`�Y���u���������r� �_����)��:��w6��;c�<���s=�7�������n��A�K�;��	�+Z����4xX����k��&{�r~.�5�
��S~-��=c�6���ʉv��=����SukK���7�ր��&O�Tb�e���O�Lq�{Ѩ�����/��H��pp�ԎE+Ҳ�θ�ʛf��rH��h92�c�� p����6;~�[���@�m��f���3T�N�+n����/n���4�1��U�]k�����O_B�r�Ӭ�+�Aʷb���J��g���c!vm�5f� ���%$� �a\��K��R���PF��k��T��+鎗ѩ@|��Pjk��}�X%���yߨ�O�N�:V��"[�r+��s���FidT�v:��~�V#űr���_n��\#Ɋ�=��uU|��铯o�{��Q�3+%�`�ߍ�5?�E��wZ�G�%��Z����ܼ�p0z��p@�����]�<�>_E4���,Z�Xך��&������~��9��c��u��<���/pI�橪���*�T:����N����:��a	:᩼��,{=�|L�y���| y�4�4��R���R�V��5P��U��u��Q�%n^��y4���W��1�+_�)y�H�9�׎��록N���B�A���Y+m?OR���n�Q+�<s�{��Q^�Xi����hj߼?nk���=��g1���\�(6Z�3\cLT ����%����-���]�Xng�x�w���l� �!(�S�D���Tf$9w;;<ӗ}Zv��� C�Z�w�kxa���F�68Y1����!dx�*�)���0󼚂r0��[��ˮ���$0���cz�ix�U*oW�7I� �:[�j=pf~-���ї�8��z\� O������
]ޛ�G�]�蝯=y>�fU�o�S�H�<tTl̒���J\_A6v�g�=s�v�?`�?W��sםA�W�U2���=]�-
����* ûs�ّ#J�p��:Y�xwVJ�u���v���]pV�%1�qF�C���� ==��H#�l��<��+4�uհQ��z�����BO9*U�E�Kk�lU3h�R�������]|�I~���+XGǻ?#7��|��_ݣiS�"���������H����hy���J�G�t�����٘�5^�K?�[���dd$�y^�B�7/�E��rR�Owc�/�"�g5�iw��d�7�Tח�6:�)���q�����2;��7�:,t�~=[�n����6͜{�Z}<qf���Nm�\�-�&tf�'��H� ��)�qٍ3��[ޯyz��mTޜ� Р�-��p��Za�Ϟ��A�B_�e��b�t}jz8�N�N���y-k�B�A�O����H�蕬K}t-�Z�PH3��#�s*vs��u����1:8) �����.6}>���,��;Ϧ��*��޴\�{��޹Ƽ�m�Iu�g�K�z{�5�+5vcs:���������ĹS y`_�I/r�}��8��]屓9c�!<?�1<�s�5}��R��0� ?!�ă��/+a��u������́�#i[�J��R���'�};�uX��C]H�b��!��E;��('��g��
��ky�koS�I+<�-��cd���#��5�G��Հ>=X��Tު�a�uT�g4�=�C�ڧ������ �VM�23H���Y�hi���?���sz6��x�>�PCf���x���cE��~�;L�۷��lU���� O�����=���Vnܦ�����L_��@ϔ���M|%�r���h����0�
��l�/�~H���ܝn;���n�!tF��'��ٰ�5����w>~fpy�Q����pBO"��h�w��*ޑvb?.k eݱ�RӭH�F>ix�%����j��O��7���'��W�;����v�=Q�gY�e������|�%$�G;u����b��5r�%F�ҭ��0�Nͬt�ϰ:������a"�Cl{UD����1����6���?7���1h��74<q���g�V,�p�Y��M��������Ϝ������=H�ⷵt��[�4�s�>4�=^��������'���Z���|٪!�IE+��{u��|ԡ(����}/����{��(*	t}�ڲD�̦k�'L�4�����Ѷ����أۋV��L��<g����Ǚ��&hAfq��k�͕y��k���Ɠ��E1��?=��|V�b���Ń���C.��۩�O��e��EqM�m�Bν�38
?8��H��-`���m����=s'D}��hЇ���H��驶���S��jD�A�QZ@��)�/����� �p)�*�v��|v��������s0��:��*r-^�i0�ty�$��3�H�	d��̶�*�;�+|��늠�؛�m�,�׷���T���/��\�@�����. ��Ӗ0��_*Qܡ��0��[�,�zG9y��%GÄm��]�T>�%�!r{��=��R
����0����'`O\�9x�߾|>�܋a�OP`�I�5oWB�Nב,���G���F�;�]�To�E�fl��m����;�n��2<��]M��ƣ�)�ҡa��~�A�d��dLM�S�2�A){�s"iV��Ce��w�L�6,:�֗-VG�ο<FE�Qۄ�\�����dg"`MǺ~Z+��_�Pu�q\��db.i a0[8)X豗�'�w�2T�_*��H�<suⳂ�N=a�4i��(��9�AV^�)�_"�
�ܚ��\���oc&T��x}\�@r�qB1Wzzq�lA�+�.u|3��dą)��e��=F�B�����"N�v�!�֧��Yxԗ�/Ëf���MH!Ⱦ�4��s��4Fz����|�1`��k5�W�vK�ӧ<�>ȑ��{ϛ4��y��Ez����{iJ�Y��:y9^^6��Þ����,7����N��/�� �-����л�Z�f��1b���cT�6��x1(#��a�_|6�,�:zĀ����M�yаε8��A��o�qŜ<�8�������p"}j���k]����u���<\�@�]�ϋ��v��8�����Y J��>��w
���P�A	�x���7�a�*�zD'���k�������u�Ȱ���$�Q�j�y��|&1�L��T\�@
ч��o^܇+	�_It�P����ݝ:�?d����a�x)q�l0��1�����O�ٵׅև=�"֦���%v/d�Y����ai�1:���[X�����P&F�[�'�
�B��\)˳�[
����N<��7��/����e�g�M|fg��&^ Vlk�S�^�j��t9:su
��Ϟ`!]�>r�]����c�ڞ�H��z�6K�<�3��I�d�\����3�`bb��8*R��yB�kqv�_�'��Oz��*�)a�@��]='�_�4�6ɻ����{���@]�)�u݂�<	�U'�Q��T	ѧ=���y�c�n�\�q��G:�y����Q[H2C��<���2�&��:h\<����:w2x��b��r^�6E���#{zY��ϟ�)�z5V�<s'�kH���~ ���hΌ�4�<�V��88_e�MLLL�1=��c����;2��޴�J�y��yq\�@:<���aǣ��x�(���R<��4111q7XK�B�/�@
�[��$���H\�]f�R��&V���@cJ��%�T|r�_�@B����m�cr��6����MLLLLD��^QPO��~LRxM<c��%g�s���/���֕=
5��l��]��@y�� �`�g��3�t�OLLLLLLLL\�����Q���A2@�s�{��í��}2>����[��9F��ʪ�����޲����������cD：u����/i m��)��J�;̥���kn�l��=�qpꎌ#}.�5#�[�͸,j	/@m;=V�Қ�����Xx�}�&&&&&&&����[�{���4���;l���N�6c�@����4*�YJ�s���������χ�0��07nt�A�qW���6浶T<���b>��ܤ��O	�<g�&&&&&&&*H3EWӠ_�@������$��=y�P�=1U�Y{�0ڨS��J�{s<LLLLLLLؠ]�.f!����h���3|\'D֑��6+T@o�=�!�3�j�9L�jbbbbbbbbb�x))�"q�g�w��I����#:���yVi��E4Í&&&&&&&&&&��KH�C]>�H��ul���Ŏ`m�P�NB�)�Q���@�L��J)�Ŧ'&&&&&&&&�(�N�x��w�s�q�?WI���$�fqĄ��݃��{���sibbbbbbbb�	��g�1�޸��ٞ�4� :T�a���x����I�.�/w��V-���:�2����YJ���&&&&&&&&&.k}>?s�2�M�Փ/i m �`U�'�[5萶|Q����9yǄ��[xW�g��]��W�����ĵT�!����������/�[�s���K��z����/k m��$��e֎����0��7ȪL�hbbbbbbbb��h�9h<yw�]��kH;�چe:��v�i��Lb�H��OLLLLLLLLL<"����M��l���zX]�n�M�!۰<�Nw,�ڑ�z�G�׉$�L�"�_�D��k�%411111111�l�si�����M��x����/i !LÂ���
{��O�@��S�b�;�I''��J_qNrbbbbbbbb����q��{����R��ƾ���S]2nZ;�1�	4;6l���#��7111111111т���7������3���z�~yS�ř������ⶉ�_�o��|�K�&_}�}n>111111111�P\�@��iT�q�M!0�Dt�)���r��R3K��kH���{�����������d�i4MLLLL�j;��(����ϊKH >lv���߶���d���po��nM�b�"�<	���%f f�V�I�4����5L#���xw�ۇH�#k�&&&��Q����da�1�"
M
F�d?1���Cd!�������H��|�u2�N��iM��Pټ�=���� a�)܎
M�'z�nbb�ʘ3��l�*V����NAW�/<I�ث���/�	�3��c�J�Qk��i����ܘ��軭@�i,ML�jLc�߯��@�u�⹁�AgNLL�6������ع�4���jt�wx��� <4u����sO�'�3�mu�{&�_��m�D�M�	bsj�S��V�Ia�z_^���������Qu���ʭ���$���4;�x�aH�=�P2�I�7@�,���}PN�+���3Ad�Vw�s��E-i��a��>�2�g���7�O��>S�}m��~_]\gJ_��jvS�X��H�6��;�&��ow3+4Cܓ1���c�!Ȁ9c�˔'
`�<��=Oo����KVRV&6�� �&y��la��,��>�z�]^��z���I�y��r�LX��� ��p����k<�z���_8<���4���6���-��3с��O�[X�.Cq^�-�"Z#��t��w���I�<���=]��ML��᷒^�H���y�|d��A����|=��I�4��VZ��0hN1R�dI�`�|0xC���-|g9�\���E^���<ǧ;?iX���t/�O;'9�_j	樹'���C��9�(7�b<������W�[�t���N\��¯9I����=�wd:(�.~�&.Vƀ���\�@��GA� �5�����y��-mM����=p?Q�	טM|.�!v�T�bn '+]P��!�;K�k�*��_�O�d<$��є�=s��J�,��r��s+mR�Q���91�)Аuy@��3UH�g�%��� 6��^�'�a>\g���I��=/���Q��#	������#kh{�`�Ӄ��:(�^C�Q&xZ�	���x]�9� -Q! 9��~�~��$�����z�ɮ�L17q��\^�,I=�X$-�GD��a���+����G

�\VqI�׭>����R1�2�;t�^<8!Q��l�N|V��t=�ilu��Y�q��[�]=�P�*��~�Y�JS��ݖ#+�����9�EQ�W{���l� ���X�M6,~9�<|�{�(.g �I�4��J��iY�#�F�̮���N�p4T��KzM��a�]X��_RFk�W���ȍ�>:{�t��QΓ�l6F� WB�x�+�}Y�E$z�_W�Kyd����k�V�ɯ �Fw�k��{N��Q�f�4eT
O��]�z}�-�	>�U���^?e�T%��I^~C���f�z���87��v����⹕���d���F\�~ur*FnR�Xi��+�q��8���|�|�ͧ�r҆m��v�Y�H��y&����S]}U�b�<s��۫��Uu��'�K��B��-"-T?���\�;q	�@p;B6�	!�����*�=u��U�Z4�epc���̓Q��_CR�!J�ݳ(�^���i }��۶ÜO��w��%D!�~g���Lޙ�Jů�	k�^~��m��|���qB���j^�F�/[֪"�ʤ��>ϯ��

�>#��a�ܫNՖpWF�>��\x��6_,�����[퓴΍{�h�9��@'K����e��Ō�����l�KR5o���!��$ ^�j�y�kx�F�^��D`��Q��Sad��s�l�=���U}���s����N��qd�%�a���W$������� ��Q���O���q
��&H6�{h���$����tX����^��}A����{�L�t�b���Xvn�#�h:ST0��'OȺ:|���4��z���y�V���8	w�`1 }}=��\��]PQ�<ْC�|�~��Bf��tP�s/���-�3����j�Ԩ�Xj�.�kR�b��LD�J�a���XP�&�̯g ��Ĥ�0�h�@6!�ԯ�}y�J�?F�h�	u�x�ԁ��6����բ�7��gUl�gRjIBv����n�e��	���e��U_O�f������/��L��wu^��������Ҹ*��ϧ��KHڈ��J��H+���m��g�^�ȹ�&�)�J�ы{
V[<����������-q/��;1ȻԞ��qe|q�G�o׿���������R*���*����q��e~/�ԦO�g��!/�Ό5ڞ����Tޞ{�W��Q���� ��q����I%�X�VP�f3E�⓪�M��ؚ�ꎡv�u�wIC�R����T�F;�~�]x�v��d�J�e����N6V^�@��yށ�ɕpM�@��w~���*�F�Y��܈FB��N�{m�����t���@2TY�d�x���D=��p.��=�#[(��|&���;�(C;<��~6�fSxP�v��K���L	^$�Y)��#I���Q�C�P�+�=7ft-]��7��6�V>c=hFL���L�a���ق��3 �Y*}�
�
֟���-%�GGR��N��F�1�?���Jr�,�TwS.(u-�B����6��߼Up�V��u�c��j�~�[ו�ͿA$s����Y(�hޓ!|�-�����V2�eIk1�ڕ��e��?��Y����7����|�&���5���L�*R�V(e�.ΕmD��d�/����5��^�Dh���w�3#j^�/�n/F�#�.���Ӷ"6<]Lՠ_:w�}�,��/$�S>7
���bW�.%c��s)��ێ��e�k
(��F��,ǧP`�b�RGk�*:\��+d�%�4(�ޠ9sxL��b�K�udZ���\`�FI��������1��{P&jd�S�~�3GlƱPo����w�mH���d��i�+�J*��˶dł�ۋ�4�ת!gY����u<�>2�g sW�6�����v*0�H#+c���g8a�z����N�{���GG��x�лG���X����=�_��kH�ʹ;c�r�J��L�ں����E��F���L,1$]��wx��m{=���;rD��ƽ���b6A��G���鍷;�dȐ�d,��'�����>�P��έ��I���c'T�e�NoP���Df6K���S�Nkawۦ���?�d�]�,�xq��F����p� ���{��j�����D��]����g�����W��6/�ʵh�5��'Ք�.��^�[sV����H~��Ϥ�s�ei/X��<0�\mۆ�Zˮ^�A�q�H���$i>D�Btp0�Ն �/�)}M[s�s&�{[V�H���#�ڶ8w��'��E����ء�����O���v#�UEa��T~�E=G�[��=HR����a{KWk
O���X:��;��w��!�棭@�4���A�y�{{��NV���f���� �Mg�a~��\������Q�����6�X�nc.�x��3�a�8)eMf�U_9Q�$%��a�-�H�b�>*�i��!Н4RI'���4���56!z��D�)�����ʩ!��#an3���j�KS!y�;�QY�.��^S.�v�c�"��$�ǝf#���D-{s�Z�*>�!��9Z��0x��s=^WF���I֦z��-�׉o ��uj1;o�Uֳ=$�������.;}#͊��@�ls��V��
=u�1~W��\_'(r��A���H���~�,w��X9�B����Y_h�O��0s�+g��X����Wp{y��u9��B�Mc Zr�+{��j8���~��+�W4	����᫚��gM�C巕���9:q��.���1U�	�v?X7<W0���������X�������$8N|��M��^�d��`��Y�|��5D�ڤ�e��w�ܘ��'4��������{��*2*#�8Ӻ�z���4��y���D�w`'��.FZ�f�P���3���i�h6<k�aB"�ݩTG=P�V�7y�<,�U����{�:��<��O2h���R���-��<���G�-��qM�]>�)-m�Y��Fۖ@��F�%|�SB-��n������*S��^r��ԸX��e������s��c�]ь9s͖��NSy�Y�!�=0Fķ��E"�n�&R9�"V��M��-g�����o�Q[�/�����H�:�`� P�tX8�s�7!қC�u�z�M�cz݊�$|7� [I�C}l��Ϙ�@ϒb�XU�EF���3o���:f���Xߨ[�٩�	��V�1�彚Q�G0X��W3_�d�����bKѦ�fuv��u��9m6��\�e�9��χkH�$�oх�Z�#��Ǽ� Ex(Q�M�G!��Qh�
�x�����j!���#�ӳR)uD)HU�r����4򵍦�1�+�`�:`[�DR��TW�S�P��~X� |\���,����L���~�nb��
E��q�HG<;���ۨ3	0꼜��t0�I=��{���,�)��IJe�B� ��;��ō
���M��y7¤Ē�LƑW���q瓕���U~o�	
�T�h�x�W��)`��5�H�Q�t^�C�t񲡌�h��;>󌢷D3�6�t�(�U���K���Rn�b�7�@�}�z�3�ދ���9�Y�W���a�hjڬ&ݓ��b��q[�|(8��O��u�bQ}O�|<��\o���aq���t���kH\�{�� ?3QM��O�v��F��,a�bЫ����ƕ�>	VN�w֡����wUX��I�QV�& ]C>sr�2G���}C�R#o0�ɒsC��Z�[b«��:��2�g����da����@��Zq�|<�߼ݪx��tT��R�l�6Lw�������Z�{���&	���5QL�V0��q�Ir����k����+�#�C��aXu_�hۮ[#4RV��U�e`@��~�6�Z�|��v���q��C8��ؐ%���\��杳9�J�CZ3��1�gs��l��]w@�� l��x���'�6ƍ����#k��ud���tM)�{�@RL�݂b����ϋw{�(g@�h��0���ij-��4�x����<��yw}�����Zf�"��m�y�D�
E�7�<��>���=��V��*E�:P�y��VԘ�'Y��7���W6o��^�n�M�ot��𽥕F[���Rw0o���6�=&��c���hR������X�EKQ�z�d]"�B��@���GeL��{�;N9������H�tX��e+:��ca$������Q�3�\�@����?ͦ��F�\#�R2Ċ�1�\��S��a��y�9zh}J�ap�|𺶓櫁�CZ=���&�g�s֘'��b���f�@QF��ʪ$��[׽-ـ���8cjO�7��ugh��´ێk��Q�ߴp�?�KD��.��?7�/�0�E�d.�rվ�g:�m��hH��P�1^��S�6�Q������ԞԮ��,
�㧛�)Y������֘j�d���
��f0��`�<л���hS9w���M�0�=g\'Z����0�x^�+adڇ�	VXU\��C��_�A�6���C�K�af/\%^���_Qt�n�B\h,�ߙo�RD�h+?�����
�~�{L�����]�9�<�<��^B:�C�/�t�=>��e$�����ő����������>��2L�4s��S[��vg�.'�
�@�JG�G-e��!�_�iJ�f�y[��pwM��f�9/��݆�7��O���d�Q��Gb�s�1bU�Z�Xƺ�u����0k�N6�JwK���y\{�Y"\�@JDI��n��UҒ���u� $	���.���"e*W,mϻ��TXZ�~��e�}���Σ>��mxRY�bz}�;ё�ޢ#aDe�fRj�Q1L^XǢD��%}�\)�9��TR�YV|���3��إv�J"𣏕v�$a�YS����1�TU�;�9]�kvhZ�����l�`[{���rt]b��x��B�J�Z8%�t�
���b��Q<�g� d���g�D?+7c��Pj���[��B��:��5�d��:���Z^S��o�u"�ǁ�ezg~{ڱ�PL ʗ�t9������l�2wn�K>��Q�:P����
�+S��ۢ��͛���oYIh��DO�l��l�d����e�e7�J�ֶn�:�_�Y��{j��k׬���q���	�T¨Z����5��Uf��mV�-� 2(�>Z9����üZ���ܭ�P+���퉏%�T����Ґrm�P*v��1p�^�d`!�>l��s��E/WQ�AC��s��6�|}���Z^^��(�������ѯn��at\�8Z�Z�^�|KMGNG�x����h�w��c��>�*c��o�c��N�[r���/#N���u$���]���X&�	�Qa��r��l&�-��v�7�k�r�ϡ�[������ܤ��Jl�[C�n�@���e�:)���v۳.S�m�D0~=�E��$����kN�5'�~;��><Q橁wV���-�;2u�Q�g#D�Rb�+�꛼E�c�іҤ��]�H�3}�<]g��i��-��F��~��h���a��Xқ�IWK���2�Zct����0�9�%T���b�=��F�/��˨�	���T��-�60c9��m97ZN���V��<-��w�E�on��m�da��m���>(����Q37P?�uٕY����!��Fɲ�:�w�Q]mc����7��e�:����>�N�#!vT4��4 d�	��m����R²���ް#� ip|�빚�<2���ᖐ�AR�2�r�҈���||O�\<�}�>�=\���gڇ�F�v�7����.�,�L�&B��2}���Sr�g�Db��;�]|�����㾵�4
,�㳃��g`l��Y�����}Nis)��PɊ;�rR`�)������{b�_Z�.�GƒӠ��IRQj������������5f� ��#�x�d(b�r����CJխ�!S
KԩU�n��}�Tjgݦ,�U�������cL��ݹ���aq"���.i �4e=� ��/ɛ-B�6�/�X	qh��2�9��
e�y�s6O��t��U{�3� 3���8����ՖN�A��=]զ7�<�,����hY%�� ˦�y᷋�I�XALpb|5�������0��=!|φ���<ϫP�S7�.����y�.���u��k�����2o+:r-��'|�Ӗ�ddv��Z���Q%��2a,�ߨ��nm)�� �\��}�gȖb�I*	�(�TJtvB�`y�<�H��Ǭ���n�� �g�j���>Dz*��0p+"x*:S8�`�J7�Qo.7�,��������R�et��h}A�f~��7������p��<��è����a�4�����+<�gk�%�������K�dv��t���S�7��'�P*�=#c������,G(��b�b��7����H��^ Y�8(�g���FhGW���*$oa��L�3��b��^f��o�>,0�m��U��KΚA>�|�����hm�|��!S��n��T���a��C}��	O�J�	�	π�U*����(�FTx����^�^�حV������@Fmx^i�FXa���y�@�;�O�;�p)c�>]�_���QQ|d%��tP�ӘE�1zjҢw�P�,�b�;)CD#�[Z7�������]8�Jڗ�Ǒhs�;�n8��7X�"��,���k�՗4���`$ᄀfv��`83g�1��	�?�[�w+����wծ�]ׁr(	��UC�k�V���*��-T��U�Su�e�g~���~�d`$��G)�gϾ�G��j߰�R>w+�J���V����*O��K�b~�xP٦j�8b���w��Vy�g���G�Z�_�Nt�������uQ� K�}!gnRa�Қׄd�Zр�f�,�Y�&��nAoƼ>"*C��:y����i�1'y�m�� ���	�i~G�z��
?��������)B��)���س��P�$�ꂾU��,W1��	��o0���H�	���/:?���g
�l�����+<e�2���<T^L���o��.pzQ�����'�dP�)����Py6PN4�nT��ց؋��= ����rz�t��sB�h�f��u����՝�����먬��$̰e	��Y�.�b��w���&��[ee�쭲��[i�r����!Ȣ?��4�
cRsI����q6��H.H�/�h�4q�cO���{w$�j �,��^�;�y�d�wq���H-�M(G�_茗���(qC��%l�>X��΃b������(m�����B�����������w�
]P���$z�rWeF[��C���Wm���R�<>��Z��k��EY9	b/j���]��l�,��'17�s���E�m/O��מo�Ђ�ů���v(z�e���Ђd��e���-l��
��fF^aQ�(��U��fqi��ŕ�GC�c�(����%���>�:�ذB��<�����8~L�8>�o�C��4mEOR�[<k(D�����e����@��W�S��Dz-���l����:�>%���,ԗH���DdYYu�5���bM�H\�@��,�\���:(��v8К�����k\��R��W�t߷��.�w(��()�I�B�N[
�G��G��LՋ�)k�O�Zq����gd1��D�!`�M{A%h⥡�t��#�7j�_�{�W���@dIe��C�:_`�"{#Cx��~d���}�i %�#G�y�U�C���aL�T8e;�A�m�a���&r�E8������S�}���6p0_���%-Z`,h�yj�Kw�0�'A�jukܰ.��߼���y��mm�M��JF�1��A�-Y��P�e�[/�}f����r҇����/I(.�� ��tH�����]��><����B��"/I��؎�R^���Y25��#B��Q�����`$v���%pIi�nٵ��+������2X*g��!/LL��I�g�Hh�.N,���x�P�š�}e���؇#FR���9��D'=]#������X��z������V�����c����U��
`��PM'��U��ߑ�g�ى�<����a�k�}�KH{è�3��ռ�������qՖTN6=Lڜ'�����b���8ȭ�׿>�v^�z��f���#�a7��IS�Hn��� =c��ς��Z�����=�q'�4���Xf��'��БZ���t���5g�:���0�B��_�o�����~�����B-`:��O�KHP�U�yI��=yG;0��O��@^	�9w�-�L�(<�sTDK��w~� @�o�rW�5#Lb�&$Xd"f$�8aC):u�n���?�J�2#�h۽mԂ�>0>�؅z��|}jK6��X�Q����;*SwUjN������q��׃0��"�(�{���t�+|�#1ޤ��JE��@_9���>jLc9w+o0_����-e������Y���Z�z4����I��Ռ$A\H�f5�gU�T|%\�@j/�M�zލ����̨PكQ>ފ��Ť���U�۵˩)�`I�F<d!��\�=��2P��a��9�:7�1����<�J[u�����;���_A���Ե�CS���9�g���}��س����ſ����k�#�ﺃ�9�xG����b{�����.Ry�|��9:�D�P�O�%$D1��_��)$��t3n޽��h���a���3�fŵ��3��n۬<�ȶ��Mи�:��v���ο�1����ҵ�<+��THx-AS$!�����3h�Q�޺cw+ZǙ�"�������O�<�כ%��bx����^�6��y���O^�|�0�/�����?��m��W9�����[`2��~�O]�N��B���"���(m誁<
/�Yz�$V��W����YC���|���A��eO��}uFh;'@TśL[o�1��b�m���c�w^EzX�:F�;ۀB�/�coG޹�u:`�bw&x[I��%�]\,��?�2��������[�ts��C!v5liVv�M-�n7���G�d�"�Z��T�|`�����٤^^&/�J	�w�)���y��ݹ.�B�y����Y�����q^)<���5U1��R�܊[u���zӋH��O@V�Pq_CS↷ițS)���B�ὣ4#�LT����!f{�qzf#Eq+:�
�S�崂���Y���}-?���g�F����)����u�k�H�pJ@R��]]�qJ5޾��R��Y1�l˪�rF���P����3g�r5��dкG^��2�I��{�s��=Jw������:!����ԋ�!��ߜ<�E��8݉��k4�M����ϑl.t�J�G�I�]al���φ��L�oJ\t^1���3���32����O�$z�J��-�Q�F+/LFgLPB�.v�h�Y�YYJT��kT$^��yV9�s�i'h�����L+'|6�Jcw$^<
�ȇD�ڑur�k+�c d���ͬ��_���B���X�K���)P���s�.�-�v�����Ry����V�ɔ����Q�l��`��/��6C�5�J����#s2��0��En��<��C#M-_A'��urd ��
8k�-o���S��������Z���b0�VeO�������ӿ~.,���W������g8�_���{�������r��?�g�3�O����տ�+wU���;���k}$-h�?�=���S�Z��?�&�������i�{���_s/�_�����甬���o��}F���W�/��ݽ
����ι1�&��?�~�~�[�r���w�&]�����������N�����o��s��,�����O�k��?�܏����k�zҧ�3��C�|}bbbbbbb��`H�Զ_��&&&&&&&&�
���h��Az9��b311111111q���p�وW����s���ך��������8�@��0 �ꖿ��Ο� qbbbbbbbb�50�G������8z���u���������������4��i]����Ϲ�q41111111�1��	���8���j��OLLLLLLLLhL��SH����C�����!������������������~����O���������ĵ1��;�sHW¯�8n�}��6��'��&&&&&&&&&��i =s�2��_��~�!E���̹�7711111111qmL�р9t	��ᜣG ~�݇��nbbbbbbbb���ң1'���_�c���?|HQ�����?5�}bbbbbbb�E0�c�=���#���=��m�h���;�y41111111�*�ң1-����C���?xHQ�ݯ9�������������ċaH_۬�6{����S���︉����������4�&>=�?����=��u���7�MLLLLLLLL�&��4�����;��_<�������o��MLLLLLLLL�.���h���Q���/RֺF?�[yOLLLLLLL�:���h�\�o���3�����1���o9��?�&&&&&&&&&^�@z8��]�a����:���)~�w��nbbbbbbbb�s`H�����?��~xHy��~��w��&&&&&&&&&>��4�9��Çq�{ο?�8�� X���������NLLLLLL<�@z06��Av�����m&���O����׿�{�o���u��U��������~���G�o�i�~�c7q.�ҟ���7��?���_�������MLLLLLLL<�@�B����o��_��/�����o�/�����r�_���������o�����������Z1+��>��yX�^/�����0�����8�w~��{�/��/�Y���������*o�{�;!$!���Л(E�"��}����^VaW]׶�]A��{GZ���PCi$��~s&�	JI�{�����<��ܹ�7����?eee ""s��u�N��H�@Bd�� �A�V�տ�����х�����#�Ꮎ�0}��K=���F����Z�����UJ8�����Ѫ�?n��n�!p2輺;7��3.�.��4ֹec4�:��r�u �zsG��*�z�'��0 ٛ�~77'�����Q�lTM����D�M�~ݎ�'�pT��,�|�Vgu����_-���m��~]i���w�m��)�X���J@�!������ہ�<�l�NTWl�ٝ}z��6�_' 4�<%�#�ѽ=���=���e(�G�TBQU`,NΠ����#��y]�9�)�����>U�����tZ6�H���M���84�5OA�n�Cоy �X�3�B���I�OH�f������U���O��5*��i��Mv���v��^���
k#��=ʡ�.��k�e�*u�u٣�Ƈb��HM7�4V�4?�>:�{��f����0�gol����w"d\��<���D��h3�ps�����/1�~؊���^I��͆�(�E0�6$	�~��m���x�ɑ�~�|����j;����k@�d�ּ�������f'��[�w���1yAG��|0�)�n�ؼ!FrMB����|��]u �pa��h���� :;�.&�>��;�Y�SW�GE�����	�}��r���2��v��.��\��{�jr^����ϑ��pT�z]��fX�(tV�!G��A�����_�Ƣ�	�3�k���@�^��O�fP7 ��]�}��O+u�G�HO�N̑s\
Z6���j���?[��[��\VOX�Ѩ~�u���H�lG%F�&��	�}�+�N��I�b?68���LDe����56D]�:-�OMz㵱�G%~'��/~��3�5rK�Ād`�A�x���j�7G���&�߭��%��t�*O�s����߹:;�%%(N^�߭�_x'm9;Y�uc��n��٬B�=�꘎��C�h~K��؆����ql�3��m���O۱ ��db@2(����7������)ה�������G�W��󙫼|��;ڡ���N�./ �o�{]D�*�m(��<{��x�Q�j�sh�h$E�٩�YbY'�K�߆$�)TM|OOFX�>[�D�0 P�ІxqT{x���w)��&�����Z[�������kz�QJ xeLG�����3%��`�N�<"ĿpS{S�N�)�;�ѽ=1�T��k�
�tu�JXk�\�Y%�R��j�Ӆe��'�la�����NGW1f@{��۹����U�)���q�}kE\���wF/N��;7C����f�>���KœÒ�Q*~G_���^�_.�nCc���[:��������X�U�LD��V���*7�nMa#�����r�hݥ��Ĕ:1�����u���pw�X�V�g�Άv����'��)��}�ڻZ4��?flQ�Gm�I���x��Qh䉡IJH����,2B���P�pwuƛcS�𽖞���Δ`�Ό���� P	G�,��e݈���9Eذ?d{���t�.-�kY_��	�e,nk���q��1����vx�U؟Hꖬ  ��IDATY "{a@2 ы�̈d4�T��{%=O<���8z2O�������'��x]֍��~aT;<��>�mL#���:�VG4���C��ΤW�tBP>{jK|v���	&�D^Q)��� �R�=�4Ս��^{�<2ir]}��-��i��-y]փ��+�6&*�1]���ǐd[�3).�ŀ�*�����'�Z��r��'�c@ҹ��qs�P��5����_�X��*�Y�/����T?|��N��u*#�C��3I�xjx^��D�ƀ�c�2���Aڈ�Ĩn�YA��Dyd�wiC<��(ץ�(Fڈ�W��8�"C��������C*H��ᖞ���J�P��?�%;��Ȗ�tJ<؟��-<��#��m}Z`�ޓ8p��>�J���zr�����n�����H�~���q)ps��u�?9��9���0�~<\]��87���#7�ck�i�>S"[a�[��t�A�p�W֚�K�����J�Wr�]m��̓A�"O�H�_>\��rNo�+�����mY%����Gs�q������ZA"m��'�%ᩯ׃�V�tH�P�Hن��v{�V�xa���u9��m�x��w~���'�&�E���3^��M^�R�G�ё4�c�6:��v?m� �-0 ���-8$oc7v��̵�S��a5uS�f��ic�ۆ�k�x]֞�V�'���G���n��uG�vk����ze,pC�ckG��
�e���|�۞X�p�� �`�N�Չ�_bȶ�u)*^q�v"}qG_VUԚX��t�q���׆�[*9�ȶ|<0�K3^"�`@ҙ	�q
����֥�xn���T��N�f��G��y]����������A�l�Up�fM�{-���2�{s��!�%� ���$G��j�>Do���-8��*���-�	�>DC��kb��M�����o�ND������L��Puĝ����U��5Ť5$��KȾ�I�gK��T~1��F�D��G�D*SV�27'u��l��-0w�d�>yU7v���ޮo����cA��V+��5H�>�ڊ������a����t�~�jc��K\�#R���*Fvi��p�m� �Р8<��F��Y �ø=���y��b(+ڑ��$���s�Gv�7}���O�7\i���:�ߵIa�t�nsn���=���I�!�ي ������{4�1\iC��)C�&����{��p�u�� 9��ti⺼A	�$�(�~C�(Vh��:D����~D `@�41��h�#�$w���Li�I���|�>�M��P�G�?Àt��1A��$O��0�K��c�����D A�Hv!�b}�r�d��%i�I��G�����bC"��7��fi���$pM�l�1*��9��b�&1��G�  6@e��?�
�KT��rw��RN���c@������Ar��6M�[�x�tj�$�a�r҅n��CT��t�d���y1!~jg������skɎc �/$�z�6V~��^�)?�j=����RD�4����h�Ƅ4 �!�7�����	�և�G�!f>0 ��$���^p�����sz�^p����zA��w\S|8o'+���=�������H+HRT?U�,4�z!���G4r��$��V�� �hސI���ĵ: ���~vɅ���tU;�H�4��M�Ym��I�����%�I?��0�a82^����ZJ�`4�v��-6�I��H�T"�HR�HT_HRT� %�8��$E�g��Rx]VKV��bZ�����xM�O����6�~�d�V�6%G�ƪ7!��je���8��� ����R�y�]9,��Q��ڸj��&]\]��=�,vak�)�THX-Vu�]�&�ĤG�ʃߑRT��鑸_8r@��tE�Ƽg�I�A�D�?:��n���d���[���ř����$
��F�z����p����{����z.�З6�1�K��tv��E�����p,�o��D�À$���t�덕j.<�q7��rs�u�Sb��#��<�/1M�7z�G~^�-f����<	#qqq��;�qǾ_R�1 I n���W���t�-A�"7�-�1�Gb���J�sϙ �VT��2�(����	AHTOl�`Q��%6��<��ǃ��r�������^~�Z���۾��C�`��m0�� 9#�ܛ�ꋭ!���>5r�}V\]x]ꕗ��v�x�9+���?1��6 �9��w�����kVVV�(���$ow�/�~�$qseCT�\�!�l�u�W��y���zP�E;n�Kw7��/�Z���f8�����!M�JymwW�ҡ�a@��ՙQ�%B6��́G��<�����㎸;K�aFFE& ��GH)� �:����V���#7D���X�?r爻n�x:n3B�����? 7'zעU����;�/ǽ�I&�����D�2���������G����F�e��ym��δ�-�a�:�Yp�����WI�ۓ�[�^A��WVI{m'�ϣ�ptM���yN�����S��M֚Mggǝn[S���*��/C�#p��~�������&�]��CQ�c��'�0 IRYe���..������������u�����&)�xxx�(d�9�;M��O�:t��EPQ�� ���,m���J�AT�{g�I�FUVy��M������7�������D@�U�Ǚ3g�g���9�;KZp�i��9�4��\]��R�s����IHݼ	zШ��5��m��D����I��ry�7% �u/��T��Rǽ��ټ��\P�)�q�]_ϑ����Qe��Q�;����Em**��/E9~��NfBD��C��Ѓ�J��E�Ā$�Ŋ2�����^T��9}z#v�VR�7��J}��aa8t� �JLS����_�I�虯��z��Z��{q%��	H�<�YR.�Yѩs�X��R�����#}j�y��'m0 I`�ZpV�(EhX�.��M�.�Up��H'�gA��Ցβ2}�������/���ա$��#��I�qA�:�yd�@����]{�ĲE�PRR,�{�_ǔ.��rމ\�}��6�����X����H�ڱ]W����U�l�v8����T?�[�j��۷B�ZĶ��k�.���9�),"R��qH��ɩ���S�s
K���v� �_�����D5�.�{¿aC�ɩ|9a�̃I�S/�{8;ə[/����t�#wK	��Kq�t��B����M���7����QZ��F�yQ��0�$3�q�U�ƅ��c��m()��^L�V�^���q�����Sܺ�聭�7�mz���L��^^��Vw��9��'m0 I`Au(:����H�>Z�n���(����GM��BN:�м��"�"օ�:���ب�]]]���$嵏8�Rq��Q
�Yll�8�U;O��
������J*������,Hj�^����k���UĽ�y��j��^�
;z�q$)�{Cg�����x�X1�idKj�z!~.��ȩ"]$A���8t���1�)�m;ie�y���FxT31ھ_�B�?� !���� �H�:�2����~y�(r#�#�3�g�.j�La(�yZ�����7�..+G�}�< �a@�h��t�m"�{S3�=���\i�C�����,�1�e^�,���O��b�u蔂E��\�Hg��P�GDJym�f�d��l柕���u|���CO�����"�8��]8�Y���t��_�#��qu���'��X����������UzV��i�dHmMϑ�-��g:u銥��\BŰ��FHL��z����pt[��3p��@���z�2i�ƋM8e��5#V~ދ�$sͦ � ��6G22���r���ڟ��Q5�JU����ág�:�8������ܜ��Q��K�����NK���xF�y��R~ۗ��b@��\Cg�Q��TQ	7�sx�ˮ�{`�e��~U��N���u���� ��v���|���~z
E���d�ʋ���G�>R��󺔿fSHn���yҧک[���k�d�±��T��Z�d��kJ���G�a^[y�$0 I$�Ѯ#yH����߅DOQ��=�v�*TT�~*�ht���z�8��a�=���$�=z��*1�d��vb�H����}���d����0{�����QxF�Z��je�t1-9�L��OI��=��'�;��ш��we@��c@����\� �C@�w�~j�0[�Is��ڶS7����(3���	b�BoI��>�\���u/��L�]�Nҫ4�����z�&��^}�a���4%{A=�kw�^=��6UҌfk�i$��u$WID�ŀ$������;N�>����#_�V���Eڮ���ԋ9��m�#8$z�z�	P���O���q��15��u���s����������OJV�𺬦��q"�t��[	�춉��r]v��C�i��?�IX�v7vn�o��n�K�ŀ$��#H�gX,r�[���@�Xޱm�Z*�>Ğ	bϥ�b�g�U;�[����et�RZ�ū�Ɋ������~S}��"J9_T��:KwU���x�cm���nb��];�۴�Hhx����Ug���A�ET�
K�)㎦��
����t`~�Q��W@D����R�`s��1��<���5{ �ƃجNlb�-ww}?8DHeo���o=��$xxx�M|�z�k4#��2Oָ؈��CC�լ���HoĦ�iG����6n��<t�	���m
�""��s'د��T���$u��ޜ-�����ՓIT�\��G�$�m�I�9��8��,�~�\���N�#�p�ς���塰��������������F"B*]l�������^�$�0�C(..FQa!Ξ-B�z�Ea1����K�{z,H=����H�/�[@����u�1-Zb��4=r�^��z��6m�N&�Z�7K�jb�\��'1 ��u����sm΅���Յ��:��U+K�s��U`uZ&z��g�ؚ�����r��E~ܘ�[z��mh���v舄�8z8�'N�����1'F���ս�D�׻ջ���Bb��c��5׳�(����+"�0 ��̵���h~��������+�)�Ň��Y�Š߉Τ�CٺE��Xw)�m�C#��e��:���rX�U��
W7W�8�订�ՔWVb�>��0�kṛ�d�����Ā$��1���fjz���?��5fSQY�)���.m��<l<����وiu_-�uy)Kv�0��(F��=�� �Ub]lE�	�.D����Miy%f�g@"m1 I`�̚����UR���ܕ�c9E���v�0 �ך='��m�y2*�6��Am��f�Q3���k=.Et�M]u OK��/�2PXl����q0 �p��$F�DŪ�a���K?m��U�̈����ѣ+k��l�xY��)�K[��(�vo�Q$;�GӔPJ�5$).��㋥{1q|
����<�^��tI޻�;������uy߭>�����l�
�f2c�Au��.M|6_-ߋgol�����3\CL�c@��
u{7��R��O�NqY9>Z�T3;��q]�g�Еe��c�$�¢�e����ѕ-�v��E 9:d;���5���0 Iq�`�S�=Z7��;<��ْ��͕jN\�)-��[�{��x]��������h?�KW�4�ս��v||_/��p��VDg��rKdl�Kq������=x`@H{{��a6+�Ԛ�.��0��m�Hv!f��\���s,��(�l~ژ���<s�A��=�=��="[b@ҩ�k⚄��t���i*���ڛ��0$�!)������PV�����]��� 8;q��>_����ji�}��O�v�(��sv�Ȗ�d�����7c�=���r�Z�`�N.���W�߄/���RC_.݃��A��q��l����Q ��s,�n>��W�+�7�ݻ��������'9�l�I�^d�Ť��1@�'�����ONa)�K���B�z�|�^to��Ͳ����������u�[	����y��bAb&��1 IQ�ͪ��<f��Q?"lN���^���=S�WglA���Ϻ�+*ŗK����� ��=��@u':�"� Ou�~�@="�$)j7_���;۴!�"���^�����5���D8�-�����th�����2�`�ߤ��":��ޠ�[ ���f��j�	���-~�����_���ZK�g~���u$�=q]�}{WD7����� 5=�� �i� !�@�W^Y��flV�WR�����^�>�xq���(��T�5��5�D�$E�+.������G�wa!76�q]>9e>�K�y�j�E�y]jL4@_�~�kd��4�ر�"<3e=�u[�sXC�����7c��S �'��J`�uYq��k�52,�`{�J��޻�;����7+Y��� ^����F�5�����8�\����ՈN�ջ���[32�c=����ˣ��ǃe�/gֺC���C'Ϩ!鍱)�.�`��ü.mL4�ž3, R7���㭟��lG���<}^��#��>^�ƠN�0 IP�zU����1q\
�p��b`��ɛ�;�ץx�s�ܟ}�l�X�d{�ۅ�@t�	�\Na	^�����@�����5xeLGv*��()��O�0��I"$4��==�<����@^(��R�/�y$��.�d5��	�B�A|�� �-�2}3޹�bB������b��%�G������r�>c3����LHv*�X���0�:4w�R�@���6��K�K��k�܍m�-6�L\�����^���r<��z�s|g4�]�(���W�Y%L��/�j��a��e�h�<=u�:e�H6$4�R��<�4n����ig'��f{�i��Y�͕�AL�ya��Hi�{��uȪb{��)��F^����/��ͱ)h�؍��%����A�^I�l����R��V�eb��8S²�H& ��L]�;��๑��������z?>[�[��D�"~>�b��._��8��4����AEUH.1�������-ЮY�w"���F���������֌<68~�����x�/܍k�HO���Mc^L/��x��x�l�f�]P�I��a�N]�;Qy�^�|`@<�M����򝟷c�ޓ �()���S��7�C��&���}�A��$�khw��S��"9���Hv!�1s�p��t�I
�M��),�K�mRn��x��D���CIY�]u ��d�%)(.�?l���ø@��΋!3���+���)�3z�ۍխ�ү�CNG>o��\5������b��]����pm�����(�����uS**9�N�Ā$���Ѥ�?Z���0�WKx����]����]�|m2&q]N��J��;�ie�i$⺜�`7����o���� ������Ֆ�a��4uj�۲Ǳvon���to7c7�Du�9��Eij�������H�̈����G�MoL����񂒘F��=�7	��qC:�8�뒤�|0��o��0����ퟷs�#�S��U7�ӭ9n�	wWc���;O��{�iuDF��$���	�E�_*7&�`�HR��ޔ��� 5�����#qS������>��9d����v��#�'��68�������|0o'��>`��$�'-�vSW�g0"�a@r 6H�%��R��6�,(*�������c8p� d~��v�~��-�$���v��.�˰t�q��|���d~T�;1��oC 3��;m;2��AI�3����I����Z��,���zL�ŀ$����A:{�!��� �A�/!�~rʃ�WT`���X�~7~۞�R_����%��w�e�ec�z��R�k� "i�rye%�����mG���,��01�A��t���༣wK�/��X�����s�|D��oV�S�M�:q��������GPZ�+��喃��:"#c@rpG�1y�.|�0���H�j��сH�
��z�6joF��9��{�c���(��!�����始w�%�論�MV��D�h�m�����D>R�O����8��n�L�c���X�4�����-�u�Uiy��� �a��r��竇-lѤ�r�T�	���f���"���U�9��2����FdHX�V�e ��#���c��C꿉R�э}���x#��w�*�=��cY��Q��Hf���8���>�EtB��}q��P��.#�0�\�굩|�պ��9E8z��N�h�Y>U�=���H)�yC�*A�m8�o����yEe����Y�190��#��ǴU����G��kX��k��7kSO���{��8��;+�},���L�I
c쿱?3_=�H����g��	�.8�Ú{J�A�FeE**�v��#]Ε��sצӹ�Ս��_�uYũrtub4F�rqĄ�aP�H�K���~
܈��9�c�֣ ����\���d���qq�t�.�P�<��lbq��M�SD��I
c7�����h?̒8j�si쏇$9� >�I[�3�_��ù;ѶY z�A�V�����S��&��w����p���ET7����q��]�I+L�����Ƅ��U߰?K=����N-��&�-����]�G�(G���)��V�o��ȶ��0����Ƅ����s=�EZ�6@d�}=��|�T�^��MnQ)�J*PXR��J �wB���~�+��iD˄ĈDD�s8��z��1 �`������8Ŏ����$a@���@��g� IDDDD���D��'��}LHDDDD$�fl�k8*�}�����H$�!S�A$""""`@"�����$� G}�������H������L�IS!0�"""""GĀD��p�� �&m�>HDDDDdH2p������H��$�r��,V�!�HR�pIӷ�xDDDDDr0 �`�:�V�>""""r8H�-C����$�	��Śp�������I�	��S�L�������d0a>�4Ԙ��!""""C`@��Ȧ��֮e���Vo?���RYK��&��z� �� ")+����&�����ڜ���~��$R��M=������<��������a@"""""":��������$"""""�s��������a@"""""":��������$"""""�s��������a@"""""":����C�ǿ��\V
KAN�_���xx�T�*a����TVO����HY�r���TV7w�/ DD$����6��),.����5�-%Ű��=T�Ƅ�/L��NYG59����% ")9��S������ �Y0 Ia��X�<�	?""""2$���	]�j�i�����H$,&� ��|DDDD��HG�D~4a�$""""`@�@D	� -G�8EDDDD�0 �`�t�1~>DDDD$	�fL Z����!""""#`@��sȈ�����I
��p �����L�I
� Y9*FDDDD�ǀ$�ՄC$Z�#f-""""��I��#mY��H2�p��b�p�X3$���D��tDDDDD�0 �1!�H2��ODDDD�KH�C&\�EDDDD���$�\���$H20 \�����H$)���������da@��C$W">f$""""��I���� ]$���$�Y�F�������1 ��4J6`#""""I�d0�����#Hf������H��$0k�_�/���1 ��q������H$�:���F�bGDDDD�0 �v��╈�����I
�"""""=b@��b��3"q ������I�9S��ለ�������ŉ������H$L���>HDDDDdtHDDDDDD�0 ��&d#""""�c@����дyc�'�����da@���	@��e1m�$""""�c@�¤@��e����$�Y�I�9$	�Vs	s�+""""r$H2X�:��~>DDDD$iF��b������H$� 4�c'Nc֏������I� �B"""""cc@"�1gx$""""#`@��-W��DDDDDr0 �`���E��g�χ����t���c�*�p�������`@�C$�r�9?""""�?$Ҍ����1 Ձ���A�����Ȅ����$1	�!�6̻O�R�o��)$����U;�~@DDDTG�Q���� ٟ���(��\V��Jq��wEye�U�;�z��mX����<�7z'E���Z��r�_��c@"�� I��Z̷�Z� �������A���[�����z���_/�s���%�u��gK�Qt���Ҳ�����V����b���C�r���GQI���j�I+��jZ�sȮ��H�|�=���͚���(��7�y�aGK^��X��mv�Y�g*�)+���C�� u�T�����IC��t��c�"Z�kҏ��H<=�΅� 4Fs%�@�\�{@E���ѡe�?��J�+�#=�N"�`&R�gb��lTV�&DD����V��$��9��|WD�������+G���m�H����1ᮼ��-���yť�خ��LlQ��Jx��4C�1�O"�!��h
��]�A"���F~蒬�����������<�]ѩU�z�WRV�M�N`��,N=�-�O���̋�,WF2k���}�����ɂ�1MлM(�&F�}\4\��@W���nq���̘��/*��m�X���o<���"�y0 �J�v�5(�r�#}hD�մ�/��o���#>��-����g8�K+��gcI�!,ߞ�U;��k���ȸ�lH��tU;���h�kL��ى(�=�k,Ftk�N�����ZG��C:��h��#J`JWC�(�@DD�dC��ҡ�j�֊Y���5���P%W��q�pb*�B~��9g:c��]�f�v���-]�}�"D�����έ0�[+u�������A��cۡ�����J`�-,��'s7#�L1��,Ņ@e�&�zz��D�.���#!Zc@"�8ڒ+"Y���k�0�o"�y��/1�1�j�Wo냹��ai��t�'����ل�'rA��t:(+��\U�n���]����#8���v��׀1�㺶��-�����3�v�U�9g0m�|�p+��* ��M]�c�2�&}[D2�"1R$F����G� _��s��������M8���n""��l��zx٥M��� ?<0�#�^�/wW�y��i��w�o������f��H�r��u0op�Q���*KQ������v�Q�mO�Ai���(����MX�8�b�v��GTwb]�#J0���f���Gn�K�{�㹛��-8S��i""�2$�p�^_G}�Du���{���C:���QH�����~�_-܊�
mJ�ѥ1 i�z����b�&���|DTc)��xq\o��Y�.@��|�-UG?Μ-��Z\����׳��VX����K��}�|=����~鯗�7Q��eX#�M��&��O]���oWb�4TY9jODdH��f"�,5�F���G]v�ٹ�O�EȄ�7�+��VKv����<TBЁ�8����9r�D�ͮ����u��1,�͚4Ds�_�C��l���@�z������K�|[:�H[�Π�9��Ƞ��u��|k��VTJ[�T.���l���-�&m�3�]��*��ȮwM"\��`$Ǖt��)<���ףY�w:�*wO  z#F�ıb{Ɵ�"d���,D�'�P�S�^�BLɜ��(5 �2uRd���������$�+?�Ǝ�r��c@��s����9��e�K�lE"�%��	M���1n����X�[��W�u;�_X�Q�:���˶����'vd��>��H��_���^�QX�3V���߮T�Տ1���x����v�ū��Ah�/����k������T	Fi��Q�ܞ�/OY�����6Z�0�G	M��z5�G��~ހ�߭Bi99��V�6��|[�Gd`-B�{�C��p����L5-Q����ԐD�.8���w�� Jo���7)Z�?[1uS��ҹ��|5�Q�1 Ia�)vD����O�l��uFb���+v�����k�v������u��r��n��+^w��C�1���j���X���"Q�1 �`ڑ�����A�'�4�_�A���Qb��5{0]	Fkv��ǒ��_|3�~�p�z��aL�%,�Q���ō�[��v���7+���T�'"�!$���2m�#�������ҥ�d���԰�kv�l�ȩ�����ѡeS%(�ax��h��!�[SG�&�}-��MĄ���I�u""�c@�¤	I˷ee�"����=|�Z�[D���P$������o�������1�S�Q���)-e[���5��O����&]��l��L��F�+�H��]]��^��N��_��0u�v|�l���ǜ�������vm�ۮMBR���ӛw^�Acp�{sp"�������`��U�#"�jߢ)>|h��MEŴ��~\�O�m�[^Q���W��&KQ���3!�߹�O^�Y��@DDc@�c#Z�+�9?"28QB��q��~���ƿX�i�v��G�G��@<:"�z�I�>�ڹ��k�7S��B������1 I`�դ$�s~@dPb���������vH��^�ײ��b	���W�:u�	�I����ݿ�:��]o���3ADDH�%MG}��HĆ�>t=���������ά�X�� �|��>�g>[��߭ƽ׷���!��Ӯ߃�7i����>��7p "�ǀ$�i>f}_��4��Ft�ӣ�����s>�mM��J0Z�����:���W�S��θpGx�����섗o��I����_p��DD�����uCd2�ԉJt����y�xΖ���oW���xvLw��'����')��_����y "rDH2�5HX���O,���썈n`��=S\�I���ß7�HL�{����߯�0��k�j�׎j쯆�[��֥��a@����M�.���C"]��O�:~^�v}��+v��/�";�,�.�==�����c����hn����<�Ë�����;VL$"ÀD�nI��2�@�����x���v]o��H6�p6�;�+��a�z�"O��f�Bn.����A�n�I�W���Q0 Ia��ە�#�Q�����]����E��Ǵ��d�fՆ�ff�܅7�ꇑ=���5E ��c����*�>���.��$�9��Ί�C�lO����2oHii�ל�d^�jrK@T����f�ٍw�� o���ؾ�h��y�g�-��1 Ia�ƿ9s�����>=�[����v�g���'iEL�[��޼�F����뉪�s_��^�^-"ADdVH�-s�I3$�C`/�za4�"���zb��D�� �5�{�W�\���h�Ѥ��@,xc���g��Ȍ�H;A"�h�kcѬIC��֩�"��֏,�L6�h�A�<�	�q�5�;ަ��$���:#_����O���l�HCZ&$!��������GK�R׉�.(�=�Ѥޟ����}<�l�Z�����cp�3�j75&"sa@���m+kϑ��P$I��ʔ�xw�z����=�z S��6��F�����	*�l��4��LDv%��5Gbz�-�>��~`!�.#+=��9޺�:�~]��^�ݵ�dC_|:o��̀I��D�;ҡ����T ?/w��΂M�)u,�Lz���6�(ޙ�_��/S^a�Z,�����d��tI�PcaB��k��^m�p��g�1y�&�ь���b
S���N؂�ł���e�(""#c@����G�X4~���Ȏ"�`���x��5g�S��GDzv�D.�<���f�[\�M^���	�?>�^��U;Y�����I�IG��BQ]5n�^�~��{�c���sJFIY����Z�	6ywWu�a/�-,NDŀ$���#W�)vTG"��#1�d+s7�ø�?�Ȉ�p.v��k�����Ey����1n&KDFĀD��t�՞�N'��YS�l�����}��%$���O�����%�zb�s�p��_!3�DDFD��F���)vT;n.���(���7��¿f��,ߖ�k��3�ߛ�@_��ࣆ���o "2
$"2��>|=��������߯�"3�w�4�>�%~zyZ�j~������p���L��W����HCZ�YYȎj�Q�0�s+��[4�n�4��iC���FE�3Q�R��vr���|�Pe�VU��J9�(��BIY9*�x���������j��-�j~�	����p�?g����H���jJ�'��d��%��t��Վؠ7*�Q��Ղ�W�V�MK��~2Yy�8����|�g�aW�)���j&��C_��o��=�@���SZ�q��ʔ� "�;$)���*.A���R������g�*\���6]����5k�ظ��T����C!1dA���ѱ՟G>����H6��R��V�,�f�4Q|���᳿��.�����a)�<�,�""=c@��j�ֿ��;1C�U4��ĴgG�ӵ�&Ѣ�(�t���0�Mi�>ʑ��\Iz�'q�qDD��^�zK��GPVQ	�ݝo����_��}5?����W;�mM�^���fb\_S�cGW��섯�������u�x��-r�� oOw���J(R�Ȧ�/�71�%��tT�0�H?��JPZ����#LPKً��k�I�w���u�LQD�iƪD?s���޼yW?tn��y�~-C^�������	ɭ#�@Իc,:�7S�)���
��,D=���g�p���x@e:[ZG��G����;�hz^?/wu�%�FIo��K0i� ���S���-��$����q��.��q�rhM,R��Q7���$���A�1�O[u��*���>	�!�X~�h�z�>G4n�,���-�wH�m��=rƾ9K�NH���
,X0$_��X��Ɂ��a��#�1�H{�~��W�������:G�[n��;��߉�K����Ft��M����T,�z��f ����{}�:-QK׵o����de;"�$Ҏ��'�L[���յ�6��5���e�	8
7W�	cuF�v-��#�<1o`��!�~:o�Y�Mut��e��wX��x��iznQ�n���H�^0 Ia�ƈ�o���h�޻�ڣ��{���:*�DC���qxpp��՞�������7w��+w��9����)���oj�K�0���jYu-�R����U#�H7�d0��ߗY?"��	7tP7����`�4�����Z��~�s�n �?���/I=�n؏|���AI����$1����M���F��=�#�.0 Ia�$���;��#�:��8����������T��(8pϠv�s@;4�� ن��&��5cRd¬�RbM�(ܠ�^�QxxX��{ID$����q�XҘ����C����yŨѫSW���,�ѿ-�ӝ�Ȏ��9���KS����Ǻ��ju�)O����O�;cӾ� "��I�6���ҲL�k��QG��$��uGf�-.����Gq��,�:�P+�}�0���Q�V21Z&�Iz����St�|��`t�3�����c@""]%���K����2s1~�l�Q�F�J0���[�����5�F���;?�Ç?m@YE%�d��m���_��윑���M]Y����b@�¬�#ڍ�3��S��=��?0P����ב(�]l��iwWg<44�OQ�$���b���7vo��>�k��IO��ۄ#A���t��ջ���I���$�I+��m��==�;�Cjz�'>^�=G�a&��C��Ѭ���i�MD�9�݄׿]i�)d�N�+ߺC��v�c�����3SL7�FD���$�Vs��hZ�۔�Հ�=�Z��f7�.���rwU0���N���0���|����;�4�o�������WO�윉э�؈Θ8}5���I
�6hXŎ�IL�{��A�N���`.̢K�0|������}���x{����5��2����{ղ�w\���9U�،���\9���8|���hѢ�Ν�	&��Ym��4j���9���Z���cԨQؾ};�iH˄d�IWt瀶��e̲����/��ۯM��Ot<qS7��=���c�g`t�|�൪<):L޺�:�;9�O>��;wV�<~�x=z�>��&�~���1x�`�ϱ���׿�������1 �`ҝµm���3��U؞�]�s>>y�)��I��D�> s�W�u��t1���	#�P�O�+�u�fCz&D��>	�v){���o����������ޯ_?";���L-0 �`��_���Wn�omys7�S����~��t���o�K���큏��[4��_/CIY�JL�{��y�~FZyy|o��n
��@�H\]/�hpww���{���5�\��wrrRCҴi�@HR�5FX��g��G6�=.û�jv>�h|�~���)Xo��_H���]��q�?gz�ͬ�i���}��v�y����~�D��U�V�����D`b@�ƀ$�Y��,�c�0�>>o�{����|�������:="A�E�_:�6u!#O+e���׬������iز����-Z��
��Z/QrtH�V��:xtxg�4��|�,���,U|T0�<5�U���O������B�1"��w��7�kr>1��ϻ����SLQ��H���,�j]b��#�����q�9� �$�'��s��p����/�d&xߔ��㳿��o͎���	��/y���`Db���y[p׀����mL�k��H�7.�( 	bIT�st|
�`1k�v��j֏�.�����ݢ�G>��ҥ>VĢaL$��//��A�^x�e0�׿]���Vjg���?���Q$rH�z�BE�vE\,��3���V����m�mD7��n*���=X��0��ሮ��!����'?Yh�Σ��R���2|�� M���7n�d�
�Du��lۊ�}��1 Ib�'\Mi��L���{al/��jse���t���j���m���ߟ���*�w�v�6%ԤĆjr��Fu��Ui(8[
"�Vpp0���c�82$Ҍ�#HTC�#5-��ƴU��+��0Qm�ԣ|<\q��?���F"���{�.M����n�d!"�ivHD�t$+Ӗ������k��C.bg8��ر�=;c�1�P!i߱�x������N����a)�b�V��-�����Gj�������1 �.Y,�ɬDk����C̅�0Q}�L��{wA��%��Q=۠qC�z�KTz|dX'nKE��޽{�l�I16b�GZmh�������q�4;״e;�۞c0��q����3Q��ؽ�����`ť�x�����񡚜�k�����8�DD�c@"�p]�}��59Waq^�j)�$6<S��Yq
rlw\����W�,�Q��nVl�PG�ꋣHDd+|J�`5����U<9��f�zYi�.(�QD5����G���DZydX�Z�俿l�Q<��<l��^M��Q$"�$)�$�~\�d>b��[\�&��u�>��F���/�R�i�����ȩ��~/� #+_]���&E""[`@��b�ƿYsiB�Ma��#Fb�H� ق�łɏ܀�/M�ƽ�a����^����>ר^�x����'��ıQ;g�ępv���ͳ�5a�6י3g�������Ɂc��j?��Z��sj>�^�k�ja@�¸��W�)vt1M0�sKMε��I�ܞ#k��yz����Ȗ�H�7O߈��N���\������6hR򿡏n�6�P��L�G6�1-)��k[�޸m�9s�`������y����Xp��_yE�z����gU>iG�{�YC���:jU�m��k`/��nq ��F~��������(���I��lR�Pi�.�����ͨ��mC�H���n�޽III�;w.&O��$�%Q����1��59�����a�@T��� ����xi|/CLC�(?����\�s5m�!�[a��4�Eaa!^z�%��1 �>Y�hb푘���I�W�����Gn �"��M;���ֻ�~ިI@&�О��4��D��;�1���m59������]�;�`^�#��d��}��~�Q���e�ŧ�6���}��-��C˦�)TAD�ŀD�ѲH7�5�^��h�-���:�7u�dL��S[�<5���*����O4	H��<�����������T3whT�[l���T�]��&x\	HDz FTD`��󩩇��1m�M�*��
O|��\)_"��a@"]b<2>QQ�_�暜K왢w����_��S��B�E[a�>}���=k�&���C���ۥ�ADTWH�!6�w7�������J1z�Ԩn�n "=������_"��zu�x~Y�7�������ŀDD���D��r܇.p�F����E%eг��Ƹ{`{�Q��_��/x��Y�4	H]ۄ��9#+Df�����d�i�M�6���,��`�Z����'N`Ϟ=HMMEU+_iF˙E+��YBT0�C��l��9;Y���ԯDz%��}2o��?�J=������+1�^��"�~'d[ ��pww�ȑ#1j�(���OE������˗c֬Y�1cΞ=�3$ҎU�D�usmF�~\�9g��gMQG����w�C�����MY���I٣&}���~�4\\\0a�����?��>�rk��^	!������7�ҫ��\E�X���˧(HW���{� �t�����y#"B���w�3���s7���y���~~f����C�ǌ3��Ga�����������Ab(�{;<���s-�~jV;�^
ƴ�e�@h��àVk6j��puVtzm�?����F�X�p!:v�(���+W�g�}��cǊ#<<�$�Nܭ�Y����O�&�4�a�u�YϞ�Ύ`L+>z���@N^�('/+���=�)>������5i�7nD``�Ş�M�6طo�C��q@bj�}�5�pQ"����f�z4��Ӓ��^�4�-f�x���;�H	H�B��_���Y���X�n]���ڵkزe�7���b}ѽT�X����С��郪U���j�[�fڶm��W���q@bq����X��B��k����h ��#�:0V^^��m9��Tu.��s��o�!�rE�����6;�i�fͺg�9s�X��bŊ2M�������A����C�fwވ�����_����q@b�H�GEE���k�R��h<X���nMP3��i���3�=�]�c�m?��F(�	�mvL�jժ�1c����s�aYY�0*((�ʕ+�~�z��\�Dmv�N�<	[��I#�����iҀ�r�Gs7��Zq���My���}��I���zJJ@�6;�UT����l}��͘8q���H���L�4	6l�]���Y}s���J�S�l};�o[Wʹ�x�W��8:�c�!����t%.G/ŠU]eӹ͎im �o~���p��s�; ����q@b��Il���m�H�Ҥ�?*y*>ϮSW��5����"�7'���z�u�J�բ$�9���w}����ҟ�^�"%�,�$&�̶8NG�ӫem)�Y�C���z��H/m�7�l����,>}�����jY�,�ƴ$//ﮏ���J�{����l$k��"('$��Ny{큲j��W��M���WTe)%#����µ�������j+ӌ�Kl�݃�hD��y�>OϞ=��X\\l$+���Hl=���)���.B�Z��"2s�FC:6���WgGUW���Ni@�#��Ŝ��ۓ���{���g���c4���EJLL��*Tk��m���r@�юƁ��À�u�D��ZM�����ý�c�ҽHNφ�l:!�<څp@b��a�ddd�����5k��;G�Qt�`��hܸ���:�0��q@�h��|�S�lV�zʫGd��+P��U}ѩQ50�Gn.Nӽ	�[}jCm��qlhce��u�����<�iDRR�������w|�nݺ"$-^�Xl�z���2m۲eK<�䓘0a���������{���HL�S�x$M	m\]�9N]���u.}r@+^2�t�������ê�/h��H�ɧ����3�iŻﾋnݺ�S�Nw|���	>��8RRRDH����͛7�yj�

B�6m�9�Ç�7� �dE�k�+�
�M��_������{����ޭ1�3���lQ[�]���:}��	U|��&�9 1M���ŠA��r�Jt��垏���F߾}?����1x�`dg����8 1U�!���AF���]b5kG�ӻ��Qe@�.J�ڹ8)�d�ܸ�*�+Mrr2z��-�)���K����z~�x��/�ī�����8 1i�츄d�:7��6g�Jg`��G�Z��t!J΄,�hU��hߠ*�Cb�D��)S���ӦM�E�uKk׮�;＃�G��݉���4��C�U9ޛ�O4���l��ک>>Y���Df���!1�;y�$����@����ѣ�w� �>?!!;v���m�D����������k��t�5���C�����\D���%�;74$�큲S�E����i]LL���{qZ�D�����nj��A�94�����p(�GMhZKNue�J��r@b6�n�B�+#������Xdd����Y�y�"��LH�R�	�T�#�	mB����	vt�H����10k���*R���nZ�ڳ�1�o������T
��h����]*���#f���60��P���"�F5��T�,�yd��$�J\@҆��U��^7�]]0f��M�mv2�*�;�p�b4c�$��*Q�3��р?á�4T�D��܊�l����E&"9=�<]��n�p@b������տ�R;�u4ڛF|�̀�ua�m�̆�Hm5��m?qE� *A�]s6cj7v�ػ>�n�:ܼy̲8 Y	_{1��\Y�9NF�A�x�7�um����9y�P���RH0_aڰp�»>�~�z4f��r���ի��z�k�.dee�ݍ��pB*O�S=�1�ۓ��(�6��l������������$+>G���;�YK�~�0}�t���Ke��5j���o,K�"͜9S�/''�6H֢�2I���t��)"F}�6�n�8d��э��h����E���O� cZ��/���������y�>�����Ʋ��>F������U��	��
`rɚ��c�TO�]Xw�emR�1
H�Z�5��(�<�"��iٷ�~�.`��_�NNN��xӦM�{�n�o����[l���@��N���+݅U*B�-v�6�eL�Ժ�ZB*��y):U��Vc�,����l�2�k�����?���'�bŊw�U�V����.]����IO8 1�(�q�ѿz�z��\M��Ș�ǘ�vRt���Ę����cժUEzz��ǟ={���Ø1c���5k���w���&M�W_}[�����!jq�M�d\\D�H��PeL�cz��J��vo^S�9��WczЬY31�nȐ!(,,4����x|���駟�x�b1��x�|��w��WW帼q@brIZ��K���_��*\��#��Ԥ�?�&"V�{G5?HL{���+�rӘ���C��&O�l�233E%��J4����@���7n�-�d-z E��؁�������շ��3��f�Mk�0 I���$�Eyyy9r�J6��������|���&��B����:$H���^�NH� Ū��Ԩ�c�54�&ho�B��e�\�!3j@��1��+U����?�;f͞=׮]�LE��[��6c�HL*;Yc����Ůf�J`�����:A>�~j!�#��"�o�1��J�СC�u�V��ܞ(����E���}���t�{M��T�r@��n�*�ӯ�N�hOQ�H�v�\��;Ѡ5$r96��Ш�W��,j�{衇Ġ;�����ܰz�j�&G닌����$+)*���2� ������b��.��}�DHb�݉����������9�4k�ҥ�̙3�����6oތ�]��ҥK���v��w},1QΆ�Z��j��"� )���ˣ�nNP*15jS��Z1vO��xCm⒍��bL��VaƬm֬Yb��O��it[�l���ȒG�<����Ry�;HVb�c�Jeg�� ����򷍌�<�M5�j��=�q$vzV��sxy(���{)7K-a�k�ѥi����9��R����ǔ)S�q������ի�uJݻwGTT�]�G�&�~�o�6m�Z��xnH;�::���5{�[$�gyR;H֣ŗ`9*� �V�b����٪����3P7Y*�s@������~���S�Ʋ�i�x�QTT��'�����=��ԩ�ݻw�JѩS������/�/_�*U�����/�	yja������L�v�|O�q�I'筅�z�:ɨ �/ �Wc�n�*lE�q����+Ӌ��\6۶mC�֭���h#�cǎ����>G��K��:u�\���Lҋ�_�����
M�b�ݍ��8:�#��j�.���-vLcjժddd���OKK�}��'4�h����F�S(��$4oɒ%`��G���\��=W'��PcI��*�����i��yݦg˨ q@b�Bk�F���s���7n�gϞ���?j��j��4iX1�"`R��	��k��#0V2GC@�z^��b�lTNN���$''�w�����/���}��裏";;�$�Rz-�i���M��8�΋/�+����QA�1p���D�V�Xa�c)�<��X�`^y��o�Ӛ%>{�llذ�N��`-v� 4\��A�7Z���+H.Z�+{�$m����g*wk�"�--�m������Ճ��'RRRfR5�Vq@���i�lt���)I�$�X�d��e�q�Ņ�2�[�z��seff����`��w��i�DR���N�Br�cc���^])�o�0�,���K?z'�N�ڦ���-c�R[���
�Ab�����*q�H����1V2�iHJ�R|^w�+	$�R��a�ns��2U�c�%$�JeϯƘ�d%T��Y?D���Z������c�1�V|�b%vz�� ���/<\��&4B�1V�B��F�]������1����pBb�/��T���1�((T�{�������|0�ؽp@bRف;��MF@�p�Ę��嫫�"�=$'�c��8 Y�Nc��}�x��j�H�*k�c��Nm-v2����b�+$k)���R�G��XA�#c�+TY���u��b�+	$��iI^	�阧
� тm���{+���ln�c����ը뇍��}��+���Ԍl�y{�1v�\=�A�
c����+$L�r%\T���t33�c%P[�ENI]��1����+$��q᪕����*�p3#���Ѻ�,�$����e�1}�d5� v�*c����Bzv��s���v=	�C���SrZ�F�{Hz���2Ƙ>q@�}����A�;}��*\����ťd@mdT��S��ؿ9�zb�m`��ު��j���d5\")�,�
����j� E&X�M�1������2n��k�1VHV��:�����Y�k��q��{�KV_I�f��*�{1�ԁ�K�"$�Y�E-vt�8���A�+�� -+j����{��������)�c���J�	@�@�_��ةM�J͠����>�U���X�ETB��j��c�t62j\Y�9�8 1�J��Z�z��S�l]X(�3($�GU���1�hR����N]���U���<��1VHV���L�hѶ� Q7�jC��9 1v[BJ��Zњ�P|�����PO�/cL]8 Y�^g4��|�#�CT�N_�ǰ�`�;uE}�#�>+��u��Rp@������I�d�ǭ�|�l��ā1v�R]	��=c������!s��r��k�\QQ���ߣ#��pv��l�����5��6�&��"��72c�i�?�1��O�d������+!իZ��Q+����foT�t��i"����T���Y��Ȧ#9yH��Alr:.�$�r�M\�5�����,t�ie��I֞A���*�٬�Fj�� �5czp�Z"�F��EZo�c%�d5e�C���&��Ѵ��XH���{jSr����nO7gq�jN4����8�:��g"v5�y�`�$k� �������_��Ę18wM}#��J�r��0�XI8 Y��RK�EZǆU���p���y�� �q5q``�1
GG�^��㗰�D8������\0}�'
��o��	�v�2�d��k۽	�u{�F��nm)U}����+H���p@R	Z�@U�":��3cM�N��м�8^D�梧.^+L����p$��!-�JK���#$��fϙH0Ɗo����G�!tx4$�X�8 Y	��uѩQU�QM#oW蕣�=Z6�!�g��C!Ά_ai�1�q<7x�>M��VJ�[�h �%��S]n�c6n�i��,������Y�X�8 �3OwW����wB��Ep�E4=�qݪ�x|dw�ݸ�����M�q��U�
Qv<ML�dL��q7������lZTb*N_U�;	Ugn�c����8;�o�&֧������)�rE<5��8�F'b�!(-8|M��c�$c������M�����ZOǘ-�}Z}�H˺����cFp@����n;�#&팺��LS#�/N�g,�ڃ����5S�ᗱgP��ձl�9�	}�������٢]*|ϥm+ZI	H\Ab�����hP��a����E]բ��|�g�!=;W�sD��\��Fz�Q�M�d2Y��1�cq��9O`��Sb��>
G2���D}��kP�Ɗ1-�+(���6]�2�qo'Ƙ�p@��a� ��`_���延�6����$��ld�ӳE�u�dd�|>7C��ɕSqp����U�Ѡ���(�j��U��#=���m�ժC�����DĬ���R��6�s�#۲=�9 1���h����6�%���,H�1�8 IоY��P_��d��S(�p]�K�Ɇ��^MDZ�ܪJ�!|Б��kC���{�k��J��TI���`Ch�R�׀�К
J/���ŏk�� Ȭ�pX4��6Pt�Z��5�C�s��x�/��͎ٖe��C�d��x�c�(H
�h�/M�O��c)1Ii�s�Z�a(jۻ��Utl>!��.%����X�Z� �U�E�>>����PL�F��oW�d�� �hQ������tZ��U$fK��~��p�ME4��|-��1`�1c8 ��_��xi��jTS���'��ȿC��X�Mq�CNnv� �[:��'���N-C�=���&��I�����D�]B
o@[^�\M@vn>\����ti\Mu�p��5��F���NNgmp�c�p@*�u����B��R�K�E�>�%;��dD4���f��^qws���-0�_;�h�P���t�g�o��}Z`���v�!q��,�ZU��� �p��ղ6Ԉ�옭Y��Ԩ���BC�q@b����	��W���bX����oiFv.��hۉ��j�6�%�������[�F�m�Q��C��� �0���w�c�Z����d��7�0���4 ���޸�5�;��v����__Ș�Q��CaP�.M�W�N_�!�1ƌ�T
�ئu.��o%����gE0Xu�:��5\�2���4|�x�8�T���0���UQ6-Ч�~v��*���V�8y�2hP�� [m�,�v��	s7�@~A!Ԇ��  ����1f*H%����<7 �C��+&!E�Ek �f��Xa%?@����[��x|��*q�:�F���n�.LV���7G��%{0{�~r5I���r6�5�߶���К@�ߨ��+*����(�H�:��g��1�L��_�oҠ��M��Iٗ�.�g�ۈ�k��V���	 {��a��,|�p7^���0�\���㺠O�ژ��UV)��Fϟ���&5���[Sˍ�W�.�o=�'�czE��4$H�:7��Wm���Q`��?T���/B��7�3��0s���R��8.d��Q�����F|�t/�����Ѯ~0v~>o��� /M�g��ˊ�C���%���'4a�-C�vs�a՗1����Zu����?J��	�JeGvi7����kS�<7P�:����˘��zlګ�q��F���KN�������mź0�]V�Θ��}��M���z��)�ڃaxah{���._�8 ����>㩁m���P�h�qu��-u���I%[��g�
G�1�s婥���`�`b<ܻ����q�<f����k��|a�]�~�pf.�)$�F��^�e>�=3�����SW��9����B�?���X���[��kG{0�'_�yH���=�H��8���V8*��:H����=��!��9�����Ǯ#��7�*d�J��M�g-ۏ��c;��Ae���[���������w��W��j˱��@�yhR�8������?�_T�wdLMnf���MǡV�z4U|�ys$�'ر��+f��ڴ�~��X�o������������v�ILH&|���h���m����Y퀲=�_C9:5���f���X�`.ja�Fum��~�5�u���|o��V�ڴn4�r�硛7E�����p�J`s���_���X�`��g����+p��y��Q>��L�t��3W��_�X��xk|�2�z5�];>���؄%;π��5%��~���H���Q��4��5���15�ꑚ�3���H�y����S	�(7� K�J���G�{���֫���=�M���#ط�w�h1�Թ۰d��eg)�x7ˣ0nEp5��j��؟=��Bζs@�ȱ�N?��_���ʽ��c�0<�a�>�֣}��@�hQ��v�ܕ�����x��>CW���Y���=�ۺ.���6�QHR����~/t�f�0v�R*G9���l�YiOUd�"�*��:��{���D\��:ܬE�n:!�h�ddC�Z�$�In
�䦢V~:��g�j^|����p��5Gw\s��UG�s��igo��<`9����L<1�O�wͬ�����W�>t������?].�(���9�8 ��]�6 Ѹ�;�`lw9����W�h�u|(u�R� ��V�mu��~��HC:6���}���4Z�B�Cҙy�!�4�IG��8�&�݄��6�.:���S�pʹ8,�r���|��Am��+����a��~₻,z����o�ƃ�,��e�j��⨴���/~�j5}�^�V��HL�hr���Ge}�.	Va�o���t�h��z�����<��
�$Y�$ZT��H������Q�SW�֫0��	�%א���W��s��d;3��$�!���f���S���DoCH6��BU�u>�Q,�c̸��dqǶuH���x�9c`�zXs@�7W�R�ժ�R�~b��ѾG_�T�8}B����U|j�[���̲�p8be������0���e��oW��ZVɉ͡����d^G�|mmf�lH6}S�1#/{���V�R����'���Pk�֓8f���65�+��y4v�BҰi���?3n��K�ݵ�j���~<г�Y�p1fM��ۮ������fVIh���x�wX0�p��H���E�>�]����u��b5������Q'C(����2��W��և����.����_�ev�2%����({#��$�8��������[��NV��º����iy�tk�a�]�gP�z��D�K5J���ǋv�'��1������95%��n������p8bf�]@�]�i�QY'����/+ǻM�$jQ�v����Z"k�3$׶�i�xװ���:V�!{��\��.�i]�S����4��hS�?���.��Y�®��dk�=��m>	����8������1-x��6C�轶{�ϓWP�돘!r8bf�U@�!s^��Z�)���PZoT�c��
3�̍�`F�E�mu�WblA�8�ڹc�c0V9V6|�|��x��W���Ja��.X��<`�t��L�4;����D^�yV�;��ݢ��5ե���l>.&�2�f��ሙE7���?ֻ�����0��M(/Ջ�19�:F�'�	��7iT�����J~�0�?}�GA��_#}��a�[�Lޭ���	�^����5M���m9���v������6��zU+�b�z/�v���<���YRZ��j鵵�=ܻ���,�v��Z�98�n��O�5��6/����F�W��$���Yx1�:F$�_B�R��/�.��H�~��!(Y��k����\Q�����Ӓ7Gb���系�H�wp��Q|��m�g�Z5{{�6�iU������=w�IjF�tCD�̜<l:�,����*s8�#]���V�p��竰r�yXZ�����AI�-SL\��O�.���X̮��y�F����|�S2D%���h��)h#�?��ƈ��pH*�����to����A���QQ |o���cjCm����ڽ2�����hoZ�Ę%Q8*���=�#=�|@�}�ʲ	m�I����ʒ<�
�R~�ʏc���̂��i�<q�"&���W�kZJB��g!~�|��X�U|<E{^�)��dv'��{-!�����y�k��6B�~�r}[��71���s_����h^�jH9�#��̡�D�nޟ�����f���ͥ�$����ah|~�ȋ����lm��*z+����w}Z����Ş�*�o�OƋ�;��xZ�4��:m�ؔ��Fwp��+�C�둾-���{��5{�uhZ+ �˰�c�DߓT%W��Ft�r����|cL	���5����C�pS�&��.���*E����^)`�ΈB��8����=kZ�y>X����1��>&=�m� |��@L�l%؝ҔQ���PA}fP[��G��n�c3Va�G���Ę����7[��]�`tjdZ{�1߭>��mc��4�h!��7F���L�x3S��d8����"T4�������\|�B{��]t�����ɭ���[���rr��X��o��cx�U�����YO�+z���]Lz������P|�d�m�b���e�lQK���3�؇��l���K1�d��>�3��Q�xKS���#�=�IJ���<��1�����;e��c���w�zb�E�<���Y�ḯ0VC!����(�����$�9(0e.L3!33�������zg�`o�Z����<�[�9f.ۇ@Åy+�O�d�1��}�Y�۾[sXJ@ruvĤ�m�Ѣ�P;jl��e�v�1r�D�pV��ۼi�Q�������;ƭΌ1)4�h�����X��ՒS��+H�����Lՠ
����y�WG�SRss+>��BSZ��#��6�jҏ�{�?3
/���M{�6|-�u�vv7upì��É�8�o�X���,���Q|�����+��j������у	V>����x��-���9y�i�=��`D-��1&��-Ԟh8L����-���CQ��]����Q(��[a��o��opu->����;���o&�}�e���G"4+t�aW��2*���7tiZ��c��F�C������DV\|��� ��O��=���e��_���?��
���MkfL)
	s4jV� ISi�f���2ƴC3�Y� |�Xo���?���|
r���_w�(y{ſ�i`�7U���J��%$ qq_�P��?����6�WA~[����a�����1T1���A�����ZXX�����>��Ɩ������G4�JC��g�\��^�,m��+���q��$c�%���oW��3��M$oW�2e�Xd�w�m���I�s4�M�o��P-��#S�"C��׷x��Vџ=8
n��つ$Xj��75+�Zg�A)�δ�S���#�[��=�ZU��>�֞��=����
����tU|._/w<Ի9~4�$-Xw�ޟ�S�ߝ���G'a�t�LҤ��Fui$�\t3Ԓ�w0��n�\��`�C�'������Pk�Q���u��ŭȂ�b4d��D��ڨ��V%��$��W�,�z�Pz����P$9�kmJJ���wa��������_��g"q�b4Xq��sCۉJM�I챤��H��r� oC�k�dK�������_�b��ݥ��oD� ���]b9-k`H�CbX�i�w����h/��|�'��\f�T	*���.��R�P�jqP����e�cK���0g/i�JL�v�!�gG�j��9�e�h}���N������F�O����Z1�Ǎ�W�2�7c��0�?^.*HZѵi�����5q0�+��h�{�HT5���i�u&�d����ء�&ƣi��r�>D4؀���e��Q5��G�w��OL����,�OQ� �7a\�n8(qx�sCm��>���c�j����Z`I����Vd-x�+��|g�&@�

�Ч˰j�84�&��M��X+*�Z2������S�{N�����?�C�",�TEv��>wO�Il�g�c�k�$څ���܎3��JǢB|�p �үB:��ԩc#c((���FE11R�(y����m�CjH�6N�ۧ�	��h���S�X��<lMv���e-Ξ=�z�6Zq#5Kl=����"<3�uLh�}����}�S�Hkᐕ�=*GK��_BA�P�;{0FT��to��!A&=v��=8p����v)*�Oq{�?S��
�ƈ*'�|��TQ��;��ED������I!��*]�ݭ���>>sv�x�&�G�*Җ��Y3cI4m�B�)_7cZ��=�a�֓Њؤt1��BRO0f�1Gc���V�[�H;W�t���8�{Qe@����L\�I������$틊�e���Ԯ]\=b%sw7.~�j�JPHZ��{ᨫ��;�@m�t�k]�4�#��mlU�h�'��r>
��\���,P��"*I��#%(2�������?j�V�p�H�81Pe@�
I�������#�!�M�&;P;ݭ�T�q�5��;^q���"�.E�X����9g9-��E�
�Q�[ƞ����q�s6�d���.��@7�h����1p�����$��n�{���nYڅH;W�t��S	��΍�cl�&&=��Y��pY^M:�GR/I;��5hP\ae��T����rB�Oa.~�فA��t�I����.X�4�����8'|�d_ywlMޢ�/~�o��.iklDL2�U�jVc%)(,�m�T;�?�xJ�`���#�"�
H�v�&Ӧ�ѝ�-�.K{�i��J�i���RK����j�����<�㲫da�!$���7��<>9�O��n���unR�z4{��:�@�ĀV�_U�����=_������ߚ���G�z���d�%+'?[���,3���h(���ɒ�`:�ሩ���ý�#$���j�{���Ҟ�[Vf%�s2n����׼����������z"O�H��i�p�.�9���w���/jjSGK�;�S݆%o��r�浫���hl�:I�����㗗��V$�n�5{����c�E�]ǫ��V�u��x�#��p�TH5�����5m��{�w��24�I��q��TT��d���-a��)c�p����e .N����$bF�!<�|�R2�}x�gS�#l}����<�����[�_#�ex��n�s�i�剪�?�Clo kM�m4�c�G�p!*Z��3������jishfGL�T������f��h�������ݨP(aR��3а!�7�4��Q�"����G��O��pg/��nh� �'1�6��p�Ra���evͨ)Zl���_?;c��;���j��X��	�xzP0�u""�>X�ɰ�S[�,3���z�����" Q[���[����^'�9�b47v��+?��+Ш��.Oի�#��俙t�����=P�v���e{�axh運6��`w��������6��q2�iU��~�
���(���I~󗭆���|Z��v���]�3_�UE��U��X(M��v��Vxf}��ʩ" Q�)w�Zg#�<�ǉG�>GB��_�����W@@�Z�DW�f�H?��E��>��|�2UD���#�FK3,�������xغ��ƈ.Q�M�M�O��pJ�_[bA�ws�E@%�P�V�\�O�gT�fu.N����0�,o�ق�<�_L�r��i��R��~�B�j3�2O��Ĵp�'���xR��д@��_����̫0s���>CHʴW���KN����{��F��<�M��غ��L1.]��d�+��e��nA�_�F�W抐���-#;��߈���B����锄3ȜZˬ�����iw7�qo��UL�S�??�eL���F��q8R�P6$�8$)���(�&޿q���*�#}���иF��i8���{z ?�=��]�it2T���o������L��Q����:��#;��������ոZ7�S<Ի���QՈ3��#�!VHtah��*�q~��{�.�����B�}ݴ��28Z=_�[||�5�+W��*��=�a����i�m7i���cB��mH�anĺk�dؾ��>��մ�����]�ϓ�G�O������:�4�~�utS��țZG�Zy�3��#�1V��a�i�?�}���{2�"�e+\�@��2�#�	rr��E���p���G�����PKȹ�D4�^z�I�Fո����5{�~���,?�Kܡ�-ZG���gO�5:��[LR�|��7Ջy�������:s5�I��Ϭ��� ��:A>���x�("&YLS*(?o$�Tv1M����:�NTE��Ϳ.(�^y�״Ɋ��d����1t��R1\1�sC�5�G�@��­�˿hz*�-�j���?1w�I�|�>Ԫ���<o�	�3w��V/h�Q����Η�_�I_��2�p�4�j��D�0f��R����Q��JXZsě���;խk�������㩗��B-wQv�N��RȯX�����
4���њZ��r�Xi礯���{�YI����SW��O�����AZ["�z/x��u�w.
zҿm��/Ӭe�E�i�#�aV	HU|<1�K#����ɿmQX�1��a
���sa�G!��6�<Y\M2���y�a��;{E���؇��P�c�<iPL�a#D5�6���7�M+��"�"�&�J�d�|�d_tkVL�h��[�������R�I��6�e��i�UғZ����E���ʫGE��T��://�Z50�5b�Ν3{�]��$<��9^u�Qm?��㻊�۽�跧�	���6to^5䵐}�L?��w���rl
���څ�V���\�V�<��9[���6�^jtϷ���:�p�t����!�����=�'a�]���Sp���T|�mJ? Sڧ*8�2��嵤��ݣ��-<��l?>}�w��quvĐN�����`@fN����7Ύr~��r�,���yHJ˂ެ=�m'���a�����vgE'/�a�/�t�����F˺�R����=�Z�e��N�{@�Ӻ��y}�7Bvn����-��f�ժ�봫jUÕv&�d����\�x�,��i������xet'�z����qݛp@��(�.��>�U�9i��o������74��F���)�:�ʤ){&M��M��S�-���F�#:˝�H�����Y�#�#����hb�1�����*~�gn��f��U!�vQȭS��M�Q<�O߼���!��M���U��΃�J}M�jS/HV�.�:7�f��KS5�����i��WQ��x������ ���B�Y�9~��^�R�w���Ol#��tC����9U�Y9�#788;��rC8�?��hz�)o3��*{��w�:FG?`($)�W�-.l���V�����U5k��~p)*īɧ1ٯ��?��M'�$�H����.����:��(�=���Ҵ��t���ѳ˱�x|�*��c����5��^�4�~ݡK�T5��pw��}��M�)��T���_>z����f��G�4�ž\Ҩ���$cm?���^K:%.l�V��w'�&�af��Ci�һ!�8y�\)�X��<�t,������1�p����/s�D�)?l/�z^���=)WTZ�L�r��߁g���}�����y6�#[��AU\Zw$�]����s[��=���rH�Mh�G/�(z�y���l���Z�GTEJI
��i�������E�%;�H�.N�צ���Q�@_�6����<ث��0}��F0�KlR:ޞ����݋��aL��hf\zV.��:�����T���0����~ދQ7D��i��<0���rH��TB����۬|ߣ	i���,t��zu0rq)���̩v#ӯ�C�f�vt����$*I�Z�h\3���3w;���>9�1�b���}״"-+?.��_��4U~�
������9����($ٚ:A>�c�h�8ɽd����	���E���@�s���t�oҤ�ە��]�1!UA/8�w�l�3S1ZW��"���OS<�n�3xb@�RӧUm���-^��&����X���'����V�ٓ��Fj�ͬ%��Q�xc�Vq�P�z4�}����3ZȻ�H8~�x�Ι�U���V��w�J��g�\#*HLc81Pnɔ	J�OG��%&��û�̻Q@�*`:F��h}��N��JM�eg���"�����p�"�o�?_��o��o������v�N]���s�q�VtǨ.�1�s�;���D�N\{I8�������3�ɵ9�_sXTԙ�p8b6�\RHpe1���pT±�Ϧ(����+�V�*U*�4����Z���i�1ǫ��O<<W�RP3����7\�r@��u��0{��0���s�7/�#�ԕxزě��v�!qT�tEh���ڴ:z��%Z����*�����@LC�jĊ�Z�ߧ�2�>e���]�iLy�#GǿFys8b�Q.�WK������c��󊞧Cv"���dWW�re0@!�6�5��41����D�m9���K���.H]����0Ң��D뺁��D�AWg�~<F���IN����Ah��u���R�:U���������g"���Ul?qa׹��^��n�;cм���

�|�\��2)�pT��YY���Ҫ��5��d��M���*����&�)h���S.��E_��р���".��7���茕���W4��q�`���v[bj����q�UiV�
Z�S�:Ň5>О:a�#<:������Clg$����rմ�bp�l4d�����4�
����Y< ݺ�3f��0E��S������d�P���!�)�����ƕl}#M���CK78 ��FjF.�($�FԲ�:e(^�n�n>V��i���[hZc@%O��!ֱ~��]�{�x���Wj�*��F�!:�'�"�p�$��ZB��*�75OU_/�zoj����*F���������(�$
GΎƿ�w����yF�_S���k�l����ͪ"����|[#���̈́w��4�Z��l+���d����|w,\�忥�|�>qQO�������tД<c�-؎�G���~\TT�ׯŏ)����6�JW;����@��o�+�9���#f�,�Li�;}%^쇠��t3�N�Ho��&U$Ϣ|�Ɍ�Z��f?���W�ܐv�>�n���W��X�h�ؓ�W㗗���7;^�Y��Q5�Y
@���8���5���ݱk��t�,�~LCt��^�AVN>�~U��H����M=��҅�5���*;ɼ�}}�G?3���\�"~����HEi�9� а��xe��ق5.��9[�ѣ�,r��{7��.�1��=�~z�~1��(}bHLC
�S9zj�jD�$��׋�;��]��ע�.&�0^��}�̵C�q��9��6Û3���e�fE$��<�ۛ��pFv.^��v��K}\��@,���?�="FR�2:�"�Ծ�h������0fm�m�w�f��SK��1)�:ƈER��UMjw٩pS�J�3x�4-�0�"���ͮkV��6;���рdB��Fw�]�-�G�u�k>��-ARZӢ�^�Q]Y��4��OW�8o-�p���,�L����P%wb�
��1F$Z��W���^�1���ӑ�<�S���*,Mh��m�4����vx��v��f���1��x}����b+K�pD7�J�4��cw�l@
1��V�z.P���)Bk�(,�Ĕ�S{e�*zjڗ�6Ivq*��HUX�S��}��;s��mh�%��K�?~X��o;��6L�,=��\��!�m.�4��cw�X@��:�0И]�#=O�L37���*n�c�����g $7a�^f=-���篣K��>�i� Hf���F�BU�~�:
_�8�i�� cju�����e�s�,(���Ñ�p8b�,�h잛	o��O\Q�<��fn:G����֢��K��ͷɹav@"�fg, 5��Vv�EE"$Ups���{Z�ޭY<��r�Y*cj��c��x�V}ڠ��Q\r:�Fp8b�DH!�����~���o/�/h�Q�fŊ@|ٿ';g�aa��}�����iZ���($=1kr��1�{�=m��{ƣ��n㑲�Řl�>����b͜%Q(��"GZ�ሱRY, QK�1�1I����ܛ�F;����;T�`V@2�����h�{4��j�����MH���Z�{K�$Z���b���?oc�ҭYM��������Q9���J���cFY, ��dʅai�νY�R`�d�[�ۉ���T͌w4o�+q)FCk�h���f��c����\��=9�5:5�&Z�x�+o�i"m�hi�cS0�%�W��3�U[�.)��8$��^��ؿ�$3�!5�M�3�����V.�1!��9 )D!�՟6��[:$�M��3��_��ڃa`�Ҩ�������v<<c>����`���$\��Ė`���8�j��X@��o�n|x����9f,3+����º��*j75����9Y�+$y�:c�+�������F0f)SF��1���\{�\Ø���,n��Ge�h�]Fj`go��H@���"z�Q���ɯ��w���0v/��\ew8.��nj�Mf:
Ia����=�Kl*kI��kB^��M�z�ǵ3y�����l��,+��Ǥ/� '���LG���ER5?�r�ö����^�f~�f~P���,1�u�����EDL2�NjҶJԪ⍥o�ºCa"��8p�Իu�sCڕ��}��0��u�hUe��1�X- �����9B�̼c�����̓�^��p� YUtN]���c�-���h^�����{�XY����_��峞�#
HLC81f6$�k%����5s2�ױ�88�5���0��ȴ7�%u)ڔ
�A�ڋ��k���D�Y����X/2�G�6���)�}+���cD�����Y�x�uX����p8bL�� o��	W8�����r�c�$;��,\u6�A{�������`��$��J�w�Ġ����9�*Hmw��㵟6�HpvO�nΘ<�#��.N��tj?�a
^�r��1�,�N��a�J�lf��K�|3G�r@b���Hj�[8�
rp�h�E��-���3R2�_��JGS�&L_�����{�ٱ|~��׺�7��/V��e����MZ|eT(*{��Ϯ��"�،U���4��cRX& �0�.3Gٛn@~�y����Jef�.Ȅ��F�ҝdH����c8v)�_*�2Pe�F5?ܻ9�\ys6Cv.%[տm]L{�;��SP&Zo4㏽�h�nƠ5���j-v����O�5efo��l{f����h���&h�
+G/Š�˿��^�������T��{��ݚ#�q��f����$����}оAp�?7M�}z�jQ=b��1�,r��_�x@�P��\Q\`�:G�fV=�$�����6m^j,���-ħ����i+*Z��y��f�3��Ԩ��N�[Z��+�x��e�J�ή�LG�Ig��-gG�URA���uH�f~��qI�

��E����5������^��_����Ol�y�O���}��Pҋ���:$�*�Omt��y.��kߴ��ca���L$�"Ĥ��>1���L���;f;O]E�K?c��~�צn�??��'����'�0�˱<]L���%����T��$�d`җk�����$G�Y�E�������dn���L�h��Bit1���h�ɚof�6�q=���z���:C_��L������{q!J��۬|x{����x����*�J�Q(�p���l�,�G�Y�E�)�4(i����adf@r.R�?�)79 ���m����5�yy��
�ڟcXhq���;N���SՇ����XL�+�}��%��.؉�V�)uZ��1��PɄ�����,\Ab�0�J�e?����`f���S~�䑝�0kj[?H�=�k\Ģg��`����Sc�hx�V�����q-É�X0��p�X��А�ؙ{׋� '��c3M��[������b��s����ذ���8ؾ�8hd3������`�W��c�7����Q�je��5��r����#㵌�c��")7���br�2��	b��9��	�e�){999�A�_����YFDL2�� �j���a�fٖV��U���9,�q���µ�,�Cک�tk���ա6����7��\��q8b�\Y$ Q�qwq*�1nJ���'�NYu�����1?��Z����Ob�|�Dh��Ii��	ǁ���^�����iU[�+�6D���s�
0s�~|�b��=�0G��;��������3(��%"�(3�4��	Y\AR?Z��Ч�E@zB�����o,�O�'Z�v���޳�G��+E˺�mT����Cê�������x��u���q��
�$�+�S���(��fv���1S�B2��Pqsv2���HZAC����C���a���b�߷���$ڈ���ݧo���\�*ڸ��!u�@Ԡ*<ݬ3ҽ,�Ҳ������� �#Ƭ�2�\�/f7E��;���LQ`�#�k�\Mh�3�-�Y�6���Ğ��c}�Y����x~h{����c���5��=�Д����Ԯ~�CT%�
����2���q�Q��c�y�G�Y�e� ��bg��mnOb��3��Hi���)-v\AҤ�ix��=���B����UM��o+�;*1��'!<&	a���>2�&���������_C��+�~U_h��[��>X�S3����:U��$S����9��KYW#q@b��7�J��0 �r���Q5��˿`d�Fx}lgխO2����8�7�y��i�iDL
.E��^.Qx2�z���e�� ���}��?!�!
E4�O/hs��~�,�|LG81�
	H7M��T��M�s�ppAPA�.Ǽ�4{ekL|*�x�;}�}�Y��w�{6Ŕ����9Z���(B	�BkcҲrE��͌l�^Zf�S�J5���;�������_ oW������Wwx��ww�����_�k�d:��K�b��0��pĘjX$ ]K0^���R��=���������T�̀�,�����[C�F~�x�����ۈu?=�;M	�
n�`������bש�`:T�����81V
�$���L��	����5'ÅlB�?�.~9 ��d�W�LpPvq���Q��O�u�o��PUp����u�q�����Z�6(���`d�=Q�HYK8czg����a�1���U�"=`���0�s�m0��d��xG��W��h�1�iY(�I������������.EU�A5m`�m?qE����t��c�d��eR�](�df*�G�2#���vtG���/����_��x`�G����|R=[�¤Amį�6��Y�����/�G���e*Hɖ� �9��2�"��"3Ӭ}�"�=�)�LY���e����1�Oh�]��L_h@ů�N���p%.�p8bL�,�n��V��Xii`�D����݋X�@�	$���v]�J��6��_�bx熘л9��Ӷ�Q7�㺣X��`�%�S=ˌ����ɽ�K���S1I����θi焊Ee�ԓ6�5� r��.�����1��Δ�'L�h�Â���AU��z7ŘnMxB��Јs�p�i�>	fc81�	�v�Z��~�3$���D��VF�,3����0v���Ui�([LO�c.^S��BU��~�&�!`T�F�߶.�:�>���`���E���pĘfX, ��o4 5���
F�v13 ��p@bw�=�(<�Q��8d�^T�e�@��	����e��⠍U��'��unR�vv`�Ac�����?�h��0�&������#�4�r�h�s�kWQ�{�a�L�?1���{HM5���:{#G��{4��X;*M6���J�����[O����ѹ��X������G�E ZcF4��1G�i�E[�iQ'@�sv�w���6@�����Ӡ�?��^���O�Ӛr��ld���$>%߮>$
�ݛ�D�A#ë�*[3�n�	t��FQ6��ٝ͜81�Im�3�V�Jb�x�`�l{Gq��I�!�"(hLG(|�0o��n7e�G-j�|n�cJ�E;���{o�5ѫemtjT�G�����q8t!�N\ƺC���=q8bL�,���e����.}�qӚ�&���{�RR$vM��3o��a�돚q@b��rl2~Z�,��!����Cêh� ����4v�V$�f�0t�b�q�R�hye�T��4�$r�pQg, 5��, ����R�����NE��-�%`Za溴k��wT6bٔ�lN]�c�B-�t���80Q@
5�u��~��b������� ��aŁ("&��	�#�4Ϣ���.�q�Rӱ���wpR�}��^w7upt���!�؅����`�b�� " JH+�!q�u��������ۚ����ϼ���άw�3�w�������%A*��03?�B�2�_�u�#��`axݟ^��b�@}Ti��0jq1-7K�^�h\+T�R�!h -u#�P7*����l>��#�Rq�l�ă	�C��JX�잲�b��i.�꧰����n�rlE�Ͻ����vUnӣE����u�H��NNfAb������ֶ�Д0o�Cg�-��c��-(�f��5�� -�� ��a�b։���x�ۘ��d�#)#W�{�IΔ�l�M��,�K��FVX��$H�~�����I�g�x��(*H��CQI)<����M�"m;r����*R-$*�\Xxz�qbRR,{��[��l�*f�-V��2�P�oZ�8�{��"��A����@�����.p����ګ�vu��é�r��aP�^Y���_�o�bT��a
E��b�����]tki�O�H���0;"5�Q�c� �!}�t���Mm��f�s`{�ft(l��q8X���P�B��6E�ޚ���cXf���� �q�9�0K*�aֆ�uon����3H�06
��8$*���T)ɚ~H��av���3��`�����?�#����a��#�qX��]M
�U���.�:d�qV�D#?��:NT4H�b<��\P庂�^��o-U���	�0cc9JTQ�"X�FE�����s�i��Ҩ��ul`� �i=�OM��M0��4H�Y$��#b��q��
*�ܨf����cA�/�aF9�ʑe������^� ;�Z�_���:��J�T�����E�#J��Z$H�"9����޻<�q�ú�/�;52��(��/�?b��X��GW�C+sͣ@�B��}�"Hk��3IT��*�����mG->儜s�A�R�4������q.\�����׷���:50�͊'�D�0c�)G.��!Gc��"H�����Y�I飺5�J�('d�^N�g�Μ��8��ѡ���@�%���:|�����0���^�0c�.GQ<a�jDA"(�Θ j_��H�ʷ�8������,��Q`Qp�Ry�o�1���$��_]!I�0�gS���a�.��0S�T���1Lu�� ��y����h�ȮM��;->N��;f��aR��v@�W�����rͨ��Jb43���o�>-�n�v�i��0�T#,GL5�������Ǌ+��w�ɶoL�4	7�t��/"���j�������Ѳnd���yS���*��:OKJ~K'C�;�Łq0
��=�ٷ�\��z4���mt�ջN�a��FX��j�o���ѣſG�777|�嗲����7߼����;&N�����q�~���jAjX#���`B���It��l��x ��*�M����T��		��|���pk�fF�I�)�����a��&X�`�����<x�`��W�^��<v�X<��(��?���� ���޸��=ܪ��֞�0e�:���QPܙsʲY$��)�U+��� $'�����_\Bq�V�� ��Ÿd-�xE��1�0��r�������L!wrq�^�>>>�޽;V�ZFeAʗ}�m;�q=���N9S�oFn�e�"�"����Ĝ���T(ԮN0v߰�01ݵ�i�(� �-�Oߧ��m���k��a��X�'������{�O�>,HWPU���W�5*H�^�P[�X�ͪc��cs૳�DG킃I���1ZWj��n�K���^�iI(�L�����m�>���R�0è��D�Y���s$HL9����E~�U�#���ٲ(,��D�����Z��8qh�B�M���b�B����k\�۵}��%I������8�B��x��� �a�a9b��cǎ�ܹs�Y����Z�j���`i�d���Q��Q?ߺ�w���x��~����;�:��0&���X�
�:yh���A���O[������$]���$ 8�dI�<���m�8Ò��7Jf�a,��qRh�{���V��-Zg�Z��Ч���h��G��[-HE��7Z�2i
���c'PHݱc@Y�Żأ���.�g:I�h&	U��޻"�|a.��0�2,G�ѲeK�]�V��ժU��sfǂTM���] �Λ�NZ����^cE��ğ��X����������;�B#�,U��{]\6��X���2#�����&o���s�a��D��2ԭYm�F���4l;r�s�x��!�Sm�5/���nW#'�'Ft�Z���C�a����7�;rh��6�蓩FΞ���7�K8�hM��$��z�3^�cŎŅ�a�Q;�� _O���H�os��� �w��f�iРjԨ���[īM�N'f��M��V���1ݛb��CV/��$铔�-�	�mUH���	���\�P�X�9��y�X�^cH�&��d�����aF.�OX���V����k��[���V�a��f�fϞg�ZK����6�����,��� �ZA"��ŢO�%��;k�N�?���@3I�ܭk��LRR���{=� �_̄$�I�\>�80�>�5�:�=�ʎc����_7*�^Hǻ�T��U�H���������GK�Ʈ/�a��}��k[O��ݚ��(R5���H���E��9Z�@�B����vi��;��v4�Ը1K��@�O��z7���n��yfڌ������F��\�Sm��vx ��Fi����;<�*��t:��!+�g�3���Й�J�3�A�V����Q�x�<7�ALnjS���Ş�V�x�I�u���׽�!q��_���*W2�e�+�@}��k�mDu���%�FRy�b�����믿гgO0������"7�����Y�7&�²��Ġ�2]�q_xg���V����C��g����T#))�حd�6 �F[������8I�A�딼�^?&��D�vq�d�~H���9��ێ��aI�������]�JI�.xtx{L��j�㹱]*�����X��ؙy��b�46r��߇���0Le�]�L�E
���4��Vs�g�
n��ӭ��*,dI�NH��b���J_���P�:��x�V�f��[�Jдv^��/�Z֑e���zH�b������߯ރ���0vI��p�G��>�H�o}P��T�nd�ݿ5n��\�{���]�Sg�(�n���uI�ć�Mи(���YaI�F�nK�HRt�GC�h�	�������a��@�G	I�������^�p�Jw��":�o���h�'�X�-�΁qh�H����� �އ���盛�M\�[��H+�������ڈ�Q�b���&�&4�4{�^qr0�ǏD�ǿ��O�w@���_�cݎH� 5��jA�'��30�-۴�Kq��-ЫC��}�yg�}=1��UKޥ;���~�H�c�_�>�P8��b����(������]�Z�F�<� �a��&�xg��ܹ1B��N<���G�ŋk)и`|D7����e%��
7�LR����B���c��:��%�\�	�Y�i�ǘ��LI*N'�7{Dԅ/�����;���}.�B��6,G��1�����,����p��X>�3�`3���]�W܀Oht��u����iE%�+����;an�F�6�	YT���"#����:zȱr��
�݃�Lh' ��Z?���=�n<�Bjf,����w��W�U0�}}|��0Ѽ�������FlP�*�.�;���\>���]�v�S���)�޽�:، ���������@��߽�/�z�,�]���BZ፴���O�Ő�׮-�4��,��Ǐ�����W���|7 �ڴ$X#Iq�"���L�����"��r���{e\K~Q	68��."5+)�y(,�<��xx?/���^-c`<tt@�8L����b�a��#.��X�]w݅���
-[�Ċ+0u�T0�`S�D<��Z�z��	�C;6�͝a�֣��ӀF�\�g3�oH+�������9���b�������\�\<1"�Γ�(��6=��c|���&m�b�~,_����F�ۺW�Mjv>ޘ�ii�9����v�-�RUPI�����{�0c26"Gr]��lpn�?�}��	��='.�����vF��p�}��D�9x'�9��2&e�eb��z%�� 5j�Y��啗�1�6C뎛�{���`�$EB��h�$M{j���ݮ��/�X mv�h���^��/�w�6�O�=ӗZ�?l���b!A�H��En��������9$��0c6 Gr]��-ļ���������H�0�alN���ތQݚ-��%�>?���E%��n���E��s
�A�ii@����/#Ь�ŋ��d,�Fr42�'���p��I�H��1���6�đ�{3\���2��)�F�j�`D����9��	�.F^��H�aݾ���m�O��u����ĳc�`�W��8$�~��jǛ��-�.=��Y��*�@7|�[��l>�o���IA��S64�*��h [��a�ţ��T�/)BT֪ŹI��\��'e�5"r��B��yW��$I:I�`�$ՌƗ��m��O�M?\��S.I4� K�d_CwKJ�p��d��
R��1��X������y{��R���,0�ݠZ��j��2 �U�I��*�@a��Lb��ߋ�֗^.�Wy�@9��(�M
A���+r��A�7��K�5�$)[�G��ɶO1B�M3��qݺ\�Z� �5�tI�]�j�1<����("��N]�C�9�</�I�T����E�ݍhr2�+���������\�ݪ=�7�����BL�����ESn��U����K�ׁaF�A�������<�~�^��s?�s
nw)=u"*�N\L�0�a��D<��*�������r�#���F��^K�+o�$�&Q9p*�@�I�� 8$F$�RW*�E/FG��i73�"�$GI�tI�$�3y�IyG��Y+�q�a���堌�a�$Ս
Ց�����	3ơ3)�⏝xbDG��wi��X�d���H�����a⠶V]�\�oV�ƚ�'M:7����5��oW��0�aӂ��W��>X��o���3��H�'��p���'o�~Y2�����Ç�E�����lfP���g�*s������=��b�]>�($I�ە]}����q����r�ۑ$��R`�$uiZ�ຝ�/�\J6�`��q�����\(":��b�ϱ`����(4��놻Ftm,�f�Zw������*B��!7�XQ����6a�?��a�iA"v�{�/�*���A�HԬ�w~��=��[y|���:��$W	��'�(Q���`ǭ�Y\\.FT�T����0������^$I���$�\�Z7���_�Ǥ�f��7f��8U�_� �I�Ϻ!V�8���/�'#�4һ�]�h$�a�C%9��ջ0�W��Y~�B9�[�h��-��ه��c���A2Wen@�բf͚�������4|�~�HUs322p��%i�$�I�����xO�>�cѶ~��m�����㡏���=������0'qj�*t�"Q�������� �!���_D�����ѷ.�k�b�Le�]�%)Ϋ?|^��&�l��?"9ͼ��rI�I�R�vb��:	jR� �t�0c6*�Ս�o�����+Ev��/��.�,GL�j��ȑ#1p�@t��	�&VH����_�����cɒ%HHH ���2��@�v�޻�>�F�ӽ)R��������������7�]Q�fYΜΞBC��S��Y%��HIRSe�J��p�1�ѯ�����ƒ��#����Ղ���}K��+���:��|JH6z�F5C�+�ށ�$��lV@�0D�h�O0�TB��B�sTta��EH�(A˖-��o`Ȑ!b��\���a��2c��\����
v��	�z�B��3�Y�hì������C�E9⏖�-��Hw����>x7e'���X\tˈ��I�����TRB�(ʥ(C���Hr�Ą����
�	���o�ߊ�`�~�GO_��-��B��t����1T=����j�ڰF>~d�֏?Ӷ���m��ZcU��M����ť���yqQ�	6UH4X��2��8$�Q��D�:p�-ہ?���4�b�Ic���z�'O�H��A�x45`� |���x��PX�r_���L�Qo�I7w0i�W��!�gRM9�Э'��c�W�%w5�r�xP�7Z���+Ѭ=z{W�����K��L��W��!B��\M��1_/w,~u��2��H��ŝ/|�����h
%ёS�$y{�����,�4����>��a���w8v޲YQ:�eI��Z�)���9��zx��D-������㋻�Q�M`�Ѭv8:7��c�RU+��8��8o�ҥ�ٳ�"�'Qz���/f�R�7c_�D�9w�4X��N�`
3���|E�)�k�48�4y;�+�s�T�fg*fhH�||�[h���S~i��R.IP^^���nC5�6�{ş4��A-P���񮇛+JBѬ�iM KJ/�g���s�C�LEHR���������^��)�����Տ�N�* ���J�
��;e�&��H� y�����C�P�Ƶ�����&���删�ä����X��$�Y�[�ed9puuŲe�н��ʹ�G�m�6\�x���ǢZ��;"66V�6�˴b�
q��ý���$�Gz�����&\�<wn~}>68#������1��T�!<�un�j� q�(�p-�4K�$Q�oz�6-�3-���������f��ц*������x���RP���M�uD���B�8xZ���)����J��7â�cp]���uƠ����AEnA1��|j���T�����9��C��5�;r��|:*�,��k�ҍ�vqb�&�T����Ĭ+�X
�铣��||��"4���+�ޠA<��C���{+wh׮�M��I�&�ٱ;A"�J���aݻw"��ۤ��}nn��+6<+��)�h�Nps��[S�٤��(�]�8'h�]�Ӄ��+����2�BEf-٤���T�]p�p���bQd�F��#���^b��*��(T���XLHFצ����ٲ��D�[{53�^ΪaL5��]���9z�U�w`4�mx��q��x��>�rkw���h{�L�Uo�Vx ⢂q�|*.��q|�����OVz����3f�9b�~�?.���g�᧟~Rt->� �y�1#��إ Rs0��������t7���#&��6w����}\��D�=j��C��y>J�Lrbvycrh<x)v�pX��-����N�%+�2���� H/���"��D�Ij�:UPUO�3Up`����������,�єbBߖz�D	�q��C��j���3�?��'��bp�6ڱ���4�au�M-Ų��y~G�R3���>f<�#�67�Ϝu���7kDY�q4hP��-�֭��P:s�}Q^�֭[ѢE��ϻ��c�С���/��ح � ��<����~�fqg�N|J1=�)f�������sJ�%sik8�������>1�oR�<� _O,�$���M�Й���o(��6M���*{Q/��$!@�!~z��I;�U��O|C��Ɏ�W�>�:���4�����pW�V�v�E�M�}���ip��#�D c�؈]�3h	\'Dg��D��\:5�!�Č\��ffK�����C�|���{t� )#��o�PNЍPȝrTA^^^x������C��,Hv��mG1��PL����|�`D��[{_�.x&,_6��ps�Y�kcT�$�xᝠf��/�e��lP)��HӪ�I��m�ۿ��u��:�bU$�	�D/#}4�WW���:tF��L�C�*7:���k�]O�9Z으b���SF��QCPƎ�A9���S����ap�"��KӚf:2�ώ邧Fv�I4�D�K�Ծ���Y�����Jϭ[�N��P�����&�v/H��?��$̑$:AQ_�MR��n~�7�3>�D�9I��p��12�n�"�>h�B��Q�_�ƭ4�PA�t�����ǂ_��$I��ۖ��G0�sS��I�W��4p�}�LÆ�	`j�`H�(�s�1���8yI�>hԻ�FVYj��;o�,��l\���BH�o-k���1=��y�
*lss�Fb��/�)-�x�E�_;�1�z��'.z>�%%�-J���uq��2����D�$щ���Th����R^����ƭQ=Ф(�dĐ��P���}p��K���ѯ.��|4)<l���Uޙ���!����*q�L�r����ኌ=��+5󤦞J�Ȱ�+��9���l.�h,�|�o����0Ƅ�a���"G���ʧ{`p[<=���<ӗg��&����э�L�3_��s�¸��pπ�"��\��yFB:o�A|+�R����Ȇ�%3���~DTPa͚5��U�V��KI����#�0�DT�̙#IC:4��7oǘ��Rq�G �슸�l<�ucs��4����#�h�$F%���o�"l����-�/Gh�咔�M�2��݇��	�����qX������op���qL�|�N��
���WO�c�;`�_�j�I�2aF�>ϭ�EbD��۳���e�����J{Ŏ��Zr����+v��fW'J�40���C7�����ڊ�4����[9䥗^av�/�wtʔ)&��p(A"H�J���㺚�
���]��_q��:}4N��cRX{���Ob\��,̓3��;Z��zX�cz�!�x~l<3�t�&H����i��I��I�����\l�w�[�Oq\7�Ԧ�u�Q��ԏ	F�u0�s#�pl���"$��y���<k�;D�p�c{�ͻz�ʣTD��o#�vwCT�/�����J;�_�k?n c�8����g�By�w�k��}[�Pds��Z��P�ֲ�2i8�ߍc�4�|L�8YY�U�����̙3EźY�|9��$b�/[�Z!ޙ����Pr��w'�;�j&�^p������R��ܚ}
�r���9�t��?�����zHӚ�&a�>�5yx��&�A3F4sd�U�ՔK���_���Ǡ Q^-rA!N_<>C;60i{����p�#��-h^'��LڞB�h��۠���n�`w8�]姾5o�]��;5�}۠]�h0���:u
����yt-#G�D۶m��ob�ܹ(,,4k�T�{Ĉx��WѸq�J�-[�C���qHA"�2LI�e�k*n�x��~��*�|�\�^2T�z�g�X�m��I1�(	�˲�k�t��O���S�<���K�f���Sëll��c�S1���"��lH�B���_�����_��{,����L�#��R���]�1�����/���o6Y��f��z���d�'��k�^E�,��ۛ8���i����/FF��+�=������:u���o����ӱq�Fl۶M4v54������h��ǣG��_799�>�($��d���G���B�37ϸ��]�}��6yZW��
?�'ã(��rл4}�2Ѭ,��#��M���;
�%1��j^x�P��c�ۛ���G��֩����
I�9ܮ��?,݌Go�	Jc�1�]��C�?��'��4$e_��%�2��l���L�nd��$L�l%^�>�w�i�{����:#Ð�P�ؕ+W�-� B��ə�2dΞ=����>Ig�3E2~���u
���W~X�Oہj!8E�$m+�`��?�Bm���I��s�R���0�@��Mu��~�`�����{��V���ώ@˺�0���/V�SN����+�de��/��}�{�Cốy��碒��\2�@�B���%����nT�"ǡ����Z������Ȉ��ѵ��'�+>[�}Z������5X��qn�`Bǎ1o�<��v�¸q�p��	0�8� {O&b��s0�[6�4�z�Jw�}����eJ!I�.-���r�)w��"�
bʊ�B��&�|�.+D��s�#ɔ�L�y�Z\p��o�w��	�"� pT�W�%<0�^�~^��:Q[E-���?�$��$�X�Р��l�Y�G���,�zT��0��۔����kv�º��q{�"߂J�b��DSM.�m���>�k��-4�D3J��n� _O0̵$$$�k׮x�����/��ȕ�yO�:���~HΌm�l�tb&N�+$����������GK�ƴ�[T�3�	����@��@��7��+�.Ң�E:)�h���9ʤ��,�/{z�r@��U�s��
[ C�����G�:�f��f�h�h�B�*$�f�䒤f��mC:�Fz#�*�/�~?�ݏ�}[��#��z�H�g�����v�XZՋa�T�����&�r���`B2��K����p��&X�L"!)SD����&����A˺��ǀJ{��"�h����BϞ=i^�Iц�x�b��[��Y�����P��7�����2����p�t⢼�;ԝ�4&I�(�D�Ds��Bs���.*�.'�@�f�l�)zu|QZ���A�F�w�4rJ�"�:�SD��e�W��:Q�x~�������F���+1��mb�KM<���Q����ɸ��ƹ��{Z���,>+t�<,��^��5��t��7}��3��\��#�),.��u�BU�V�y;��1�QTT���hԨ�X��Cppp�<u:�fff�ҥK8v�>,�c�Ʃ�����L�Oޒ��n�f��k���Y(
%�#��P�rI�.6��Vn��AG_� �;�Wc{6��{"4���g��p��E8rV�>XI�&-I�{Z�f˞�\�s��ꡑѥ1ָ��Jw�W�����~O�0�9е�f�ia��#����Ҳ2�k+�wr�'s��G������
>�u�:+f�,�"C����y/�[�3���(��6=IqI���g/ٸ$Q�
���ļ��k�p��f������B"$�G��BSZ
�4X���"���H4�)����?��Z;��1���k�!�P'2P|~(��c2�UX�d�B�*���r��l`%qZA"�9v�'���-]�\(��;z`�M-1}�6��� �F䰐$Ѡ��y%�f��Y$�[JjV>&}�+wVo�!I$�E�K��}�yR:�
aN4c&G�d�5y򖎈
���)�!}���8c{4�g���3ܺ5�����Q�0f�#y�����٫����0��ԂDЬ�},ÊN�&�>�W<�����Gu�9�'��'I��VP}^��vx ����jn�~��}.�d�-�$�,����jF�\b:Vo9 $�^��/��e��!Ϡ��䩔zE�<�V����M[$*�1�ä�K̒h?9�#�~)'��Hv��c�(�gߖ�K���_�7�0���T��[�`ۑ��n�0Q��h�>��<�>�u��R
5%I�_�gU��D��g�t���ͬ�U |�ǿ�͊]6W2�\��%I2�GH�/~z�!�iR��sGN]Đ�f ;��>H� bt�}�o�>�7&�Ϗ����`ԍ���y�����]����x�۳r1����/EIL�WV���_�ƛ?mDD�����7�0Ut��sD)�G����q�L.K{#���<��LU.JT�X	��$y���=�$I�p��2M AbD����hj����J�#�,W����Á�h
��l�����Ѹn4��/�~����� F#}n.KR��XW!�M�(��+�0��>�\�z���v��8�Տ	ƈ΍�(m�E!��>F��sq(!�O\������d��f���q.���NJJ�*t*����pM�1�I���1���d���ό��߉y -ۼ2�Ơ��.X��+/Iڼ��$$��.���B1��*t��b���ढ
����$T-I=��ϛ��Ȩ 	���\�jzVHR�����=�lg �(K��7v~r�ȋ�\�	]eT���r/��	m�$2FT��X���+"$����+v��5��[E�ۃJs���o��)S�X����p���"?��Ն`A2 Ug�8�7�Z�<����W�� R:�>��XV�:��&Z�%I��d�7�Q��ݛ�[���M�y��${B(I���� _���D�Q]�/�:W
�4�k��:G�r{�0�����t�ܰ?A���ǵK�Z"����d;ǕU�I�Q�P�|x �Տ�u�t�{���xvtQ���e;D���_|ļy��~���7~��7������X�v-�z�-l޼��� aӁ3���xhH<��IT���~m뉅B�n=&��A��d5W$�¦P��$�f�p;j>j-�=�[c�������b��$L�b�x�W�$�R�)��8�P���l��%0Lu@ax�;5�=RbV����^{ݝ{:�>��((��0��r����F��!���������X�����`B2�Z���;�8q;v�0�u�?���#�����_��{L4�e�aA2j.����X��޻��K�c-t߷�X��悍�� �5M8��nPZ�49�$I��L��th Jj__��eo�t���0(Ic�(5����.��wn�s)Yx��`�I�h�=}p�����I�0�x�v<��
y�N����K�,A||<.^�h���ԩ�����u��ŠA�P\���P��mS���Wn�.Mkɲ_*�@%�i9y1��ŖC���Y$g�90�j�$�L���J���(�I2A��֏Fצ5ѵY-thOy���\���w㣥#+ϱ�I��@����G�U������cAR'�� nh�U����a"���0DGGI�ѣ

LK#��x@�:�Y��Op����aA����/bث?K�Z�Y�\�Dԋ�]�Z�����&��$K�4�0�ԷG�$�|�J�� I"�����[�E��]$)�ب|���rU!F���C����J�^�$�ޑcV�F���2!���02�r���vf���>��-
-�������1a~�5�Fᴉ}�~)ڄa*�$
����[M�~���"��$h���p���E3I�-ªU��� Y	��W�
Qz�����TP?&D,w_���\����yi��~��I7��.�HR�zѨ_;Ƣ~lH�5N<%㳉��R|�z�(���bt-咤�ڗ�a�kf�\��ˍk�Јr8�Q����{�.)3�V���mGq�iC�f�Mm�at�&hWua�hSa�#�R�,�8�ƍñc���k���=�-͛7��ŋQ���i#S�NeA�,�(�q�(���خhQW���T����k_�|NAQ�4I˿�8�	:5;�y�Ȼxy9y��1=��������ye�@��04����"�06R��6b������	�h�˒����r���ٵ�E=�Ԯ�ǘ��ʑ��<0@����ҍ�����] �n|�|�X���[w�F�X��wW|��0�~v6򋔍al�C�����k_?|��Wq��Q����&�����ׯ���'�YA�֭Ųg�83,H2B%�ii�0w��R�PRz&����<��Fʎ� O���<i�/Dv^<�ݮJ=�����NM(7뇵�1w�~d8y�<�$]7ʋKJ�}�IyF�n���r7��-��0�A�t^���j�4kFti,�<h.jT�c����9zhH;4�bp=��m�"l=|��c�>�<����O��hp;jJ���0m>�evFRSSŌі-[��}�����s�Ήu�r��)|���x��{�ĉ����]�����=��ξ-ѸV(l�!Z��б%h�h�֣�����.G)tG�?��*�)9�#�խCL�6�^Cq�S�_�9�H��;�?�? ���?��a���Y%���fkop=U�������ČQV����nĹ�l�d����]���oT4 �<,��_�<=[�1y��ǾƩKp$�Ҙ1c��ￋR�Pe��K��s��8~����[�`A%A��;{��[:�ۺ��}��?6�7&�������K�z�bVid�ƲWps4��M�k���y�	�����؁L~MBR&&���
	���Y�t� ��*q��
8�cz4Ex����/~���rt-��<*�WT�Շ���N��`����E���uχ��`�ʕB�M����HX��)��J�=�(��f�Ǡ�8Q��O�X�(��I��]'�|�	�R��,�d�>�{���	4m����?�}��(�F�˞�D�čl;b^��&Y���(���q{o�w�)B�$FI�Y�E̔
m��,H��_|���8L�<���ccc�b�
Q�;;;��~JJ*糹��|$����7%~vl\CT��׶.ְ�0<5�ӿ�'`��SX��.�s�s).�,�@n$���Y�:1�x��[�#��ɯ�-���|��\Ʊ���/����6���h�Y�i���'����ߺR�W��a9B��W�9�o�ۤ�{�p��g��b�Q#�_T����0��3�<�����t-�Z�!xT�;?��P̨���ବ,8;,H��e�Haiy��"^�_�8�m+������tZ��\���;�:��K�[����Kf���E�Gn틧�/7�^C=>��ی/����qL��JrsG�hT#T4Ϧ��K��U��Y�y��yl8�D�*�Q�S��	(�Ck�rݱsi����L���5*���褋�wމ����u}9�nݺ�F�C�EQ���7��0'��QaA�!(1�/i���F5C�	����o��� ����}$;��?Ҳ�B2J8s@N���s����E%��x���Ӻqm|���hgzձ�[�����B�m'	3�C�q�/�)����˓_��+�׋��������6N��UZ�F\GC����G
R�z<�� ���1b6n܈-�oh|�M7a�5j���F�Q�SO=U�yڗ�Âd��y*V@��5��s��ވ'Yj-�#Q+"��Pݤg��RJN�IƎC���>�Pi;MPt��`�J��yn6&��k��Tb��Ǳ�\6��_oL�&��a�n�$�e㥙�����Q���(1�ak�)(Ʒ+���fЩ9��N���22�rtk.����Ɏc�src��0��4[�nE�Z��[G3HT�n������o���Θ1C��]Kzz:֮]g�G6v�����X�%4��!~����i�?G�"��S$CS�$z�p3�O��WX������\\L���dZ2�>�<gzGoMF
��$+t���~��Io_�I�,����wm�w'�Ct�iX�Ɵ�l+^�t1�s�+�iʤ��^�.D�$W>�0�Ae�i�V	�,�$Ku"x0�*ʑN�2�#".�pj®&ǫ8yb���߿?6mڄ���g�)��Μ9�Fdd$��>t�޽�~>��C:w�I�G5@jV�X��J2i{���hĬ=R�HYi	tɗ�cY�r	%,I*A�D���랎�z�Sc0�gk�wu�l�����;QiI�F���P�$F~�W��K��oێ�'��]�3FPY�t�y���0 ��(1ü|;k�\O�J��q�<e�8AAAb�Gg �Jv��Y�Fl{-u���T�vڴi`X��:��%0�T��Y��$��/0
��S>�tE�+^y�f����{/.)�Gs����+ſ�+�>7$I�����y�87��+r����59�1�j�#��G�����ǹŨ4���*{�vZJl��"�<XT�3Į]�зo_�ɜ~Fiii?~�޲���Wb�]�$I*S�īMOFK��H�T�f>xx :��g����O���'��h.6:w��ȘH<���W�9%c.Ԝs|��pSKQʘQ �#��L��/*Q����7�~��8Jv�
��Q7��\��Ín�{�nt��Q�5k����4�4d��<yL9,H�uh\�%I�v�<�DA�$�D �G������N�4��ɉ�_���K0{�f��S�F�|��ՙ������v��O8y)c
ݚ��E��ׇ��)eF�`9����0s}3�>��7�lR�� ��32Br��,}^a�$%%a���&m{��)����^��?����y����/1u�T���:,HL%H�t�$!-QIJBY0K��tnR3��1�0��7���3�Ju���}C+��E���q�*�`�j?������>[GϦ���v�����x�֞�E������}�b7�*�\*�Qˑ�J�'��P蝒��g����ܜ[6*���z�M�>]<R��ŋ1g�����w�b���*�~�mQ��iӦ���Eff&:�-[��-�Ͱ 1�puSG�t�$˝N���oL��{���Ĕ�H�����j���ٵm�Ϸ�3|ag��-c1�őWƩ?�.�����v���i%^7�Kcx�[~��-��b��8q1L9R>2�й\���b�%ړ2r%A�,����%��������QSFlT����~Z��P�X*�@c,H�a*$��1t
K�$bT��%�rFti����#r8L��H��u#��r)��-OJ��<_��RR��וQ���u�TM��7'��(	�/&�g�k�z����{�d�QQY�1��rD3Gv,G5m���?�ٲn��KP�}D��f�����7%ذ1�S5��$��cI�Jd�~?�mS���NHƓo����W.��F����K�CФ��|�57֔���b,�xH�5�fLDm9�Ӱ�k���^-��]�:.J5AzjT'�� Gϥ��<kj,GL� 1�qS[���;��AI�n��v���i��K��/[Eo��YYP�p�F��Tƒ�
���y*���o�%�=�(I�^������Y�Y��/\wK�Ƙ�h���AL���h��[����#�,H�i\��KbЫ$���+9I<�����&�ps�z�B������g��[���h��eIr
����>-1�gS��[�:��D�w��`�i�`37�rd1����2���ڍk��S�f�ܙKd�/f=s���t��fRa9bL��1I��D	�De%�Ԓ$Q�q�b��[ŊEu*$IT,�JG��{����Q8Zá3)�������5�YEZv�KԥiM��ߧ���~@A��� �A�vqxdX|�7�Zc
����#�DX�� a)�h&��$]�u`Ir��4�J�+�$G����b9�A�ҭGE����X	ˑ,�[�� Q����3�Y}��ԇ�������k�k����X �c,H��I
��<JJ��%�)�$]p8t��ʙ9v>?�هy +Ϻ0O�
,G��h��:�'������y��x�UVg�3#Ч�y��o��)���e�a0&�rĘ	c��J��
7��V���utФ'�,INFq�e�����-�|8FFX�d�>���o����6��ĩK��%Ą��-GP���1���XN�$�]R�0"��j�h�$G�$�f���Ʊ9����k�b��6�tX���U�qg�����!���bA��<�84��"(jS^ꢚ줸��Ȯ�����?�)�dAb����j�%��I�B#Eo&�1Ц'K�͒䈔^.Ê'Dх��(ˑb���ᑏ�c�������������E�O^JGfn�؇��?eG�5W�Ou�Yi,Gv��?;�~�L�'#��JRKq��){ ��ct�O_�S<T0�L�dIr,Υd�ǵ����������r�8�O\¤�W��G�m�J�-�#��9���zU�{�ǿ�0�r� 1�P!I"'I�È� K�`��� ���*7y��Q#"���i��&�%ɾ!^���Ͳv�)�������������(*6V@b���k����k��|J6�wj��`_���*��/ƾӉ�?��a�`Ab�$)8B�&�"Ie!Qи�GXQ�|P��@��bp�ͻ�cܠ���߲�Y��x�Ol=S��m�"0*�r�:tCj�������h��������{��ȉ����0����KF^�=�%)M��hP/&�L�%IY$a!q1$I�g�@�.��s��Ԍ\|0���t�$ۥ���o�\�[=X���3�Yx��5`���%#?B��Ō���]�TF�\���($I��	R�c�[�}HgDG�Bb:���I�YJHR`���bl����оaL��w��^U��aFxT�(���j��I�Rݎ%IY���&J2D3IrAyObȒdS���,|y4|=�k�Le�)ԈQ�#�a��%�*I�F�$Ir�z��(L�	u����t��`&(��6�7m٨��k ��
��D|4gvN��P,I��?�. �ѯqO�ֈ�ƿ��͊�H���F��r�0��u���%
W�eLb�ڳ�p�z��� 1�"�uAa�T��/�tɩ.�[���G]�zD�ojS���Ş�
�\�A�z�7���H���>!�kGb@�������v�:��$�T�{��͊�?��5����檷�rUP�]�*۸ZuX����kV'\ܴ�	������1}Fs
���_���LJH��)"����o������V㹈�Q%ܳ$���c�V*	���"�,M����/��hғ����W�����n�Z�!IT7�����/&A��-���տ�c8,G6O�ֱף��/wˆT$GT�n��cX����}���$FԖ�2�B�q�}��p�G�r|��' IR�z1z�S��\P7t1DdIrX޿��Ur�p��44���m�Ѳ���[�}'�7�셯��Ɨ�DN�:b���Q�$]��Bs���(��|�-�Gt�f>d^gvk����������|�$�L��>8��ܾ>�+��,~��x��~ݽ�"���������0��ubF���C� 1�b���lH�+�dqC���Caw�iGD��^>�Ē�PP�s�#��~L0L�Z��+2��>5����㟭�%�� (�Y5FX������Ph�R�=4�.A焒�Ȑ$�t:�|��TZ�ee:Y�u6%K4ᬭ��Ӧa9�YZ�F��4ã&#�6#Ǿ�)Y�pZ$9�f(�6�
:wO0S-�˫�)-Ii��$�C��!Y����m�Ȱx��ǩ�L�el<d�>I���r5�8���=e9�Y�^rT�9���Xy�'d��騐#y��T	ɑ��3NSm�.I�LV�G�%I}�o�����tg������e,�b]�ĺ}�1��9֩!b����aQڡ��%�m!G�,G6�,�y���(��kw��p.%��b��Z\�Z��T#���D�b!��CL��m��2O�
wԖ��p8�Ʌ�$�Z!I�I��|%)��$�B"X�!I�����Q��{��m��7k���]���J^�\e��̑k��"�#��v
�*�V@��?X��W�C~Q�Y���q��u����֬V�۶o#
8�o�F8,GL5�T?޾"�^qI*-�"I4��a<j"��uZ�4�S����.�K�FY�F���HT�`9�i��ÃC�U��=��r�f[�D�.�-T�qƃ����z|x��y�� ��利fX��@EI�H�T&f�S�(F���~W�xs��E$��C%Ii"4:e�ڼ���v,I�b���;_J̆���y��U��-�x�l�J���_1�J�t$g��s�za��9pXX���j�� I��i�ҕ=Ni1�B�h&��N�E%�X��jǫ���V>0KUG��n�.�%Im�[�0,G6OÚ!�ۦ���ۏ�ǣ�.�M�*��������o�.r���0��a��p8X����)t���mԐ$Mz�trtLI�)\�%��С�$i�s�#Kc���6ZGyF��\�X��i���%X;m���ٻ��r<Ab9bl$�� I��mv���є,I� IRYh���PI�I���)X��3��op�GK�ƅ�E�Ñ�����o<7�����Z��J��>�,G������&>��9I*I��i�d�,��B��y��DM~�xdIbl�#��m�h��/�PP\�oV�V�}|��QZ?зr�Rʍ�ժ�ȃ�{X����]T�$��,I
��Zރ%U%I*�A�M��&����ޡ��\�mƗ�Ȯ�Ҵ��u�ߙ�[�����J�m?�	}[�]ߪ^���c�� 1��$I�x_�T)4%E,Ij�R!IIҀ�T�Ci
� j�Ē�(�Ե]�h0z`9�;�3���=��&$d��El��#ƆaAbl���xTE��%I
fIR���۩!I�:���0��rd�4�i���)���dߩ$��B�K�yX�����%I'IR����ۏ$�^��k�������h��P�S��
O�@N�('��e(����SX��`9�["�|�>O�'/*\a��2r���]���y�1����:� ���6/[��TH���$�09����������j�!���ຬ<���]Eu;U$�,��b�0J�rd��y{�}>��E%ʞ�n�r����0W;���(G�h�P��U�1aAb�����*HҤ�t���s
��
�����|v~���q-�32�&&2k�W$)-�R���3�Y�a9�k�Z���-,��P$w"��9^VT�#�1���$Q�����J�).�iI:���:�z�5�����)�:6�ap��0�$1c��$%I�d�	Ό��rd�е��j��X+,���<u���Bu��Xc��is@IҥK'u�q8����Mk�]׳e��n��ګ����O\2o�W%)I��(����%IFҲ��٪oק�^�o�#����PH����;%iQ��9*!�NB�X�;���[H�t�����P�tr/�AI:p:��Qݚ����E��RP����z�� cþ�wz�L�
��F�f,I�rY��s)ʆ��4,G��V.�@�wԠ�����
���t��k���r��),H�}R��䄒�n�i�I�/�vx ���
߮ܣȱ)���=��v����\�ғD_%��$1V�r�pйK� ���p�\�*�����7�~�i�%�m�#ƎaAb�%I��]�m��N����Cgѽym��_���X/��<,�󧌪2����{�;IR0IR�*��IKD��W-dl�#��tb&��E�]צ^�j�4(�>B���:�+,���ga��1v�H�$
7�)zMQ�4h�I���~����鎅S�`��?��%y��6���^i�8q�L
o9b����rI�v
W�����q.s�`�DX��='/ad��z�umV�6T�=��єۺ\�v�)+[��bX���qt����Ր$]f*��f��#xtx{���"��S���oֈm-���n��Gueg����롓��H���$�LK�~(��r0*=_�^N�M�r���8z���aʬu&�1���n�1!���p 6	�� � 1�Z����/�F6 IS�_��^��`��@_O|��P<6���u�v��)f��f�z�ѹ1��l�`?/���j�.l؟ Y��$5����$��+-KҍPXgt�_��S���4�9<�N\D��Y�0P����x{�&E�M7���I�!�B�ݧ`s�1�p�$��Y��$��UT���_����]�ܮyl���ƛw�ƅ�����������y��!*��k����������E���(�$+4�#�ɪ I4c%��%�:��s��������	��I�0�F���Š�W�_���)��߶�}��]�䈎�t�6ɔD�Y�ճE�hQ[�Ԫ�~����q0X��D�Q�A�p�+��nIzw�4����q&mO�w����yk!�J.C)(�$�%=I��)��cI��s�BlT�u��n<�i�7[�oJF�����TE��j��ȩ�n���D�볞�7��s��L���}��@��ky������f��̭�r�тaԀ�q\h&�LW^XAAlA����ӗ���7�,IrA3Xw��Yy�JQ!I4�Ē�>�9���"��nT�M��������I�Y��rd+���U;O��zz��,Ϣ�Ǣ��?��w�����l�L=A�r޺�7��;��H�.I��y�+��$ơ���ST�$����()-�����xpp;ŏGR���]�(���	QH!-�����IJ眤�s2Q,r��-ca��9-���/�Ԧ��^sD��>~d����E���6[�*�Ը&���H�R�2�▘�쵅1����+ Ă�8<jI�a_�j�$*ڰa_޾���˯R��W����ET����TR!I�?#?..6*�,GN͎~�l���6Հ��Vܠ2k���(?c_%�!G*U�+������ܰ 1NI�.=Y4{U�$4����� �,��}��:L�4�'�����%�@I��d�����ϖ��E��HXa�>�Ja���0B2���kv����ɩgzfzz:ujno�PU]�Vu���=��]5}����;�C=�
Gw�#�/����>n|��X������on��v����F�!i2����r;!��bѐ���F��pDQ�V���ׅ�.[w�?�En��A����}���V>{��28�鼖q8�ͣx��� $�N�,}�wH������ǵ�քWܰ=�����ͫ.z�т���]����W1����Z*��d�f���g�tdk��?�����ǡ�� �V8"153~�w�2|�7_W�{�t��;5X��?���������F����S�ß�F����f��&! �\�,$-����G�6�k6��+��B�����9_|��#�'NO�C��K#�K�ِt��R�w}<$��j,��u�/��RU��ý�����;>1M8�i��:~��~�g^~��	-ɞ������}yQϽo�dxŻ>�v���\`�:.�{������ՄpD�h>ś���bgz*��T*�Л�>�j���Xu���K���f�IH�)��R�!����\���8�8p���B�7��z�L��GO��b����S�G��2��рpD}	H4�����7���?Q���|w_ }��t�p�M�\����Ŏ���Z!i��(C<\;>�J��(��:�hZgCҁbHJ�<��q�&WI�����ǂ����RH�Z����	Gpn�MJ@���o����?��t������RH�?rg��CCR8r@�w)��܄#���DS��r�������KH����p�\�zH��IBR�ͽ�-uI��܄#��ws���!)::�nHʟ8v�0Y!)��4�����8��;�k���B8�s�@@�����I���|gO }�}C��釤��!)�I*��64��m���?}�?
�3��k��t���C"ː�-}��q6$�?�*-�ÝK��	I*�pTE�3��#����7st������䉐t����}�bH�/v�Cgw }������\R��1.�H��Hx��I����$x��������CR~���=IBR&bH��2��釤�Bu;!�1Gpn�<���?�rG�0#$-+����vH��ϝ�n�X�
Iu%��	GpN�O��=IY����n��+��bH�/v`�⛞RH�z�y  =#IDAT�_����E8�s��$��|>���;R�($ec��/�
7$���%77���8��Ȑp�&�	Hp1IH���r3ө�TI��\����w�-�IH:���NHʄp�&�E	HP�bH�/��K���������BRFbH��R�O���:�y!)3���pe��\�!i���9[�!��g"焤�Gpn��M@�J,��#Bn6�ӹcH�/��y!)1$ř����N1$兤tGpn�TD@�J�B����O=$�!)I���>;��UH�����@Gpn�(�����Z����Ly���E;�5[+����Rg�CȢCR����L�\�S��\�_�Y
�,B,�>1~v�W�/�#vt����&O����G�:L���d����r�,�qA�K��^��+ P�������ձ�H  Te��=�w�XN$  ��	�Sg,'  @B@  HH   		   !   $$  ���  ��   T�m�Bxp�he_4;ѐ��i*={�P-~�333r'*lU�����#,ks�!�M�g%����|��%��hxӓ!w�x�/�֟zYx�M;43=(��w<�x�@�_;�G���\H�|��7?�&���@F�&C~�`��ߩ����;,K�3!wd�?#�|KK�^r{'4�ɉ�?v(K�O��9���Y*��.G�!i>�`鹋ALH�P[{�+^�|���cGC��,��T�p�o	��2
G%-~&@@��-������5��$�m��T�%�"$����	˂p�a8�o�X�Kx��C�BHڟjG�)3IBR6�!� �rH:1zv&i��$��-�p4?�: �O1$-,�J5$͝IsC�Na��|&B�h�o�~H�/����ް$	Gpn�ԍ��Q.Y�UNHʇ�Б����Z|��C!7ZB|̅��E:��,>I��Y1�"[�f���|�v�UbK�O{F/���G4���=y6�Z���L�5L�;��|!L��	���6���p�$ A�-����m���6ZN���Й?SGӋ���@Ʋ̣YlவL���O��=G%Ŷ���a|�=����3=aj��f/+��	H� J!ipMȏݹ�0X��p��-�/ �Ғ�����&֣��4:����\�~�X8����A��au���9* ��t�L�H��pd�/�3�u�#�0	�w�p�0qoh�? �qfiu����t�?=�˘Q���$����TX��08s0 @�V�}-���5��\�y?O8��HP}3G¦�wCR
/ ����3a{Ǟpd�/�~f��|dl��a��  �6�::�a���0��M��2d$??���zf� HKg�T��cW1$���A�*$ A�R�KƿV̪P@�b�m�{�ÝC�x *! A�Z�&¥㷅���  Y�z���X�e�H�� �G@��f�N�Ѽp@}l<s_�ϵ��m�pq�$??���v�� ��M���\kk]�� %[��]s�����#��}So���	H���g
}�G 4��㷇{��f�87	j�sf,��|8,5---���;�X�"ttt�>����B�Pz�?�������G����x8u�T333Χ��+�����}���U>�/}����mkrr�ԶN�8N�> k�]�����½0��xo�������\���Gl��Q�Sa��]ᡮ�pn�P��L�b�R�������\�B�`����㿞��G�gΜ	�֪U�B�Sy!����Ǔ�^}���ь!<��cǜ#Fz�=n͚5axx�4Ht1���O����G�	(�F�7s$O�	G����$�����C��dhd�\���q���H~�������K�؉������@sY�`�p��@]�8j�V|���֡C�J3MP1��v?�{d-�{�J��x/������9�h]���xae�ɷ�$��3'��齡Q��������#��;�GP���[�gy�#�#�Q�:��C��͛K?v8���WZ�Ո�E�֭+k�Z��a!���{��	���fÆ3��G:��S	HP#�&��*vb����A�GP�o�^�ĠG���������ʕ+SFO��׮][
��)(Q��^c������u��]z饥��F<�>��'Cx��500u t6`I��yݶm[i�Q��1(�����_*���gqb'3�`�t��Ҩ��i׮]a����'ދb@IsƨܿG�'ƶ�q��^֝y0��- ��	HPk�j]���؋m��R=����c�=V=ei���.�����El�[�n����h�M��_�m�3�tO�A��k��k��=�gFé�` ��`����s�3#7���z��O��NJ�lGNm�_Z�LM"�Lw#����>�`��"�"q�&�jDO���'��|$<( ��$X�X*�Q��+��"�FՈ�k��&�s�=ιY"�l�RZ&��b����.+���"4�8���쮷xO�ꪫJ�Ĭ�J��sa:���	�  �"��M�Γhq�ӎ;J�å"��!����W:X�����Y�X�c����b{�G�'._��(���\\�CR<p6K�����-�`Qf�|u\:r�嗇�(��;w���X�x�R��u�����8�p�}�����@s���{b#�7*Wtq���{���`�XlH@��$X���RoqT?��/e�;3qs},Nc��(�מ����Žq&���Vf�	��x?�gu�Ŋ���f��zVn�J��s�;C$ �"��f7�w.�h)w�,n����ɬC���Z�9Z��hA���+�p������-�{b�^�r����L^/�E$�ZO��H���湜�NM��-�;,�eu�+�� nO���-�eu�0��'O�L���$(��J�H�.G���ˁ�u�˔���'ivv�t��B���T��\�{���w�yg���HP���$��x�^=,���X��!����K#�dg͚5��r�aÆR�0K9����K�Z]�����w�qG��F
��ab<��*ht˷�)k����F�G�;Z�by����JNd����T�\r�%��f���P{��f�'��1~���4����$�R�|��8��r���,b��$�a�鋳v�m�ƅ��7.S�˖T�[�V�^]z4���ƽH�w��������U�����5��͛7�f�iӦ�!�Y��l�l]lc�$V��k׮]��'�Ō3*�&~�1$�>�NI�ӧ�T!�q����\�fg4���C����^���u�hݺu� n?��+-6ˌ���9.��w�������e�  A52^�7�/��h�G��50�_{mmmM93�dqD>�������ח��5�X�<^�ݻw�����&4;	��^���� �f)�P��-!?�����\�+v"�������*�ŽH�V���b8X���ĥv?�p��ť�7n�.ř�Z�$��:N Ūbi/#����C�C��p���-v��/�;~�D;�=F���q8"�ɤ���łͺ���֮]�=��% ./���f�pO�ˏki��
  A#��ׁ��T����3��V�^W�u�b����u[���t8rh_ؿ��p�d�+!������Y�f)�]�x@n<{+�sfX�d{{{g�{b�&���@�HР��b;���m�٠�\�\\6�]=�a��u���������k��cǏ�ݏ>����kĥv����T����X��k����B�]ƶ�eK1��$�9�޾�hnn��1.ጣٓ�����r�XJ_Y����d�ܸ%��w�^;�:~li)<~�<�Vg��n���d��-^�C��C5$ A����7�R���(��PH�21>Vz�N�Ξ��[����?\z?v$<����t�Ng�31$)�P���5\��I���.~l}�����NZ�I<}�T�c4�r$�
��J��J�����b[:�����18� ���xb��EEcŊ��}�#	9��2��0>9y&LL���ށ0�j�t�ˏ�q��X��w���Tfӟ,^�xm̬C�HЀb�3v�*��B\z�o���Y�����o��܋�����7b�Z����u�K�c��}�ޚ<g\Rr���p�r�Ո����������Bggwy�_lS�v2��v1`����W��G��Meϛ�fcZL��3�g����_���=����4�Y��s�7l+��XؿoWj�{̬Cm	HЀ*)�3E##�J˗�3�O����y��i_Q��7]V�����0yfqK�b�>.+y������qv�q�=v.�_�m���h)�w�����P���C�kJ�X d�c���ղpG������"5�8`Ti��x_�m�����ĸ<���f;:���v���5��l�����}���fj<jfjK@�g�*)��EFF6פTs,�}l�`1$�+�j�R\�r����������指��ٳ�,R���Q%�b]�z]i4�Z�]�8v$LN�����tV/,���g�분��8c ��G��*�Q�*޿b�����Ʌ3�ǋm�t�\:j0h���6m�<�]�9<��=��w����b���t�b	H�`��r���Q�M�=Ǧ�~=v�p��s�NAy˨*Gc���ុ��^\�$�]S��NV�ZU���٢5k�C����~�9<|`w^Z[���|�޾�b�~qػ�������q�-.�SѮ��`H�b�,���ᚔ���у���/���f	r[[G�l��a������S'kWZ>�[�O@���+Y�tv�(�Jdc��BaU[��X����p�ݷ�Ç�V������Ė'��r;�q�hժ����q6i���Z��f3IQ|�����;��w��s!Lƽn�Ol�����ޚ��'�K�ⒽZά�`�5���;5�O'�CmH�@���ˮ\74����.-q���уax���^���
SSg���U}��N�Nl9*߫V�+U�J���LiT~`xm͟;��Y/
w����ňsm��*�'�����#�"g������v������Ғ���Z���`����	H�@��r�7�X�.m3����铡���������}�T ��J:�1Ţi�3<g&�k���������{~1$�N�8V���C8{zz�ɓ���D�ʽ'FqƳ��<]I�4��n������<x���/{	G@���+G\c���c����DpǕ7�;n�jUU�:;;���@8v���p3���9<\����8q�Hh��
i��vuյ�w���E��x������r�qi]GGgH[4�?�J�X�.�l�}�z����B�$hq��\�3���'�O�*0�%V��v�ե��Ո#���ř���Kg�ь�~�3'K��!V0�y�M��}s� �j�����^|�*���+�;�ʩb�N# E��\&'O���wW�'
HP=	@\bQnu��f��U��������k6�C��㣇+��8�ˣ;���b�*w_Fwwv�;�?�Z@�b����<���V9��=��Ŏz<����Z�Q����m1����Iu�h��W��3g��c���k��#��'B�$h ����Q�r�U��B��W�\�;ߺ�K]����u��VIi���ʹL�V,�����(��k�=w~�����W�=1�x��~�ejr"���Q]���۾Z|���y��1^�Ç�Y��$h �,%I{��u�Y��G�m)�6_)��έ���؁,��V��Қ�?[11�����0�~kط��s����+V���l
��X�3��5=��a��`��W\_*4Rm��<T@��HPgq�/���+��(�35�o�^U@���-�3g�q]�*�h�����g��q��{�Zjg(��2�/.!��f��Y��M����?V�����U���kh�TG@�:������r��,L:�j$9Tْ�cЉ}�J��ꔏ��,��[�]�����V��N�֕������۳i�e���}U?����@e$����2�t&�i�ڍ�(^K��'��QI�1W����eצW����~(����W\bg�]6*�'֧�f�f���u��]�����HTN@�:�dy]�\UZ�_��x�G\�3�ў�F��T�3ϛ�f)v6�t������5#���Gﯪ"]���f5K˅�u;�mmm�g^9R����$v�=��h&�֬�>r_���,�����]��5���F�vX�zCU{��=1^ӱ�� ��]���G�d`peU�b�����(�p�f�����ʵ�/���3�ynq��b�}F@��HPG�3Ϲ��W��0Κ�ڵ+4�xJ��-�`�JR��0�.������:;���ӧ*���}�� �O@�:�& ����zhi)T�!���T�;���j;�Rz⬧A��^�.<�뾊�.�$�k[�&hV�IWWWUk�u(i[/m�+�1���fH��]\�ઊۗ|z���vV=���رc(��uRm��|S����.�"5��1[@����t�]� ����T�.^[	�' A�Tہ�KϚE[[GU_���.Ͳ��V�5����Q��FK���-aE\Z�^��L�����Tۉ���E����V�,+O[[{��
������j��v�o�A�j�{T�y�*�@��jGKs�&
H-��f�7Z\��|ܼ^���;�3�g6W�F�7l� ��x}�cjj* ' A,f�#�D3H��o�q��.K��Vp�������[L�l�A�xhl������h .N@�:XLg`~~.pqq�Y5��^�jN�j��x編��D�}-�{�v����u���f���NP����ZŶK���T�4��˿��L�}1)$(��u��*}ͺO���FE��Z�y��R�,��<i1�	;흃�	HP:��k�Y:�;�:���jcq?����d-�[�����tb��@�j�ss͵gK�ʆ�f�ăOWXv�:m�' A����y'}���arr24�l,f�O�9��R���ci(\�^d�YN}o��Z�<\����㞘	�# A�t�ӌ��f'�!��N���1�7�?P蘿1���4cg@@�F��f͸������N
������ε㞘�a���ٌ��f���j`:��(H5��fǵ���CƼAe��FK����9�a3;�-��]	2�*;�5i�3vB�⹆�qO��H�1��������fǵ��H�1oP�i�k�Ӷ2�z�Դ(� e��e�rh|~N�F#  uc&h4�l������bdõ��H�1oP�i�k=�m��Ȏk���eK` M�|׆����P	2�*;�54>?�@�� c:�q�I�٣��s�K�<d�Tvfgg�����P	2�*;�4���Zf�=�# A��jd�ٮu\�;��L���T�6tڳ333��� cFK�3ۄa4v�;::隞�Ԇk��YtP	2�*;���߳��>3H�c�(;��<dLg ;͸�D�=gΜ	�ƌe_�q��<dL@�N3vtܳ1��Y3qV�޹lh�P	� vb-�JW��݌�It��1m�LM�v���H�{�O@�:����R699��%v�0SW[��
H��f�|���ӧ���@ =1�6����@���}�%^����@z�Y(��u`�?}��(q\^�D"q����ڊ�F�K@��	HPͺ�+Kͺ�$����@:t4k�5M�K�l���eP�k�i)]�N�
��i3H��n�|�Aɳ)9]�B�Ƨ�H|��6g?[ZZ��0��G@�:�x)����M�O��f:jH�6���Nb@R�.����3U'O��^�R:�@e$�oX�9~�xhf�mŃL[[[��q8p3'N��V�
�^��@�$�oX��.�����@m�=J������P	�$���{e:::�G�-1�Ңm�'��ko������;֮]�#�g��p]����T[�,TN@�:�o\RmY�xV�����ħ/.a\�zu�v�����b@����\.PFK�`�]m5{�,���=�FP9	�ha��Ҷ�ߵG�	q	��T;����t��X����3�x�Z��
���Ύ=* �H��<�ȑ#a۶mf(k f�A�Fl�7n,�P����b�~ӦM����jvv�ԩw ���ٸ���	H�# Au$������&Z�H���ٿ�L��$ -^Hd#�-�[�x�����Xf�xf��-^��[�Zf�qy���l��- -�{"TO@����D'�zF��-���U����Չ��rE���ׯT�=�' A���tb�799i�>|X�Z�C���QZz\�x�����	H� tb�w��A�/ ��Xġ�����H|}�v+ UG�����A����-[BKKK�|1�\���\��[�.P����xO�K��+���T����zr��tO �*���u��W��/n掣�\X�l
H���+�sO�\�Y��E��R�)	C���L�pqqOB,����v_.���+��W�^�v������؁�g�؋T��yU~�|����*�o߾@}�{�b���yp�x���Sh{���ʴ{�n�*�PN���#pa���
XcسgO������x�U]��#h�b�Ӌ���m��L���}������Mc���'^\�F���(l_;��%$h(FL/�Hiubсx �Y��G�)5�ċsO��)l�? ň酙=��Y��3{�x�/���Va�ځ�p~��p��W��H���p922:;;Ou��q�G*�;v�I���*\�n�� 4�X�)�k]�re�	�=Z�Gy$�ܹ3��8�&hL�beܣ900xB�&�yBmF�z����w���H ʣ�>���B>����R�)�����abb"иv��U���xV<`<v �U����+7}�힟
@C���Ĳ�6l���Ƶ�Ԇ ����i˔��ӧO�Χ��F8{VW�C}.�ٕ��vn�����$v��(�WӁ����~�x6R�{��Jm���l�'����f�k�1�B�fW�)x�����q���x��p�WsY�����#�����.�����I�����Ҳ�f/���kQk�ֶ ͮ���޿qe�#�>�% �qP9q�Di)źu�B3�g��������\sMS.����)}�,-��u\~ܬ�������ih)�hv�ϣ��ˮ�����W�����w$�H�/�l➃�z(��x�c�K/�44�8����=t������}�ifhm�=�^���U@���Z�_��R�s�=a���9$./���{K��HW,���m�vEh&��KS�?�����kn
�"��=1~�i�����������k���o����-=�s�d�����v�+�B3�#��.g'�ix��,gΜ	��G��9�񼣴g<�z$x�0�/��?��<gr��3d������,��l��c)�I�PA����e	��^q���޴���G�m�������  ��L�-���	�잱��-?���{�G��'��S��  �ŉB��syF@�ٗ]������������ ��DKO���,K`�;Q���蜥���c���{?����N��Ӗ����l5��9�[^����������?vY �k�u����w�e L省�ys�������>�8���Ua6���<U� X~���	@�x�~����}��/���O~���y/����� ��c����ƕ����k���>�w~���ŗ���������9l�$ �di	��� ��o�/���;�}���'~�=��8�3-=a�e(�� �����ٽ�'^�Ϻd�7������𕷼���w����pN�Vl	}�$ �����0����n�|��������_4 E�yӋ����{�w�S �!V�+��!	��c��K4��������?�O�oe��S���W��������$�9<�bG���� ��}���d~E�f��V8���|�+F�z�<�����;F���~�ů|�����',V���.�����֝y0 @#���@�� ���z�]�}����Hњ�����o|���c��l�t�}K�:��N hT���*@3����~�΍�?�( E�{v�?}�����~���mx�]]׆��������m�N�4���/��/�a�ߜ��+HQ\�����M���O~��������ˮ	F�?>����p�W> �����~���t�?�r�cY�zV��}�7^��/�ƅ>����=I��}o|�O}�ӟ����ze�&��?p�E>������g?��  �`ժU���á��7@�Y;س����?pɺ��.��U����p�S�zݫ��ɛ���O}��x�/��/�����/}) @=uuu�~���M�yW�����W�v���p9��������{��c������������ ����o�N�
��zk �zhkk����FFF4������_��U���$ E�w��/���7_����3����^�����}��}o��fg$��8s����?\~����ʾ��?��]���*�ښ�h�`�����7��|힟|�����;�. �=�yO���?>��� �B�Ї>6n������������y����:^���4 -x����W�t�g��_~�]��-�@��_��iӦ���� �t�W�w�����,^qö�����_޼����<O*)�lo=�?��w��+����_�������Y�&��?���n��;�z�  ����~��~.�����,����_x�^�.��ϗZ@Z�f�{�������^�����oyǟ��;����lG�&�:�ɟ�I���?����, @-�ر#�گ�ZذaC�f���o��;^���\�mͷk����1(���?�X��3_��u����o��޽/Ф���7���E��@���� T���#���o�~��,w[����^��y��(���4^#��������Ͼ��?���GNn�n�����}�=qz�?@��I��>��χO|�a��� ��ӽ�U�
ox����p���K�~�yWl��?z���~�%k����e��l�p���س?���{�ȕ߼o���xx����}d�}�����̽��//=n����O~2�u�] �epp0���Pi����,'�-����e��j���o�l�7]���Y�=���n����#�k�o'OO��������m����gf������Vh��{{�7�o}x�?}[x����{��/�η����G+A@X�fd�O�����������=B|��G�G��@>��k/�L���t�m������=+����!����D|h*��+�����a�޽�|������{�7�����/��?۶e�]HU�$hv�֭{0>^�������n���{�}?��7����{��db~~���{�ߡ�����~M.FK�c����'/ 5" k``����79������b@
�d�Ν_okkUe	;r�'�) Ԋ�  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��   аr!� �	H���r���$ZZZ� @�$Xb�i64�|K�t  Ȑ�KL�%7�Dk��x  Ȑ�KLK>�4����[�HS��.W�y�[Z�'�:	��B�p"4������(�����|�y���|��A�z�`�ii�5M@���?@��Ғ����$Z��eB$Xb�e�Phmok� E�|���[�Z
���$��[� uАz� E�|n<����|.4M@jk� АV��M���t};��
�S�I��h{4 �������ά���R4�����%/�k�=H���� u�pV�}��%�4���G_o�-��A�2# g��&@��-�S�}�7X"���6 ����2<������	����i���"�a�2!3�P�o^��R�z���D��-	��\.7���W�~WW�]R�ӵ�;C�����mX���@f$Xb
�֓Y�f1�����-��myw�n���3�y�|���e���*~�,�~�|>����p�g-;�l	H�Ĵ�2H---��ƕ;��TKK>��'�\�^9�W��G+���*�l����f����lB}�=ڶy�Ȕ�KLGG{��`��R}��#+�hp�����3H�Balff�/����f/�l�?f������ǲ~͖��L^g������dO@�%������_�cEWj����u�%���j�!����������^��ڞ��hd��G{{:�XVV��F֯�ޱ"��hkݽmˈ�5P,1�B��ʕ�_=|�ȋ�z����T�����믾����D�!lܸ�3Y���識NG�×n_�����ٹbw�������x�\>Z�:R�+.���C}H�]~��?�* �٣|
{����uWm�ҵ�e��u�ioo?899�:�׊�ή������;���%�,K;v\����vǇ�x�����z���Sˎ�~$X�6n\�?��=:z��t_)z��j��CC}u�[ߐ���J1���暝�������kuv�CR�@6mX���b ,[�\��O������OlI�ur�|��L�%Bgg��f;��$X�n���_����.�N_�oi��mb�տw��u�hX۷o�����?;yUZ�;�ݽ�!m۶��c��5�,k1�_w�����[�"����Hu������믺��f;��$X���o}����On�������w�ށ�=_�?|z�e���U��4�x�K_�����p����ʚ?>�V���Li˦����ǦM�����k��T`�QgwzG�C�	H��m߾�Ǐ�]u�}�����Rh�kk�|��}dۖu���ZȼD9Չ�_��������/���׬dW��=0�&�,�3�_��[;������k�z�cǯ޿��+k���m���c�����vn}M>��@�	H���põo-
�w�}�;j�|�|m_�[���U���}뺷�X��``�Y�r�旽�/������$���КTK$Z�Ǯ�b��{�w�����K^�����>��C�~�����𚐖���ζ-#�
@��`���+�����з���ߟ����9b ��
�ݽ����]3��7�[�8\����������n��ѣǞ]��C|)x���7s�(]�c�O����4��D�9Ϲ��]]]���w,f4�{�k����b��j��7�V�G@�eb۶-�q�����~���{���TJe^T�LL�-�wm�WYQ,�ύ����C�j��ӅB���������+^���)��7�y�=�>y�ԥ�~m,��;:��ϧ��F�oY��u#�)�v.@�UW���m�6��;��}?���T�������r�Z�/Z�f�^�m������H�����~��o��cϞ}?r���8zt�Ƹqynn����{���ݹk���_޺u�ikk=^��Γ�&�95>q����+���6�����+9�ϟ������;��=�uw��3��mٲ��q���5{����Ç�<wtt�3g�_�R(�jmm-�::�Zi�E�GV���-#�Y|�� O�ٹb�s�{���x�u�Xl�������w���Ǐ��ɟWhm+�����о�3�r�T�>}�]�pɶ����<46	��8��~~1��.�i#>\��@��q��ٷ��/<��௜���Q�׏K�FFV��MV������ Q(�X�.>�����N��݇~����?���ǳ�6�k_��hx 57�v���q���g�?p�9��ə��>_�%wjh��kW}|�p��PC1���������G���c�?q��y����o�Z5��c�mk+��! ������z�o�����zzb��c'^Z�x���Ԫ�ٕ��ӫ�����խ�±��¡���Cm��#���C+��w'�ׯHY��ٸ~���czfv�ر�����b��tpj2�zzU����b[mo�_l��mg����~ɲOX��M2_�lq    IEND�B`�PK
     $s�[�z��gW  gW  /   images/3024baee-4b71-48cf-83e2-7da05d24f50a.png�PNG

   IHDR   d     �� 	   gAMA  ���a   	pHYs  �  ��+  W	IDATx��}�]E�������M��B�� ��P�_A�O�C��ϊ,XPAz	B��Ki���M6������;���;sgnye����?/�޽sϜ9gN�937
Ny�}�^?�ٕ��#���tú4�Nel� �"�_�@	�B��)�D��*�ף`�w�X%B��e7�;�f�lH�{xa�b��Ϛ�O���N�m����ԊZv���t�JC�P~��� ��}��}5eUlO�e���Q��!4b�����So�31K�x]�}�	�@�o������i ������%������#-#$��nozuݑa[�P9��)���xh�脃*�[������
���sl�O��Қ�5nPN(j�xs�@��!�S�3�+�	�L��VW�,��ms:Jh�b[4֓zhsπ�𓺣���M�TSeY����28o+���v�[�L�7�QXVdp(��G���W#6�-g`��ȁI�_D@q�ߥl�0d�O�9o��(��(,{́�rO���16��+F>F"b�S/��,�z����N�3 (s^0�����4�L<`�iٳIv9��(^�P��msB�㬋���jNlHg2u�8��ax�Z��cgl�ߞG�.B\a�������I�2yK1$� �` Bʹ&����o����3r�ʓ��3B- j;��\�r�}HkGo�ա�T�Q�:��� �y��ŋx�J/�<(Jqa 툝��b���	���T:Q"L����1�.?��&��&�R�ȇ�c�|�5Fr�9�v�ԣ��T�*\��� �2��] =�^|L�=�c���%jV������qK�@7i��R�;�XR*(UF΋((d��;��V�޶ѐ�d����TS8Ø:�j�(:�K<tU�@P�ǰ�Q�i�3�B5��p��6�̓�i�Ȗ�T�́Č���xTR!��8n���eEYH�d#q�GD'��"q�0��؃��� *�� 2�x7Fw�W�m^����x�Z�Tc���{E��r�Q��.���Q���5HB~�wбj��b���i�ބ����$K'|���y���Q�Z�}���o ��xE]��ђj����#�@0�pJrb�ttk�i߂3��	����'��? �jm��'Am��r\iU3a��GAD���i!����U ��#u4g���tY��������cV���8Qˬ@�1��l]TI��.28�Z�n�6��sN+z�OE�G�G#�c�D�|�[֏w}zss4�3?8��P9ԇ��zAԔ���y��:��w��2�|^��$tR��Y��X�՝]Y$���o��@'T�@���4�)��RU�'*DD��mF�Ċu���k/,-�~����5���/�o�o��P*}J�k�d���X�5%@kKM�蝓٦���X�3�d�j�v�wG����\p/�}2��*�C�Æ3��l��(zSi�N�K��nj���t�w�a*�*�_W�pG) 	]�s��3���!�H&5u�"j�f!�	G]��d8�'8�Փ8ٮ�C�O�_L챯C��D�����Ġ��{��g��iA���u(<�)�9v�b�H�>T?�p�i��uꏻ�C����۞HS�R>�:[��r�g1��f�E
��A���^�8u��RUJ��z�����&~������Caޗ������@�h8���W��ď�#G�7R� ��)Q�RL��B�a*��ĞF�8�:W�z���9�8y����x�ħƔP��ax%�q���QS����y�.�����PL�S4��	{�%��D�kӵ�$l��� �.��C�B���-C�p=�m��$����4{}���J_7�q�i��'���2��cT#�r;������ QJ0��jD�R�bX]y�UX°�Q�6��3dG7D��y@\]��̬�Kc!v���I����/���,�f���ZH7T��O#�>���Ⱥ�`�2!�0&TCj&�3R|=��J:.�b0B�9<��S�$�|��4gN���1�r_H���h�l��NȄ��̐���$3άDH����'6�B���� �Ż �`�(�gQR"��A���M:��%����Y��tY�A��8Y��(��T���Q6K1W�B�AMͩ�6��
�;��y�z����=,����w�H�K`}*��:ԩC<�>����D
�F�~ee���ߑS�Py(f�����j�H5l���(/J��U��Z��)@I�Cr� �M~h�ʔ0צ�8�c���`H�7~�}z�Y�'�wPzp2=Zw�Ki��H�SZ��b�����~�,�g/�,	e��:љ�ҙ���4���IX��y�Mw�ޑ5%Va u���[h?����(�!��⹮��ğ[�h]��zטpR-��QDu�h�ruZ�F�pIYXK������\E�-PBF���mg�ϧ]�a�f��*B��z� ��4� �U�b�9���:�UI�vq�R��8M�F��9$�W���(5!�<E2���?<���1���\7R���bz�ސ�f֗:�"�HH(���&]�G����,2�@�	�:C�W�E�J�IZ��P���n��,�2����BW�A �,j��Y�
l[�c;����RG��`�n���*�H��/n9p�`z�h
���]=jK)�����`�P����qR��@���k���a0^�("KP�Z:��,R1�ZR�����&�ܦ��
�y���;��H�%q �`��0%3?����e9 ��vG
M ���Ԣҭ�U��Q�ː4�}02=*W����%;�)GT{��~��hP��g�lW0�Y���x\E��=���ns\fP���e ��3�f�\��CT���bxnԬ��:��4�%Y�w%b!�3D�mz�bN^�3���wט8��I�|b���J�����^���5�9�IoI{�����3\�fe�1���^�����R��6��Ut��X:4UlX�@-GI��{Q�J���{]�C�5�編DՆ��af�E܇��=Rg�N#%�N\#��j>H(�l� E��R�� e��z���D7�����8׎ȶ����$?,o�V��!h�"��g��Pn
_GR�a�yH�؅/��ψ-�����nAU1��p'�'�$8験un9��*�
=$W(]QQ������r��1�����!2�ҝ �L)*�ү;�����BZe�����a��PH2�@�S�IB./˯�&X�rG%��1<#�G�Ԅ����SL]�hPٲ`$�c�IG%9*G����DY Zw�Cט����$��&51q�q�c��Ɍ�!"�=@�v���l��iN��}z�!5� MM���;{!����,��Xi8��ֆ��
��/	�um �G�7]8��=�2�*y(9S�tc,��v�T��T��PSɹ|	Wz�J��qbu@t����ͪ��dt� ؚN�!|�,��:c�0zj��z&��E���D8LUO�!B\�ыn~��P�df	U㜻��?��s�cW���ވj�����^j��r�j4dc�T��}����'F�3$4�I44zh��l���A��Lf;#�c�峆TI��C=�,C�j	������15���?yO�PzZ��`QoC�M}_x	�E �6�m�̴���C�E���S�Y̔�ua)�;���[����wH'
�h�`����Ǵ���}����#��WI�uB&��v�`��	ً+�Y�gZZ7^/�P`Ɯ�{�P5�vr��"7��1ڂ���S�UV�%(�;���0X��~>Fz�g}����y��{3�.��-P)�![w�����t��y�&/_�O��>�VB}�V�T��"�I�ȯ8P�c ��\8������xoNN&J�DG�W���Э�1r�C3�#�!wt�Z�IsT��tz��B9h����Q,���MI�7_W��#�){�T_.ŀ3��䬲ǽq[т+�<��� 869%�^����	�������+�mk�2z�zTH\;��L�
h�iį�M� �1@���J��|�u��f���f���C����.�{|g�g�u�#��TwQ5ۙ^���8/ħ�ȁ#;&b,���ԉ�S�	�p��[�դWO�,p��c��i08��_�� ����a�����!:��"�l�ͱ4UY?�^�O�����2c+sa#�O��q�/	�V��SnH�@.q��&'b�d�,S^dT7@r�]���*���m�'N,f�P���Q��t�8�>��[�]WS�s��ޠ>E�?��]��p�͉�_ғR��z���ђ��ۑ�C��Q���4�.8*"(!����ǀM�;�m>u+��:���@y�u���Rm����^��iOڴ�.���T�����
���������8Z^�7���Ц�f?<�+>P�u�	�S�ܰC�a�G1:b,���ŗ��|h�05�z�����Ĕ�ȹ9q�!���3��Y��mߐ=�����3�Yff8�)u�f�4#C��:���m��Ld�	
����Z_�io�\�x��6��#��*fP)f��5���$�	���Ҭ�K���?�.�m��ϸ����3��u��1<�:��A�uek����(�T�� 5�0V�K��t�P�8�&�F+w�JBP)��hL2�d�U�Ĩ��>�m��J?3��1�9�	��8�Cģ[tz9�l��빹ϩ���mh�ȑ*��S�K�i�(.I�FH9�d�X���/�Z4JL�L�=x��8
:���f��"������_��qЅ7��Ҩ%֭�,WUJ��%�C	2W8'�b�?��d�K��r�o���3�[µZz�*��:�R��kg�c4�:�
�M���'��}�Z{ ���Z��9s~e��;VD� T qz/Jf����ޜm��|	wJ-d+x���h=��_dm�X��j�g�ɪ�!5k��m���%�]����lf%nR����܊F�ޓ`��	���ї���d1�YP�FɈ�����a"6��5G,��R��I�q'<�� ��!<�8�yuL�w�9�va�}t. ��KD���C�|������<=���!��T�g��3UGt\Nz7��	8+z�'9H��;.� 25/H8��S5�Yg��w��܀*Uy��/���2������%����1��5��е�Amo����5�?k���䩯C�=7��P�S-i�a��\�+\g�(wX�c�d�ޕW'x�e\�`Ɏ�%8������	U?s�S������;>�\',���2H#�qTbг�o��'ڿ�pC���� ^�g�^�G��{������8�vX�󨳐����Z0K�H:�r��2�&;4^ӑD;��6�P�x��J2r�A[к�YuQ����<6M��s	7��P�H����h����O/Rƨ���z�0�D���N��+t�uY�k&]�K�-���%{���\���F���+�D2j�z���i��Q�a:�Y�K�����ȫ5��Rz�%\=K=��ۚ���JW�B� ��W�����ǝx{�6G��e��b�O�S$��Z��㴱\��U�)�(~����qe��(��!rE�X�S.����Ϗ;�����&uc�Gtfx��t.�A g�S�6����bܧ�_���B�iY��<�G//^z�Ѝ1�)&CX㙆J�cxr�)lgā;xt��S6�G�}#�]�&�n+ �80���;H@�ܡ@�nfr���'^���:X�#�����R�5���y�Q��p�-ξ���~a���e�FR�t��zB�=����;ax�ƹ�:L]�ʻ�]�tn
�G�=�:p,��K���N�z�I�j�I?"�jٹU�������E�/Y����1�� ��`�YS��:·�!qfʒ�[bnJ�xi�q���#�m��_6$��ڋW��ݥ�R��L�݇�5+�5lk���>�=���Y�	R#��j�8
��>̭TBJ���}��\&����7�\��l�Q%0$K
Yn@<-��:#�8Y7x^r�,�O]�� �f��}��� mEM����6I���|���*h*��S��+���ޠ��������,J
�6t1����T>@��ԙAi�`��ם�w�ڵ��)�!���)@Nj�G�|j�a��0 ,G(�!�j� ד�OI`��$8p��FO?z�z��6P#ܘb����zq�ޕ:��qZ
���Rr�,�]��iV����8&�!�rP��2�1��Y,ED<��/�2P5A��`D�pe]����rOr�axǢ<�U�"T9����{�_B&]-�mj�����:PuwD[{ܥN[$G����8�>(8-< �0�Ġ8Ne�ӝ]�r@�I� �������"Z�����	D6�:S�Đ� `����vP�j�{+�=�qG�߭�U[�/L#&s�� ���֖�:gZHw�--#�4����p���f�h���{��Gf��k1�
yM��*!g.�!�I�*;���:r�)"�"p�[�����F�t�"U~�g�Pk����׽+����h��)Y"u����Q���T�f�S+��|i��g��+}�~'R�K���z�6!���g��~��xZ��?ǻ I��M�W��*��l0u=%��I���9*�^���?v�b���IASGGD]a)��_rr)K�/F��4�D�O�"D����k���w�H��$4Ofh!Xh�mCԈ��mӀ(	����׶�uT^�y� �%h� @K�!�p�"q��D��d�X$��C��������W�u6	�p!�Y�1;��Zp�R`U-��:�9\z0'�`�����%���7��G� �Hh�/��nՈ��S)&RU��d����Ï��/q2$ݩd��U�"�C��w�I~�XH_
&����_���hC̭\��pHq�)7�Q�P��b�0{�����{���>T^����1� S.)밥���x�(_.)�)z����xD��Kz��#�;�DY��,&.�eE@+���ZE����x��?�ƣ@���0������"�;寂�Ǉ�
���p�Kn�63̵Gd29\��5�J��7�@�x~h$>jM��d�57F@�J����G^�^6hmqAv�������례�W�GD�F�g|�ы�1p�j׈�r��Ԅ�G	L%���8�'�qɆf�=���l��Ug�<�!B����0�!@ia��/sq�$����u
 i<�\�W�$��'O�r5���U?`	����Z�T��AT� ���=�R�o��u�d+��!y����͔�地 7)ۨ
���{,p��3n��
��*j��Ou��R,����e�u!/+�;�}*��w�7�R5r�N(lV�F�º�� �(�H�j�ٖd����A\�����Fi��@��$$*޷0xڑ���Q���0Dl9�+!��DP�vb�LiDw�/_6�K
��s���\;���, �`%��}p���A�W���L4|D5����pb#}+�������R��B���u"~��E[]	�-� i1� �
�u��;�겠��H\&S%��! �)�k��s���e@��� �KK���Ii�>�F|�Kԉ�A�η3����qSI�R'8���3��ܓi>9L�{B��e����o[4���掐��\~��I�`3"�o�Q#aw�k��&5��vE����x`H�!��#<Z��l�g��i�V:)��`�#;��$���YSO֋����e&V�D��q3tR�����LLF���G=9%�$����KX9���?�~��*="߃�LY�} ����oz��Z�"�Hh����1���Yµy���v�,6f;��lU�,qHq���i�,�w?$�{ي�*!����;�������^Td�/=R�p�ԏ�3�}A��nU?L;႕]s$��5�?]����1���V�Ԗ3�%�yE���7�]S�kb{��8c��<�^�d�͗���6I�o������w�~�n6�y}nl�cjPdW��(��tm�>����q�����L����n�!aOgۦ\��/��wwII�Iz��	��y�����Ѩً2��������ͅ�0����F}��f��	��_�kR˱2�HK6H���V����W8�c����O�5bJ��|����x��3߿�a�@�q%P�9��z����f;�V�$�!:�>����s*@�9�eL�������Eޢ�@&�@���譹�A��:Ï�0a7��g�(O��1��m�3�l�y��v��V:�)���n�M.q���!�(����K&K��pt$Z^�O��P��b������&�b(�"Ψ��t�#���5���3-�)U��T����}z����9k��!p�!qM=3�Q��|=�A#����B�AgC�0 �����!�?���@6R5F�'[�p�nS�^6�n 5�+��52���ZxQ�y<@�%�����0����Ŋ���{�Խ.4�ĩuM�Q0$=N��p+�v븖+�b\����a��`:�ի*����5�A#\]&�5^�2ugӇ8U�T�t��U��� ���E�h[��|�eU�+	�j�xU�N������qL�ɰ��Z�$��0䃎e���pB�C4#K��H�4���z�~�^�t�a�9 (&:(wLy{�������$���(��fi6�r-7�8��;�����W�捣�$5xu��IY�CxE�`R�!�����f�s������Î��@�&��i�hw3�<C;��&�}�Ho�f'g�Q��ڗGO.�_�B�0$�k�%St5��Y���!���4/�qU2��O��Èh��)��+�ɐ�!����T��aF��:�?{�Od��2cK�5��7�@��TV�nk � 5#�U�-����T��(�R�ة��ф��C����km�� �NGg�����|+� *��g��N�i'�#D2�Q�T�Gځ#aR9�2o��;����%��4,�-�2��.��m��p"���h\����s!Fz�T͈x��L��㪵� 7U(�[����]1��3;����[㘾������M)����wh����i6r"�Y_��.�7ӹ�@�k9F�;� G���Җ9O$&`M�lC��PO�Ӥ�xy��)	P��@4"��k�rDr��c���oY�l���~q�Y�.���b��H�7R�p��$8�#��Y���D��]&����rZY�����5��	I(���Jd ���!��T+�@�{�2x���GV$�э)�Tn��8��fOVtF~>Vx).�f3�TWl�	�S��ߗwF��?��ӟ%����)�p�GN�/�n1�o�d��B� ��z �=��A"�j���uj��j8�2�� }g��~ֳ(gH4Na�������f�D'��H$�1fX��� ?�3���b���)^i�B���!��N�A��u�bx�K�q~���&�`FM����;��k����1>Xť6L'	w��/�T�	�GSi�+�����͌�k[�/	�n*iR\lHI�ʲ�S^�4��l-�*FNF����$e�e��r���f�%vQv��ng� ����� %���aCz�!����`�@l;M,��!�&�Q�S���8,wC�x�O$�w;�L�l ���H"yf$�Y�9����f��I�{R,�]I���،78k�(��2AH�4�~��HU�óϾ�]'�hvM=�Pf��su%p�QMPٵRld#�mV�4�Y�`ٶn�G�b��ZIUk���/UZ��-6w��9�� AY�����o���=�9zv#��쁁DR؈(1*+���.9��Z�?������vo\u)|�̣���v�K�c��de���J����&�=�����Nţ��������_�Ę6EA��,_<uo�[��D8V�L��=|20�~��
�v6� �\w�p��:X�g<m�p�	3��#��ky:���r39W)�!���'8:�z}� �:�f���à-�?���B��PU�o\|�[	]��>�a�"&_8�`h����k�x,
��y�\z87o<�d�'��L�-����P��{,�:��Le���S�S���]m��8C��G�h�/_p|����@�Z�fH�Y�#����L��d&�"�du/;q6<��vu��w6�ئZH���!��>v�lX��<���g��9c~�@�	���=b2����^��1��`dn]E1����E9�����>��9��*y3�<�q���,Ă��:t����k�CL$�E��'0�KU���GϝXS�z[���Ɉ[uY�y�$^7��5jY�#��F� ���S�`b]�����B�����ےC(�a�gq���m���1!^.�E1�gLs�w�@&(�-f�����bx8 &ԖBcU)���
�p� �q skY��=	�#J�<��6s���ϼ�T�H�*BCϐy�x��*��r;an �Ʀ^N°��cPH�Ie�Ӊ�A>S����8����XC|D،��g��t"�H@9gv�{b��z���f̜�W�P�kڌ�PS[�񌌐��%��J/jgנ3jD�f͙+�]�t���9�������<pNgp(�<���423s���&s}���b�F�hkg?w����m@��ю8L�6Z��a�����H���&s"��0�H��E'Bj|fí���tvBEe%�?AI����.�u��J���xau|��Y"��!9c����� T�Բ��X�V����ol����h�_\�
�L�����&O�
�uu�����P^Q!$�٭��;`Ӯ^q�����͌Y-�(S*�ޯ���N� �2���;ab�MK8�(���٢��`W5��-��-{`,s�~,c¸	��epC�6���*���oɛ!1F�7�/�g6��.<ݧ�����w?Hl$�=K�����@/��c#�׷��7���U�Q���+*���JpsqN�ϾǙ��"M{���[����	(a͞[|�H����W7�A�����K���Z��	I�3~gc������읇�%�X��<�.T��ู�x���-���q�S��K���C<������p˽o·/;���b"Ϙ�`��t82U�m������ʪ�y��Z�7q���h)�H|�yג��tMkvx���d��I�����8~��A������A�!}�CDG�W����T8��I��F$�)ؼ��}<�n3�_��	���-�p���e���n5z>د�����	w����ܞӿGb����ކ��	k�����M���5�6XrE�b����O��U�:��Eӹ$����j��O���e�'R����3�(p����7�*I����vؙ`�Ryy��d
��>�.����1���d:�k`�aq.�`�<Ĥ���7�������j�?�����>.��$k`����D	m�.���7���&9����˲�I6�u8q"�zs�;���Vy%� �� ��;���u�9טZ b����;�{V�Ћ�ָ� cֵv��{�� ��gQ+WA�#��*��*�Qyv0�n��}aA3\�%EPT�|��'����L	##$�c�\��tH��O��%q�WK,�f$),��Z[P߻���'�ep4x"��j�	Q����"��߿��Y����+��=�!���a��W��/(�$�07��R{5�,l���A\R-)��-��$k+�ڌ�������k�;�{��%�YJ8CG{�N��C�ioeg�a_��&a��N�NLK���@�>@
-�^oX]�@��������j��a3JYI<VQ�/��E1w�Q�D�u���?�Qfk/�i���22��ݟ�;be�_NLGb:���2�o�����}��b+��Uz+�3	���+<�J�!)��|��!��h!��e��u�N��I���8�j~+���WF�i���|�a�|��)0sz���5�%P�B"����ؼs�k������DTT=�ۼ��K#��=��a��7'W���p�/�s�jj� {��i>�z��I�������'ô�Y�C��������Wê�mjy$N)��)��M����WA �i�? dP,���2؞�`<��W�SB�;�(�0t�3�s:
�=`���}g'���[;��;�������G��X�'��������?_~~����|�N(���#��e�qӯ���Yc+��d�3R���m��էM��:j��N�V�`R1��
��ѓ��c��k��|y-<���b�j�Jڐ�i4PR`���28j�D��p�3�����͙�c�I0�AiA*�j\0�
n>k��)�c��7X��XF���2Ȉu�!S�Ϟ�+��_>�����a����@| ��������~x�5���k`����I�%L��|ɱ��I�'�lk���#YP�S�	����8���9��!����N���6Íw<ooh���gRQ��B]�&�,��X|�"��X�u7\������ރ�t8��I��-��e��X�m��3%���F���Af��p�����5��>���姡op�3BL󴇒PVR
c�U�sF���@{�����P��$�#�C������9��f��{��a8���ֶ�3���3$�;�U��]�g$�|дF�5SSH�?<��x�����(�	�=.9�d8a�<hWe̘�ܰ��!�غ�{W���6���C��}/������Y��Λ΅n�;_2��diLYZ�r�ײ{�&ǩ��HE���N��w�R�Z��S�0`$�0�=\7��u���x�����<��DB#?ul5|�����.�b�j}U)�,�3�{W�y�-�郯��V�dN[� \�?��'�}9���ˎ�;�"�#G��m۶��w�T�Pl����tڜ�\ƟS�a$�^zYH��.8
��;��|���#�����#g�/�?������b��ŋ��S�ڟ<�Y��҆L���0	|�[�§�9�������;��B�3����b<�s`ڴi��3��5�\w�u���[��������b����.b{�_��ޏ�<[��9pח���?|�xx����u/�������[��'���?� ��w������r�E�]}�@#��dΜ9���k׮����y��a>�a���T�D��N:���rx��U�8����-����b��{f���Ͽr��#U�3��?����6��+�$%�~����76@7��1��?�<<��000��黌�����/C�r��H��B�*J�xІ�T_8z��(����X��Id8�9_�d��p�cʆ�N���ULJ��O8 �_�� �H\dps&"�"%�����n���Z.���o��Ȃ�
��iF8�V/����������f�N\��@��H���� �Z���s�#�+����3�fk�+K�ҵU��e9�JAO�w�y�L&����x�p�i����ޫp�CGņVЍ=z^�����ж���=�4�ߏ�vȈ���w�)��LJ�!�yw�.�u�^ܜ�1�
�%n�L\��#����^��z+�����ŋ��/�!#lBpd-�>�e�v5!��:`�&=ca4��̀��m)7�<ǘ��e[9Cp2r�JT[������^�ux��`���ӓ���s{ӥ��Ų��S������#>U.�9��
�logn�ȌD�ˌq��;�O��"�r����7�̥��C��c��C=���y��$#gC�ؐ���Y����(T���U�{�/�NW�UЋ_W��H�lm�1եMͣ�]Ĝ��N9>���a���M�R��.��B����7�|Ӹ�N��Yt`S|:���*(hTQE��= (/�ѢX�8�g !������{L0��	Kd�g��駟�;���~hhh�;v���9��%���3$?U��r�ݽ1T^���G/�����+v���6v�[�
�/Qgz�DD`�N��I�ܹ��2s�H��|ҙ���x��*����z�9���x0Į�	��"�\2L�(z���=}0���"q�Kw�;н=��Ep�M�C2�.P��|+��n�FN��Hb�.c�����a�!3� ��U�r_7�oom�7�^K����g��o�h��[�v1Wwޤ1�Č��k�8#�qc�J�W[vu�\[�H��}wO�)=��ϕ���ĉa(���{II��^V���8��^�������5U�bs��i'�D1�,-�p�YG���7��O��
��@��mJ��N:x
2m,ܳd�@���r��q�#�����V���+t>z{,�UE,��ެ�Sg?#�s3������2'�0F���gBê���4<�b'l��A��'͐O�����>���t��W?̓
���g�wp(t�;��{�|�u�M<�XR��IΣ���k�8F����Jn�Pˣ�ǵ{�?pV�����-n�����8u���`"v����΂��Y���?��}�m���h,l��~:ڠ���g,Z�ՂO����w�W��O|�
���si
�)0J�%Z��8��� J���N�y�-����l=��v�㯭W�y�pX0����I�ֶ�a�%�����	+�]ϷeؕBf�7��ɩ�'�cJ�Yg�/��i���0y(��4��ކJ{Hd�������Ȍ�5�c���?� ������3����_����A��C�w��nxf�&>㊳�o�o�Af���?���ƕ'�H�o���S4�O�_q�|~�"�q)) �^�bq�䇟:�E��A>Gסz;��i|���4г'���L2n��3�+`�;���T@u-��� �In<�0	��	3v���;_��g�gj����1��+��9.��}!k�/�"C���A������J�̟�郯���{[���%���M�X0(���yp��	������Z5��oA��ҼV��Θ Ε�������l�N�]�.��5����۟ZG�~�G�h�� 3f���c8e�|4� 45�| �l�Kw��2�c�G�Qp����?�(\y�A�{�ʼ{�Pu��������W.=�����B��A��S?�{t�5�[�����c�lH�mz�_��8�B+3����7a�'����^�G}hi�8ΐ�����g.E��æs����Y���*4� s������r�e��g��#���xܜ����#�q���c̢�������^���
��x <�|�i�;\���C#�i<_����XH�N[W?|���ߞ[�U�<X��7�*�ЕL5����?	��=|7��'b%�nT�Q�$,JJ���'�<��~mjn��L���p���H�4u* �>�g5�_6	�{e|���p	���JeȂ�Z���1�y���> ?��i����Vn�#��#��??���n8�H���3�<XPAt�����1@C-W!�V���5̃C	��oC��MrИ���чυs�X��VpL9��	⸜�1��ڸ���-�z���u�������S���V��&A��w᣽�z8~u-����\������#o�xW��r�p�?�����T������?~�4�����3�n���\j�;D⿹���-,���.�d�h7Е��kO�׾����n�ߐk�@�'�J��#���\w�xf��}&�����.C�|�1�>V6�c�]0c��1c�PC�H�^��UL|�+��f��8 �}w+���)
����鳷?	,���|�b��WO��*����7��pT���:,�9.	�щ�A,>��+O�˸X������G�`�ax̠�l�25ť���Sn��{�El}�L���;]��F�(�b�f{�0��$� ?3��j�8�Ө����6h�	ظ���ֆ�r�����!��`T'W3	������ן�p>�$��}/ö]3ʒ9�8a+2\6k<��U'�Y,��~�����G�����pf��i�?��=aJ��^����mO��3��|��y�]4���8�(��;j����f��NAF�l����6W�DFՃyT5�yA��}�~��2�P�y��%O��� ��b<;��c$��=}��_?23F�ja���!�GaR]i�sYe�S��i�#��Y�8_$?�Hh��?��K�~Go��1s���/�v�y�q-�6��i�34�8r���p��SY�!��c�h�Л�ܺg�6CgFPA�q:$��<g�[�3���;s&���a��2p._�?�24ď�b��K�9P��w�D{{}+Op�h���p���9~��JB����#f=c�ӟxc��y}m���b��c	I���$ �;�j�2��#�n�F��^�Wð
��h���vR3OG��($�&��a��XgL��s�v��
����$�=0q�L%�2�����Vm��������Df@^��$�=�{`ٲ��K ��w/���S�d���?�
�i�s�V�[`[�&�nno���h�1��1乪9�Κ9���ٛ(8��1:�m�-9<��ID	�K�����E\�@q��?
�]w੬o��"�p�}y7?�b�]r���1E�����cf�W�솿VN����f�.c��񅹾8��o�%pWI7\���Nf�m~���u�8�*h[��ЕM33��4�xǷK��d�T�PYDp�9O�_q<������R���|^x�شi�����A#�����������W��x�-��5.��
3���KK������a�6f��(�7���A���	PWU����<���O���ȫkv�`2%f)�nN8h2��v>���b���tx���������3h�p�r,`���<��z�Ez�	&�W\'�x"L�<V�0c���Ʉ�-o`����ן{$|墣���>�p<��,��Y0c��B���%#�aȌ�[�����4�g��'�/��
lo�a�����SYƧ/p�sc�-<������O�_�Q@��_�~�ό�=l4���1��*���E<�gޣ#�{q����H��Dċ�}����n�	֯_�,>���N'Ŏ/��8�e��r>r�^�."ܹs)4�Y��0�ٔ�21="���G�:1oifnM<[1	�n8�$m�çO�Nf���G ΢ګN=~���|Sή�~���g��&���~60�o��)�Ӆ�q�Zl8�}f\yޱp��g�̽��{^��|�;a+�"�)��l�28���yN/2ӂ��s{�'=Ġ ��w�񙳙�~��©N�[:�ùm��BC���r�
�"1�]��Q��p8��|6�?��)p��Yp�'~��D��-�7·�H���?�gc��`!�5&H��gY'�W�{��y ��'hO
:N�c�q��;V��~Ĭ{��G���wЉ�
sp0An�ܹ<���+��.�c�=Z�7$�G�˳+x�p����R��#o�E�Gâ�p~�F8����D��d,[�c��q�ϒ	�����r���a��1p���͉�0;���%/-���~9�|�H��o�V�C�$8���ˏ�S�xh �w���?5���2o����z�qN�[%p
���t���7n���:
�8����uk���:Uǝ�'�y^?�?��ͅ���<�.��i%�mP:$�dE-��V��:7���~�|j3;Nc��O�.-;� �t+lٱ��������x�n��o)�2���n��~� N��/+/asm	��h��T�/���(�a�@�(���7o��������� �y���=�0|��ϼ�	�����������q������-мi+�	(//��s�Ñ�&��3��<+�C�t<*s�cnb0TY>{;
���_�|2s<��TY ��������)}�ʀk��S#�>�uGm�8m��~�dx��|���a�t�Í��쳭c �����z*߰s�Yg�u�]/�����+�>���@.��򜰬V/��v˟��폼�37�.;� �<����������m���^�7�5�5��U���B^\��~���T�&����<��ƂV�F ?��G���s<������w�Y�]����Y���!S�a��o>{\p��ݓ�|��w�|�"8�ƻ�?`kɒ%����ok����=Ӈ������/�)w梜�����xq܏kLG㔆�A^�.H��<�;Q� ZQ���ֺ��5����(|����!���L���ޜ�����pv��pB�����KG82�G#^��E�z�APLY*ƺ��;�k���(���p��O<Ⴡy�r�"��U8k��`��Alk�0UC!������ـ��^�x́�0�
������T8t���;{���:?o�X����8ۋS�,]��;��f�97�*U�G΀�Y|q��s�1?-He�Ӏ�{I������!XZ[[yL�-����H7��w�Z�Xk�8o��7p�$l�K����͝|=���J��M���.�vw ��ŀ��F��i=O������-�Q���\����sS�����wx ��ˎ�0�c�"��I0����u�0{�Xx�l�c}
��>K��;���v$�Z�����){��-qћ:���|���#�5�-��Ǐ���x��$�4T���.��P��л�����;��c*ç�1��w6�S!�=z\��GU �
���E�>��M�?��t!��� �[�[η#�22�C���)!���|�/��KW3q�̞���z�E%|�ٳ;�9o{�஥E�x�/}��@f�: �b&�!<L<�Y<�Eu'(&�_����Uu�����h%�X1��l��a�FnÎ�T_I�T_�ի8�����:�-�u�%p��q.�ԏ�����ݼ~�-' ��ï�������yE�p���1�3ɘ�������Z%�|d(!����A������@e��ӻSj�)���!]��d��R�I�q�r���N�{�z!G�C|m��V5�L���$,�)��-��q'ԲXX\K��1f�.P6@���3����;�/���؛j��d�x6�x�X�e�sus7��ܦ��pQ�������Q���2�t8�ÈMS�����I�b�*�\ѵ�;�LA�JR*�P�ʧ�q4�2I���Or"`�AF���T��-GAÍ^��%��J$J�Som����(�:Ό�׮�ᒁ��;�\Z;��?d�$�5�V�3�ΦO����#O�)��`[c�b�"jQgm����Yd��n�օ��M�%�S���~
<N�/��n �݂���U�;W��� �}���:�ꁪ���gORC��洪��[�w�y�gς8I+�2*���_�|�˸o�b�P$`4��"�Rtg��m��xp}�����8]/|�9�8[/p�G���9x���P�$c�Wnv.b�H
�ڶh�w`!�KV�B���K�P���xq^@�&uh�����p���hQi��ϧ�7���j���.8�0���a�m%|bs����0���mrq$
��Ǚ���/��
����uPJ��]�S<Y�h"1R	Q�2R� YG.:Μ
�ç���1����=��T9L�5�:q��^��dEGFG�� L`��*����UPZ��<�9���N,yN���8�;;��ut��ڟ!�����Y�y�H���[(��/҄�+��T9`����Pj���!��UU�|�pYY�4�#���̧r��Ō�J�����F8xRB~p���5��H��}�8��� �F�hr����jT����.�Hw�]�D3f̚=��Aۨj γ1���`͚5�l�\�D88�={�l��i�J��rg���y��J����y��<aO]@x�ҷe�.tuC;���(���Y'���x� ��D̘1�E�1(bƹ���IH��:x��ȠQ����'��s���{�S�!	��{��%2tܸq0~�x_f�%-͜�I�&񵌖�f�Y,�9��S޷�g��8�jjꠎ�E,���,��g��{�����@���5v	�����A�T����e���q�J&=u�u�{��ɹV��P=555�g����<����ضZ[����w����#����!�|uv]]-TTT3fs�����^V�ou^ ˗-�'��gz�A8U,(+--�DK������5q�[��~p2$���$|]xm��Ę!�@�IF�Q�^h[v2� ��Q>�}cHEE�X����I�ݼh�KSP�UVt�T� �,���I�����I3���j������d���� 8�)�M&L��mͼ^{G'�fy�T���9�8:��;��S�B�E� 	3���A�㙹apd��[�^2��G�,澗�z�5z��͆H�����X�:��ނ�>'�^be�#	r���YJSEŋ`FSi�O)��\#��jS2��LG��,;ϭ��@IGw�|�(g]i���MxX�{#u�$�<j�}aPV� ��w��T�\�
��s��g�%�f�p���~woo���`a�k}}}N���.�Eh�x�.N����7�1��V������n`٧��C�8x3N_������w�������t2?���Lj�^qI)�f�F,�'���wH./����f�3g~p"�c�LC"�(8�	q��mW޻}Qz;�@�6�.��g���������_2��Z�S�}�h5`;�=�H�ݶ�w���§��0;�������r8�wCww�|��0�gg�~�b��D���Ͱ�h�mڎ�b��B���QR*ъ��[S=��3��K	z��P�i��ͷ��R���X}M�5g��Np�L���X �!Ȟ��'��:���N����y�0u�&��3���8~y"�בb�D;q���p����?����`_ǎ��/���DM��T�E�eu���D�����~�d}U����C72�u"N����d:CLk�_��<��Ox���	��Ĳ(S]4��wVq�/���aX4߀mQv޾����g�l�������8�����Z����c���b��4V�r[[wo��/�����D���;xÍZ]�aW1?�s�K҂!�T��u�1�Q�^z	ݸeK��qܣL�,�>���G.��w�x���!�d2dv__o��q��3l�x����������<rGCCCI>���Ι��F�c��g0,/����W�ylӸ����ݑ�8�ڂ3��I�0��@��t���������θ� ��>��T��N<h2<���41}H��
������2�$�����N�M�!�g�=p���jՒ=
�,8�S��� 8L�l��O����G��w���p��o۶50i�w�uv��v����'�aXKGϰ���8���a��5���O��߹����"0�-Y�Q����d�+P"RxB��r$|�O��|��G�����v��Ȥӑ����?�r{Z���q��ų�F2�t�}w'̚6F��_~R}�g�������!�X�ϐ}��g�>V�3d+��������~��ce?C����!�X�ϐ}��g�>V�3d+��������~��ce?C����!�X�ϐ}��g�>V�3d+��������~��ce?C����!�X�ϐ}����c;����##W�7��ˈ�3�m+nr$v&Q����M.�y4�(o���;Z#b�Gp�����	��eY䝐�<���@��˲6�c���*�{u"+�@i��,�n���.�C�<Ě��ͪq�t F�#�M�Dr���5+<�Ʋ���2����`�������C���e��l,�dw23�Z$�n<�X��w���[wv�h���!H���2<���`�bUTT���-+�Gƌ�ƍ�����)uļP8	F���"F��	zDeu��ǘ�XQ<z}_�� ?�7��M��;�������:�L}��uDIi�DvkG4�����_����F��_�9-�{� �    IEND�B`�PK
     $s�[�ة� � /   images/8f771a2d-db90-4bfd-8b3e-8d66edcda07a.png�PNG

   IHDR   �  w   `�3�   sRGB ���    IDATx^�}xT���{��T���DE,�"��

XP)ҋ��.ދ���k�^D�B�bQA@��zKoSO�����0�7���y9��>{�{�w��῟��@	3��wV�;%����_\�8���Q����O?� �9r���[P);3���qڣ���%�mݢ�!����f�Gnnn���|��펳Z����Yv�=�cǎ�����Q��l��wϙ3����|�^U�ӄԩS3`�Zm�+WFFFrrr�Ç�q���~���o�fV���f<�ࣻ���fK�,��p�¾?�����BzO��yN�uH�EQ��<,�^�@o۶�;]�t����O�,�wD�����:u��g���5j��F����F||<� �n74M��b 9y�$֬Y��3?�(����^0dy�'%R�>|x��S����`�k }����~o���G��5~���Wi��#5����z���Z��xM��U����"Pa�[�v{��4o����p����X,6x�n�]�z�@3���������Ҽ��q̈́	:���K|>�ǒu8�1��e��4M���Oo��$���͛�ְ��iU�&���>n����� a@@�KC��os��8�i��c���x������C�L�4���c�/�w�qǏ�7onZ�H��$IN����ݻ�;w�"���=�c��m���bذ!|�>����C~^!lvt]��a�8�s�<�g�hÖ-���#����8��O���֓V��ׯ_�j֬Y��RB�e�����E������}����|�g����}�-��g� #�4�~?H�(x�l�,�2��!>.���ߩ�y�ũS���ZNڅ�ްaCԝwޙ�q-$�g$?!#��Isйs�W?�䓱�����*۪�a?����C�ݷ�w���2�� &&��DE![�
��w�4(��4	A#��o�y��'NG���Y��ʂ��4y��^��0ܫ���J��� ��n�?����z�(���&L�wԨQ?_��/s�5Ɓ,u�xRS��?@��MS�ωlW�N��H��K����&JQT�\��f��x��^~�^�	��իW�G�������(i�d���Fk�O?�dmٲ%��~�	0�m�|-ǡ�����1P��PT?{9r?�v;��5�Y�W�!�y<X-vH��S'O���׍=�����q	O�5jI�8�[BFgq�_�G]�.��l�	n��_v���<��(QRG��6l�w�]w����u�Z�2�>7,	���@"�dZ����oUNgR�����fs���3�����e_WoժՉ�zn)n�Z�j ���q�8"噄@@�A(V܆Y�vm�{��P)�\�K".1jԬ��e�{n�4i
��A�UU�� [H�+,Aa`sB�)�40B*�|����i�rv�$�M�a�;1|�h=z������R�F.3f̰q��M*~Kq�"R��燤=�~��$$5j׮���={�/��xiD��q��w��8��߿GժU�q���7�X�/i|(M�n�����
�=hذ��g��.P9����������عs���o�7�+���ѣ���Nӧ�D���4}Up"C�� 0B;'�H� B�t���>��#FM��:��,Z��Y�N�~�����ҳ���>��È��8��-�/4iҘ�L#��wd�Z���!�!�Y�7�c,�d�]��6��Ė���Z�Z��?<R��a��U��sy�/1`l۶�r�[ۺ�7�岳!��p�~�v��&�$�V��K���=L�\�&���b��~�?��2Lw�/� �[ψ=h֜�&�9~�o��GNN&����Gr�%F(d�g�Ġ��iԊ�S������no׮��H,�o��fkҤ��������Y�hQ���~��p��7b��޽�7�ȵ~��B9�j���)���(�Bh�L����p9���3]��f�^�����Y�f�ٯ_��ɨ&uY>!���C�N��V$�1`�~{��Ov|�A��]���I#���C_q�A�P��^7ȥ3�᰻0c�l��������#������6m�4RY��s��w��/�D�m�08�E���4���9Z,
}_K�<�1����� D����^�W_}m��u"���?���/���?3���ǉ��]���8�g$%%:y�d�+�S��Gڏ?~�רY��@�$��敮��8��(6B��c�;��O���q��K�n���Z�DJ�hů)��A�UD����k��U�AF�(�0��0p& ���n���.ɦ*�bԭ[�����7$IU$�c�X@��s3Q`lܸ�OH�g�`F o��j��U08��OCӵ� #111-##���H������.kD��s���$��^�;\�(�%C�xԪUO�`Ȳ|6qV$����aG;3�OĀA����xR!`��k��4'|PRQjZB��u�͛6��q�� ��J�YQ��R��C(��o�q�n��]��pqĀA6Fz���G�O��BU�,���Q�Z]}��b��΂p'����<��<.�GO�^��|�@�7��D�l��{%g���Aң�u��_ׯInڴuF�� ��y�ru!��R?��䢟W�\�ܦM�ӥ~�%.��� U����')! ��VWR%l�ѐ�p�s!�J�6v�J��ur��|���ڵ;Sn�A�����<1���awX���آ�///111����Lbs��!F��*f�~6�A�gO�R��dfr��)�|A)ϞEn�M76P���?�!-�	EQUU5"��p�R��K�,I�ر��p�1���������M#�@�Ofv��J����$U��p�٪,������M՟U�^[�LZqJC�Ob��@�.A�qK�����[ظM�6�Ý0ATM��-0>����~��7@Ā���C�x�UfR���e���366��<t�FLBQD"򒔠�UU��(Gt�b0(��Y�F��#Ӈ}/Gd��w��w�;}Z���<60x��t]�˃)	��qݮ]��wDD�J?����@��*��?����@���K+�� ����l6dg�2U2�(m��/y�kT-r7�SR�s�\��H͚�����F�N��1�	���r��>��N�n��� I����<1�i7��3gƏ����A�XHPp��8��g8��7�STT�QEݣ��T@���Sy>ǒ��)q$&U�ȑ��=
zA��C���#:t��}E��Q^���ϬY�����gO��1`��������TQ�YK�w�yk׮Ug������nI�
�T��oѢ�Gg22�����n����'�|jr˖͹|��s�l�H�ጢ��8��^�38M��' F��m�-[6cݺ��{�v���$�R�<����}�W�疄;a!�Q�As����7z�6���I��G��P?۩�Mݵs��l�j�q�$IH��U�=/�����s_?nB������J��0 k8��p�4�j�"UU;�����O�����g�.���0;�x��<����ڥ����p',����
�㭷�j4hР��1����S��jI�+�3{�n��X�tI%�q��F�
{�zv����1�m�'���z���G"ٖ*�o�s ��ahX��c>۶��"w�Ac�Y���i<��S/0�����(�z�:uj�!C��]�Q�q��>��G8�}��4l߾˗-��{K 9����f��N�}���?|�_��'�fø�Z �E�>A��A�k���i�9���';>9x��ԷK��+\Ì�<'��I���z��������x�,0�n�+��&���.T�{o��Y3gM�R�R%��C��<x����_�J/gF "�V):�(<��3���cC�84|�r	���3y��&Æ+���������-_��2�q�T���skv��s��e_}���UwO�>�:Wf\��`#��g���f֊�����g��v��:h�ЩW[)~_.�R''Nl:r���J�����I� 0v�ޗ��˓�Ԋ�E��_�<}���U��^_����2f�k���{��� �w��NZ^v'�v�zdL��ao�;a!�3Ϲ&�7n\�1cƄݰ�cǎ]ǖ/[U�r��f횪m����oV}튣�4�^��x`ەf�0�E��̢ş 5u�1��	J�E>{t�V�=���!#�]�y��}���q�;��رc���=��c۶��Ƹ�($��Æ��vΜ>��ҥ_v��}gi^��� �WK�ʻ���<�n��Ç�~�4���h|��<f̘�ƍ+��z%۶m߳��k�]j��ΝyO�^}�=x`�QQWbb�/]��i��(�"��8�/Y��c>u�K�WB�7��ѿ� 4iz���^~�4������G�~�7�X�{F^�\��رk��e��_r�<'�ӽk�_�.]�c��A=E)u��0n��-�ؒ�:�UBÉ��F��zuԈW"�̬\���� �dĈ�O�0�r�����<Ǵi3�׶]�V,_}kIݰ�*w��2��� Y�}���ƍ����RK�b�aT pp��ѩ�C��(�؝�ӻ�i�ⵡCG���Ͻ�udD�����gqp����O���_����>���AΧ	��" `l�sǟ+���Q}z���zFfF�ys�=u�L�[n�m����7k��di�e���E�>��� ������4����CGF�)WR<�9z��r�С�Ǔ�-0�6��������Z��G���Q�R��^ ]-�d>F	q�H����CL��_~��q��}QڍuI���I����].[��D���~\ӽv��N��qƌ���:&�0j,Z�ɾԡ���e㵾>$5ƌS~�����v���pv�ؽm�ҕ%�����{��*�U�~��ϗ|qw��OP$�L�0l�/؟�:�ʶ��+9?�y-$F�x/��I6v��'ǎ[>$F���aڇ3���]�X�u��f�������=~��EE��:uo^r`������2�~Ptѧ֧tg���������[��_���:��w�dc��m�_+V����4y�i����`��M�9|�U�jի:�g����R�h~�=�K	w�l]Iy�}������[�=�2�a}"��� ���wo]�l�m%�����uú~�Q���pK���i�jպ�2�E��9$u��K��=-Ǧ��;��q�D+/��!`��	M�8������0�������t?����.��ֻصk��W�hc �,]����7�K�wc��_�\s�}��wUD֏>�3r��a6o��1�B�b�Յ�={����2|��s%�`�.�y�n�<yr�aÆ��x>�C;rd?O�������y�`��?��\��D`ԯ��':�?���/��E�uz��#G��q5���'�SG�6��A�'}hQW�=(�v��Ç�5�.~��`�6lX�l�������-VʄӉ &O��CiǶ|�տ�(iAޛ���o�1a�/������K��3kN��K�<��y>��:4uȔ�;����0�8��Z��֭Z?�ਡCGN����S�ޗ���C�����1����<eE�k��c0s�ll�c�����X9�^�݀����6�8�`Z���K�X����Ͽ����0�դ!X���ܹ+�<��!/}'��-o�Bxʔ):�8*a}"*1����H$\�X��w�ï�7;~½X�����~�b��<��EQ�2�߉����)o/�ۧo�Z�R��1}v���ռy3���ʈi���LFe.g,�~��wx|�K/�%^ހq�<M�2���C��)��]x}ĀA�۶m�mv	v�����ǫc'�b��i�$��0���z�s�<�X�_~�ن��@cd�Ra��L�d��:B�u5��e�&��塨��U��� 2p�';>?`��iaOX96>i3L�2�Mjjꪰ�3���'c۶M��i9[�XXX��>��3�|�]%�B��t�&՜R-�E����c�[X���73 ��q����b�@�Ջ��nʞI�c���<���ܩs�^tU�����w�ԩ�<��p�5�����U�Āa&u��y�5d���h�i�2�X3@�=�ݏ�\'{'RT�j�������zj��	p$u��%;;��H�(�y��=�g�v�3`���aOX9�4��&M*_���Wټe�b�d���O{�R���_꜏��z�y�ŗ�R�5�Cq�?�>���лG��)o�$�����6��9s�4�իW�) ���-���Z�k�j�$S�0}�=���c�����f�۳}>_\y�|��W�Q\�}��߸ظ�$�t�ڃ�6I}�ǳ}¦���ƦԸ�(�pUT8�Ƽy���ѣ�ԮR�͛��#0Z�h��y���]��\�н			����5�Ks�c̝;�0���}�[j����i���'Llױcװ?����O���>���&���G5|��g�OQ���0�Cc�?d^+��2�ju�����}�f�=���p%F���w=z���s�� ��%>o޼[�u�=�����ʀ�e=K6��(�� ����Ξ5�y۶���Z�jmIOO?K#(O�������t��5�S��� �-�ܒ�`���>��pwRJJʟ�� �Ǘ���.�ܹso�֭[��|E�ܼ�W>&&��0��'s�����f�c;�IV���ڲ����m����M��������7т�7τ�{���������Z>))"ˉ�,�M���tE�x�+#**��հ|���k�Dغ�~����oߞj�^�-�B�,C�r�-[�Ү]��|���>��/LnӶ�����A�ʕ@�hGQ��o�vg
���~�x�W�o֤�'͚5+����2eJ�S�Nݵ`��������~5ϋ�=�B �!�}��լYs~�V���i����~O$TI�(���U�Vag���`	 ��#"��hP����G�k�%�a�;Шѝ8r8�D��޻o=�⋃�o֬Uɱs�	��h���W;����c1�~��փ�j�<l`�l��_Y���&���#��S�Wj�|��q�>nu6 I�}
q?w�֣_�^��-�4o�|��u����Syb���1gΜF�z���xF�� ���u?H�j�`ioE	��f?o�eUM�5�w���q��j&�DA���r�4���=��9-ݬY�U7n|(t�fy�!p�XB��C�={�m�{��j�$l`p<�_~�ILL� "�P�zz�݅p8,������g���i�H����н{�2s"�5k�͆Z��-n��U�D�zqW�Ч�L��80Hb���wR��1)ap:$�`?��:-Ag���:gSp��������Bآ��`
��Cw�o�����<�SUU���`MT�x��~}���ի�Oe]��͛�Y�~�D	�1%O $Y8�lg^b�GzW�.�/�K�����dw����82{�y���OY�`AXnk��X���*��W��P^�Q.'t��M���0�'��h���5�n.1���ϡ���5�Ŋ��|n/��a9tb#G�R�WDH�x��'�u������\�s_�V�|�����0Lmi�/��T�KN�����4jamv�g�Xb��Bw���i�?����u�,@x�st@�yS�P:.��"�Y	�|���7wV�=�\u}I���E����u��uo@~~>4��d������u<x]�fpP8��P6���<	ɠ��A{�7t��59����P���;#��bpyZF�#�Η�e6̦��:u:գ{ϧz���KY%F�ƍ�n��G��v�MEe�PD:-�j���1���j�v� U���<��¤����S�<��L�С�������`H4�d���t
I�i�f��e.�K��������Pc��82���m��Tp^/$��|����`o�g��N,�$�e� �_:��O�""�*&���!(*�6<
��В�^�	DAVt]����]�&Nh=d���-�    IDAT�2���/ؽgwGQ 8�S5�#IGKK6�G�K��j*D���غ� 5:?����)�������N"~/;���(�=��^�Q����A�<$��L�X,���q��7x��wS>��0��&���*z�&��f�To@����D#!�Hz{��Ӑ��H@���;k�p�:���q��t� ��d�0x��^S��t������n��%��э<Y���~��_����Ӡ�.r��A�:�H��,�TU�+J@�9f亲J��^�f������\�5�U7>| ��!)?lZ�W�,�x�s�Y�r�<�{Հ:��!c"�q�J_}��a���`���'�<u�I��+Ȃ�^�=z�8\�g|��MU5Оӵ�Nٹ����{�����w]�y���-��Z�	K��4�W�/������ۇ32��[�4v`������7���~P�����}w޼Gd�RU���:u\_�'~�paM^Ѻ@Ӣ]V׷�;?vaMY���׮[�.aǾ}�d����W�7���6���/[�]��ӧV �LF���{�>�ǔ��H\��J�y��!\�k��n�˖�h�G��ջr��4֯���6:�x�36|�!i��_��،�{���ۧO��J�]_����g2�À��o��ݻ��*��\K�,��
�
<_CPſ8C�ҩ_��ҾȂ��|޶"'9UE�Q����رc�Tڧ\��~�駺���<� ��Ͽ�W�>�.��zŊvY��|(R%v%��սw�!�~���o�W_�hV�{��E�*�
6��c�^����p�����qQ�D��/�ce��K�A�������Оm��ȯ�>��ҳ_�+�Kײ��������5T�iH��=�u�;��"`,��v�����G��������/9k�
:Tj0{J��v�Z��ٰ�3�>>�}�բ�A3`�5����
����4�7��p�Lv�.�8������MR+�$�J���Q8��Y7l��;aŚ������n%�7�vc�|7sٸ^� ɀ_�^�"�͵ Bc��2vrn��Qg燆K.��6�e��8��q����'�`�P!@�����%�]K�0
 �T��*/��ƥ����״w�Nl����Zx�4}����Ϗ�Ӡ�`AqT�ϯR�(���$�ǥ#��̀̖Yԇ�3x�ӫP�3�=` �a�7�0�z�	�^X�BX9�z>�f�����C���z�r9�x���h��6��dCҼ�9+�h�Ek��T`��pR���b��'��(ˮd�q�� ݏ���,t��j����3X�������D��@��d� �;)��FvV��\P��l�~�9�cpp^��<��x]r4��~<M�Y����ռ͵S�����
̟��ݻw�<0ޝ��-S_�v���P��	������,5���ag�G$`���)�dx��\ �7V�Q�Q �QQ�!���O�YRe(�D�dȺ
Q7�S6��048�3hR;����'9pZ�×;�ڪ��)v��%�GY����jX0�p��Bw �.�~��ڶS��`N��؜��">Am5� :�����,B���e�F5QK8
��^�"ÈÊ�~d���t�5Oof[.�fˀ�~�Z�OKu�{T�+c��/�>�:n��/ME�AV�ΉP8X��#����A�q~��5��`#  ���*�$�����܇�MSPݞ�?V]�ۚ��Ȕ� �S�g��u�C'"�}��lF�&5�,d��灂��B%,�\��&��P٠����%�.J֕u&/q��S� ������Ѭ�7X���g��ia+��
��*��ES ��L2�^Ӡ�}H�q"��A<Ҩ:�[OB���W�ě0{}6|Q)�4v�,��K�ZOL�4�P���v�<��ilx�Eϼ�^y�G�g΋_�Jfު�������D����P��`a�AF5��T
tP8�iӿ(�I�<|>�6z�A�i\��i8�L��|>����@!`���kL�@#U"�eAjZsp{e�����9;��qX���ZL�HꄀA�i!����er+e�$�z����&խ��zq|]�i.	k��pFLF�Oa�sp���$��9�p�����[+�����N�#����N��+�m ��䎧���~��%�B���OJ�����������6/����E��={Ƀ��NX�腩���[jU @7ll�%䁇�T�����l�18PF��1�	�(�I4����"��\�unk|�=��$��ieع�"�M�^��@:n��D�	�x1G��ܜ_l-s�P�CXg�I����s�.Us_���
��	~<و5�}�7I�Ѳ�6���CF��DW,D^���s���n���!p>�Π�mUPۻ5��TD�`�"d[��[�4��&�I�h�.CV
�80غ�Ll���;a�#={v>��t0f�Z�p���n:|��1l�0`a*BD�	�� ��*g1�Xp� �1���*��t�ixjș�R�Y�4�K���2�d ��|��^f|��eK I\&�ֲ#Œ9��"!�R37�3`�]5S�����'p�|(f� އ�!rH>Ս(;�7w�p�."Yr#`�8��aͩ֜ �Rͤ�e�e�9� 
rϤ㑆5�,:�齰آq	�<M�i>�)�8�G���)0�MC�B$�$=�z�?��W:�����7P���={q��C'���p�&��mD6��a�TN�a2C�O����~�O�*,P�fãk��t
.-$d���d/�!� g(�y*�l���"U�U�"���Y�XT�A����SBe|��-�6���WMPi����Ptd��	�l�m�5������I~ȆV_��D�f���(��%$�߇x��cػ��{���4���adg�#w���x�@&�D�K�x��L�"4���|�\!D�2ȋKR%�F6�;00cʨ���~���c�O�:~�m/MC��Bfr�&ь�|���Ř����)h�x�ᇖum暴:�I8�<�	�E��I�i������Pfk8uրѼw׍F%.N=���W�6���fv�DImJM��P�4��d(A�a�>�>��n�}�Mc`1����<%�,��qB@&��U�E�P�)��B<�Z���Ƨ{`�T�e�Ík�9.5��!OL��=
2�ds�v�;V�#���w0Hb�?@����Ǟ���N ��9s>}�W��5���I8��B�m�?�	8�.�(��2n�2`W��ʒ+c�N�be�Ĵ�� �����	J�k�)yH�4��*8+� ��I�flV�ť�
/d=@���Z�2��`��xxM���p��OH����X�C�;��r��--����$�L��U4�'�J�D1q%��@�!���:�ȧ��1�.[�h�\��dG� ���ץwX��=q�ރ&|_`АhǙ1K�Ee�4�
��:o�����[�POΆ-��$K���Ґ-U��ӵ"� ��7$��%�V5��hYǅ�ȁ���c�8�%��:ѵ�k^	NO�3D� �L��9Ywu�0���X�O�X�&�}�j:p�%�� ֑�'cE�'�
P��Kୌ�G�Q��e�.75���r6��<�A�#&��]f���	A����c��3&��peU2w�=}�L�����@M���IT��`![�@�ø�^<�Z
adC��,1��8^F���Z���x(��Z���	�[;
��I؍"�u	'��E�u��j���Ef1�X[# S���b&�9�dw�{�`r����uS}Q�-�wMj�q�%��B��dc|y؎z<�������E�I�2j o�Ew�Qt�T5�\��|fwe��h�$_7
(��Td�򈗐��Ft�ߧ�y- /�J�-����	�J�R2�̙�	�;��2������8���r����R@�d�I�|��,.
q>TĲ�dՋ�*��~���B��qH�2`3<̨���ٶ�j  ��R�H�1�y�Q�Ȧ`��d�0(8Dn��CL���hp��@���v1�<����0��Z< 
pY�HT֠��rKdWɰ��H�D��$��{�y���� �f��d�yJIP@0|`̜2�}�^].�̘��Y�ԉ��!�q��ʃ�,<nS�2
P�����]�b�aQ��p��q_��q�5����p�̟��nX9-N#��3h^'1�2�1;$�sa�_��WE����&XX��h��f<�Du$#L/Ō��%�j vUA�����n4��D�vN��z��-�.� '�x��pN�"y'
�ɧNƔ,�ֳp}`?�׉��y�������F���\��Xn���,/�*	L�<�]�ޝ�)�P/�e��I���Y�� �K��^��@⑋$1��D��C�����
��ێ����F�I�
q��k^8�'�N#��E��ʰi�� �x8	[��F�%G�X�qq�	���a�ɞСD�%����xY�J��̸6�t*��H��T�P�fl�hf����9�v�8N*�#�E>�S܅t	Ezu?����I�֎஺� �����]�a�_���%�p��X(���+�;��ݾ�*�O{sD���v>��*�I%��&�t��/X�>��
�+jp'����K�����v�, ��ع� ��$��
N�p�I o�M����A�x��>��^/VC6���9�޳yB"�
�q�KD���,-M:s%�JsC\%,�n+�<%�6�	�Cn�QTP�lT���J���J���a��ȓ�q���l>	�`8�z.�	'���D��׫	���zX(��=;w�P�����l�\]�*X@��cƔ�����z�B�5�=􍵥Q%�n�0H���J�l��jR�tT�N Z�G��
��Ǳ2 Y���8�o?ܖDj⸞�B>T�#�^Dk�P�rqȀ�{P/����B�ს���w?��x�����l�3CN��MPĆ*���5-x� �1�Ӕ�3�gh�	Z&�!��CB�D'Tbӡ�طk7r�
8 �A��*|�Cr1�ȡ�A���͓=��[릀d��|�MSpx�.��8�R�%WEg�*;�+�JJ7�KI��F>ҿO��*�K�-���Si�A♀!�b1�� ��R�ս�P�?�
�Rb�
	0vI��c׶��X+ ]���Z�Hd,���A� �\��SvW�zU�-<�AG>�ٱ�rҬ7�W	�A�������t2�Y�$�wYt��O���JPO���	�q
�, 6>1�Xr�34���i��b�Ǹ���E���C��VO�&lEU�l����]Y�X���0�8u� 
�(��5pqڰ  X!�Ac�ظ0|�'oۿw���y/��E��2����:a�5�Ґ����ֲp=w �����e�*��Ʊ�����b�mIB�X�M�1�`񞢍\��O Vˆ�/D�]��1��,X� �@H@�\��J�墡2�>
�P�8(n)�C#����$`�� �3.p��;����y�KR�& ��"���"଎��M����x&m.%5�������.@��
��g�_!Z8(��Э�qT����y�D]�wF�<:.�)#�����
��2���q�"�\ɔ�<�z*�Q��D��	Y�5��a��ԣ��X�� O;������n J+Dd"^?�R�.��J�j`9���9\s՘���LM�j#{B�$Wp�,	hL[�7���B���r%\B��(-Ս$Y�2�`�=L��aJ�:�h��r2v�7���}�5�O�`��HN2�I���� t�
��"�"B��`3#�(�C�gz��R��_�i���y�O���\KP%���3xⷥ�̖���6����b�\�QT4����C�2CNg�$�yEt1c,���((�bK�C F� Q�De�y����7��O�㑉8G%��l�G�|�o�7(��_P��>~�� 0(�J�ÃX�q�A�����r47
��P9R2���#Q�8��<;�E��9�粑�d#F)��zap*
y�(��y|e�u�c��^�"��3	M��\
�'�x����U�څ����ɔ�P������%�b�T�ID#��P�N��E���#V�i!���@�cF��(Z����z�*�� ��A�%Nd�"2����	.慈z �N�W~�̤���	!�,Ŭ�p��<q �Q�V�d��Di� �?'�,Ց%V�1n8 ��ⳢW�%�r�0�hxPA�GIX��*"��"W�J�C��g�.X5�F~��&�W�J�3��|�_�N���D�a��A"�>2���5DX(�3�6
@|#����>Ί3���E|���B�c)`F�V�l��P�;�h#���xx��=�qG=y#Vv��{a��O��8�$�)._�b�՟���\D09�S(;T8}6G,�8'�C��yP�So"F;�.Y��Q�UA6�\Qf�c�Xx�� ���p#^�K��r!n(�LE@�T��_wBlP8sCR�+L��h曣Z����o�a60B�$��8/��S�iXN�v���w�D�</1�ߓȿ�
7��PԒ�G	&����w�D\�I�p��T��
�*�B6���)n5>�r*�gn+��I�au
:qY��>�8����,��h��3@@4�i<}����PMB�_$;G�fD��)^��+�����L"��^h���[0��Ʈ��ޗ@m�,��%TI��)#�������T	�n�:�k~Uq�!�Ɣ<�f)�[�f����j~'��*�A����J�'��0��M��")��4c�S�M1�����b�Q*��T���O�U7��K���)v�j9H�PS������:���l�I��Kę�!�[�&��O�g���ĩ5`���X�I?"�L ��p�jR�M�Px��4�0
gLu��Ϝ�K�"`̜��}}���]i�ϫFH\� �2�A��ԇ��E�uZ�ц� bfA2���u�x��-�i��]yX���D�&�����G�>ˢ�-Dϗ0T�m~�n�S��<�M��lA��LRP��0���Z(dM�8���������ER���N�J�z&U�E�
�XT���>V�
�(�Kd��P�Sb���d�I�!)Uz���p���=׻�y}a�1�.1.�=�	�ҍ��O�ʙGA�.Q��t�\]&^C��ГMB�nLI�ؙ���3��$�M@�I:���E���EH�9骠B�I2PB��`V�A�l?����`?��9�	��榝����0LC��-:e�%O�ĢQ� :EF���u�L����<��L�G�����GX��3糖�R���ZK�� !~��!���jHE��r�`�`�K#MF`*��L��,1����S_+�5�P<�]0������8R%",:-��efw	�n���f�	$�:Ȟ0�c����]$�B@2�"m '��<|��2�i����I�h���B� �Fz�ٔ�W�q)`�|sx��}��w*R�!���WeE7,��C��eC�QsK���䇹8t�?Ȁ�L�ܽ�f>�/��z�b�,xƧ3%G�z��!	�<#b���vס0��R��l�B��ԓd��,Cv��f�Dd���!����ef��]�%� �jp�wa�$�Qy,}�$4�b,yY�\OX��=�,I����b%���6	3dh��GKOM^h�L����G����Aכ��4f�hSi'kP�B&E8�O�a0�N�3$�qd]�dҘ�& O��Az��S)��RL2���D\�c�71�S�i��)�F�2�`�X�(T'V��\~z7��[K�˜ky>f�8Q
B��C2����Ye`p�׹���f�y�?L���'uB�k�03J)k��):J\��]4���Dxyy$h�H��b2��w��n�p�Z�q��)d����u���<���X�����,j�����=[��$�.�."c����H5���)�,�m5�M����yS�7X�g�q���    IDATY��[$%He�$#�?��x����Q�N%�f��2�fRހKD`eQ�57������I�DX�S�fr����\��h����H���o(��D�Y�{��{�0J���O�\�����4v`�����2���Dp����� ��F�IƧPX[I�����x�dl�lA�,��U�(«i����A���̳,+5��9dW
�E�P�EP�U�WĈ;D)��l,��nS�EX}��aJ�ZJ��Tc�����\K`�3>HD�@��E����Ɂ�^)D����x!Zm���q�𞝈r8 �����B�nP�Z����,�I"��� I���U��<���N!KqB���SY�������� @��6<���E�� ��^�����VxM@�G�jq��9�āW}�{���,Yf�Vd{4X]ь;"
T�\�(*E���?-�@�s~�,V�����,9mGAn&��(�UEIY�����Y�vfԒ4
�|��oƅ����eIb8H��¢	�p�0����`�ZqKEoiƴ(#�[�P��ϗ��e��A���.� dʲz�����፞�3�%G����r�gǬ��bh�yt8�R���F�V<�
�@���En���Hĳ0�����Ywb�b��GMn5p�RC��dd4�Y��$B��rq.|n�K�/�2�
�� �8Y5��"�lV��d��{�s�B�0x>�� C�,a��K���1����
�����E��IEH_Nzg���.����b7�5f|�?m�^��n�d��b����W��q�v�(�Ω���1�V(�^;Y;bccQ%�@�u�fW�T;�v~O!��*^�lD1���!�TJ�~�� ��摗uN9 �+
^)�-��B8�S��T�0�����8��6SU�;y芟5!�a؝.x��@S�QV��L�-"
�

Ir	؜�,E�\N�șR�^r���Q,֤�JJ%,Ui`�8���
fX=�.� VMi�Ç���w�m1h�aܰ����1���84QB�Chz�c��Ŵ���K�GBl|~�%�� wUv��7�_v`���3U� �a@��E�
��,4���)UY��[�%������%���w۟�S�F4��d�1��w/~>�°&!ʯ�)�y/��T�W$��!�;��l�����=����x#*D;p��l�{
�WLA��V<��N<vo\9*�������n'���m�j\)�D3�-�J�r�0fLu�C�euWM	q�D�B��Îe���t�M⾐s ���()B��_Ʌ�����`��u�~@v�p�F�8?���	����F��Jl��u_������ϻ�骓X�t�
7�M�iYb�?������a�kϠq2��$D�!��� �}�dWn���t���7�Ѩ�y����E;�y��EeK�"F����|&�N��'�2��0C��fY��B �P�����X�����jX��wtz�.8�砟���Q�6%(C�H�F�M��1"�ŅP����80��4|5�-N�00��5�v4�W�Zj+|�� ��}���Z�g������ı"	~���@$(��{�(^{�-Z��ؑ�����K$���3d�cd����6#����i��倡/<��7CF|��X4m�Þ�A�xb�WP�D���O�6h|+��W(�p�՗�⦚@�^�#�H��CŊNp�
�'�%�x�ջ�y/��;+� �ŏ����V��	�!W�A�D'>x;����a�����-&VI�S[%v��b�b6� �,�.aE>Kgc�,c��A�_��o��8���K8��,�O���CX>�N����1	I�����������l�j���д��7ǰৃ��*�X �6IE���x�#��>s/�+�jg���شu?gb�,x�n��q���
bB-���D�1��Ag|�u:f~���6�˝+����ps�
��A��1�B-L|�l�y��	��#F.D�\�A0�������hy0x�R��p�Y�:��l$�|���{�ɗ�h�AԬV	s�ނ�Na��D�D���[�)(�e�II�X�p�ˋ�T�I1�s�B��m��,LO1�m��Wy$���ހ�cּťf���.��d�h3�q�DMg�J��N3���B�=���"��Cg� Uv�A��q/݅� P�$8�X0a�/ظ�(��ZX+�Ч���vR�ɦ)�/4��y*w��O��~���20k�T����6��H�y�� � o���G>ޜ�5�5o��g�`��?�L;ܼNA�uQ�tޙ�֦y`�;�Ψ��(;_~�	�v�+>��g�ʨ�Q5	��\���Y	7��wc�̧���6��\����~�;mʅu�GdN!r
��*�����e��ja�;�Κ9�*�"�f{
��L�OC�|����g��w�|sؽW̕�%�f�hz3�o�f�"��Ҋ��:Q�H�Xr)�E�X>�$��S�!��u��T0aP#��t?��v5���3a�a`�K�UD�_�hs��5���H
��,�ۇD!���y<=�g�~9�.�ۛ��E���' �Ն3g2�v2�>�Ʒ7��N���Ե��ޕ+�G�
���M7e5���Mj.?mZ4Ľw�@�x�D�ikp #��tB�$�g��V��^��
�r����[��Q/^���I���������Q
�x���P<���STMoVә݁��~����D3;M	>���:� D]a=G��L�&����o�r���`~<K���-�|7Hc�L,�W�k�`�#
���A�M��qmp����o`�������8�)>\r�mގ�BZ�����������-G��*2����>�t�����0���r.�!���kÞ��{�v�>��V�t��We@�B�T�F]�D�֩�W���7�bO����+p}���5�����2�(X�~�"�Џ�n����S�u��Wf���=��7��}�3�Z�U��)D�X�%����M�xuc}�? ��o��>�qp:y���)�JYZ".�j�X�~0�μb�ӹ0Av<�6Xc�S<9�V��בD=��P8}ʨ{��z���c�r%��2��f{F��Q ��Ϻ�ؘ�O���a����1��� ��q[��i��?=�����dx�{�oEy��>�Wۍ��  �D�5zMrb,�'1���!��bb,`T��(��Q��J�}o�m�5�f����f1�lr���{��/?vYk��{�Sښp��Ǡ[W��ѯ��աP�H$��=PC���\`!�t�2�b̩G��6�+_��uM�z퉨��z�ch�I4�X��-z�ի���sg��e�������b��f�Y�q����n}7�ѬőN7�[}5�LNf���d���٘�����3zcƓ�1��9��H�����8�'&�p�;��"�}���w���,��s���و�yD��lT�
 Huv
A�qw$m��{(dp��mb�)�V+J���9l���g&�܁����RVo�ō��"]KS`����pbpCj�h0ۖ��~�ukC\pǟ���Ǟ�\}����u���"�t���ڽ�\8�	�>�U$�	���������c�1�� �M�vܾ��Y�_>�M���>�L��� ᷼��2�2��ѳ��Z�i�/�-¡������'~�W��k�
خ:����%���X�`Z�w�Ǳ���}/���]�Љ�s����Of����������|�5�/�L;�j�����`�7i���f�8D�)�k7��+�}�1*bs�Vj>%ĢP��#S��'	XKo��afM���ч�{�ɟ�_�^�#h߷��A���CJqF1�Je��(�Zгk0ᢃ�ry�_�0m����G�\����S��bA��w$v����N39�j��f7`�I����ѵ�Ud}`}+�����ݹ˰^�AU2�[���p�	?�N;*��������}
�]�~;����{	���mo����c�	;�Gf�/��G�����L�:��ޛ�O��v��S͆�p�ч��ú�*4n ���	��fu7�;ءg~}t?<��\|�,#�	a9/�	�.�궫�}#\A�`���B�sS�E[�& �H���JIP�m���`l�v߸M�z��^��-%
$j-�R~{#�����:#W���,�N99�M^s��$�V~��c�S�(����Ba�n9�B!��]%����L��B��j�Վ�ֶFxe6+� ��Ч_����-L�d��e8��ݽ+��V��oB}C'�c	��[��Z�e�䠐P��A�J�V�mCn�h�&���_��J����:\e��",听�C{فG�	�w,Q PmG��E���A��p��X"H��E#z�J ҜiT���d���ɷ�:��ߝ��wf���mM��H��ٔ�*�3E��@�z/�4�vL�ep#�74��H�P�\�^��"րnZ(�J�c����h!�%O����8�b	�W���V�%�h��ajUx�e�ښb���2m>���t3&���Dܹҏ���X�d;��x9�c&JtR��(����F�YJK�P�G:��lG��!���x�$�fR�|�ݲ���	��	����Qj�p����'��L-E�dmR�$U�n��1���1&�ҁ���>���9�����y�d��$-�N�+'acȴt��dWA�-�mn����
3���G6�!�Ƅ��#l(�uUӰ'ס�x��v�|*|�Y�ܶQ�J�S�6�@��]O�4x��\�\l���<�I�7��䁍�z�dP`K��""�<Kn<�<bF�ؒ���U:���(�]L��T*�#�E�"�� �]S^�	�� �u<(� 33e�Q*�?C�1Q�d[M�s���!�������7�CH~��e"��7آ	-����W�oƶI�-��!��u��x>�)�f����6TgMԷ�	9I�o���p=f� It���/�1��K�G�[3\yR��!�nh0��O~��9��Z䒭X,J��m0����.�E�%�տ����!,g�f��R�@��-@gG�qHt���'�uHPY'��Qd�P���E�;���|^f�cJj%�M��tb��N�,��QN�^�ȖCՂF�1�kW���c|��h�j�(R���K%��ǶL�t״b(]xAI���'���Ϫ��L�$�.�\oe1Z�IV@Wz�P��u�✘|�i(���h+�$C9�	![y��W��1C�AQX~Y�wT[�ZaHU�DL�e'��t����d�"D@6>Qi$�9���Ǫ7�D2[�Q"��V"�A�U2��䁂��#V����y
�<	�0p��3�U0c�eP	 ��ј�R!/*ER\:@�'˂K{�h+�u������|f&�|ɖk�)�>�_C/������!���	S�±SR"��v)'�1W�c�O&�-����8�����)�D&f_6�B�3����(���#H�g\1�q;�4e4��T !z\�.ȶ��ݾ��:L�$�/R�N�W*"��(�����tH\���ֶP��4D�e��W��u(�T��ĉ%%��R �%��c��]Au�A"��b�E�ku�ĥ
ZK�����\}+�C$j�F�at ;Y�t��/���FC�����nG�ן�~���Q�Z�+��. ��z b��5;���Ү*>�~A�V]?�=IU1�s\d�H�e���e�2���B�g�@	����6����L��;�z�=�tx������.���%[ذu9rm+�Y�����(R=?��J�Z���1��}7�2Pg�%C�l����X��2�f�`��T��mҷ%D�+�E���kuEu׾(���ld��I	�-�L��.A�V؊��M5��{������P0�P�g����ڜ9Њ�Q��,�
ꊆ(�_`�`����m��&��D��bB����R���>\h�*l��P�{ �e�%@Ls��rff��/�EˬH���ƀ(N�DgY�`x����]8=�����Ku�G�9W�e���p��b+��J����1P΋X�D��=����s�bS��?O���@1�������2�����S��/ zFv7`w�@c����z����8��?�4�1�W���G	�s�E�O!Ձ���$Y��I���f�E!�p��Opc���Q(�b�LԘEH%9J��1c|zǿ!cXAU�&|6����cp��=�d��|�vL1�\W���$V�g1v�8�<���?�F���ܷ�P��<�|�ƣ�g�8%�(f9єU|S8�=ޞw��{s�ԋ�q�Y�b]P���!08����8:mh�x���q�Ǡ�*�|�m%S���W��e#!�SO?�O�n�.GCeyƓp핑r$�"��,v����G�+�����{�$z=pᖋ0l���'^�����Q�E�Q��fɑ\��������gb�������
��I���S%-�G#k�����%M�v�c����T�� 4���cף)B�JIԇ-�=����5�*%��h-�u�E�`�Iا�g���b��y��ȼ�I���/�N��A��P�네3�����������1��?�� jw)�(k��m��%�$^�KL��"{��)�,��z��~�~V�}z9M8﷿��0bP��,�T�B�d&�1��'��7-���+����Z��.٤�N/�ӗ�Ð�&��ݱ�9��C�84NwI �4�\WP�0�x�Y��4���9��i>0��5u�$^Z>k^y��]/L�
�U�]���CA���j|2n�n*���.��H����2��C�ƽU��i�!l&#s��K�<ߚ���s}y5޻uι�D�kI��ܒ~ԨL813m�/�!�<�*�=a,�>��Df��������ܗ����0��?������JA554���o�|�<��d:������mH����t
۰���7��O��� �BG��XX��bP���G���K��㗗b}P'��m��˷�������0(���c����������%'�(=�׏���=�qH$�N��P4ѫ�����������a�%�����A��(��TU>�|>n��A�7�����#ű)]�(橮$��-iW?�cx��ؕlm`P���	W��O�A�v�
[�8�}��b��n��n�N=�bl�a���@ul��ٝ��r3
_��E3�Ľ���sr�^!�G�w��C�������ć^��LC#:��'�&�Ð�7�?V̺=�\z�)(�R�G�l��lT��-<��ۘ��~z�zW�%�a(PL��b�[�`P|.<�h��,J�{��x(�B�(�D�������c���E:H�d�����!j�,r�����'�����Y٥2�i$( k)�Y5�v��.ĵ�c�K�Z�f��y��F�
�CK2�nz��Ç.���}+F��U�o0{�8�̟���n�R��J0d�� _,�w#��N'�n�]���/���o=����.����U`�&&
ӌ�+���G�c�3��Yw�I�8�F2։K`�Κ�[�Əu�O9^�����nR�������k�t�p	��C��rXF������=�]��8�!Α��L�GG��G���'I\z����W%��Yh�(0�Y�	nM�An��X��$<0c<�0#T���^�v��̆i��}�?����h:�esVS��9ͷ�C7<t���;:[#���训�[�/A�6zVs���8��#��T�$�d\�m��9+����a��[�&8̒�@�'�d��g�c�돠W�ZQ���O����a���L�T��M�7�1�tkD��*�0c4|���h��%���E�n�-�uM����$%��A����v'��Xl(שVT�(߅��]w1���W����@)��g9P�!+.�Xt]l4�6]    IDATZ�G���=�d������	�*0���#��N��$!8w�]" 0��eőI�֬�2����"�r�g¢=�f��Q��#2�n�|�@���N�2��倷��ӈ8GC9"���'���7ջ��(������>���� �44��$c0�G�Mōl��z�����J�1����)��7�OF�{��K�
�*oL�����
)��j���������(��B�́[���/_�抗p����e�2��t�n�$�NSs
�W�ÂFk��߯G"�Q���-�d`�m������Nئ��BlM 5�RZ=p�$�����Y�A܇l� �=�Jl. %��g?W*r���#2Sƍ�2�ok�:�RcL��Y
������P�{u�D�^�\@��2u���y��w�ᱏW*;�$qL�����}/B�d5�$���u]��P�6,}{Z?z��6(�]`(�;Ճ7�1���h��Q�Ff���Z�c�;c'�K��!�٪(d���1[pc�����o���6�S.C[�V�y`�-�-x������
Ze�*�@^�� =��ɮ��kZp�3��ЩhM��zEށ�HW<X�>[S�B2��!c�K�A�o��Eӊ�� �E�/���t=n4�|�|5�C]�@mЪ2�_���xE�>c�I`�.�V/����tc`p���uT��X��T9JPhS�+Jn3d�o��p�a�?���Z�h�Dƽ���Z�a��b��|�8��\��v��.r#�IUk�������C�þ�C�슂�XJ,�J�+X��x��?�����f�!��F�k�1|�]x��T��pK�:�)_)V7k�.�:̾��ck����G�Qbjō�sN$%}tbYj/O�	�l��$1� �Wc���W��lW[T����Ӓ1����(ql��0m�?̞�k�#hһ�d�Na�Д��1mt�rX��$���� �m�K=u7A�T`��AWs�C���c$0Ȱ־؆%c�k:�H��'$AL.-�?�dZ��+K�/{<����U���E8p�uh��Q�و⁰]�`nn�_��������7�U3g
�W�0�V.o���ߏ�gޏb��pEԅŪjUU��L����%Ό��_�Y�������F��hYf��c_�b�fg���eH�t |���\�X��3��KX����%RXE��'��(�U���$�%�e��֎%o݃���_6Z�o)c��<J��NR'>Da�:������-6�O={)ӤӵHʜg�{�rM��xa�R<��2|�x�h�ȋ|�rT��@������Ϸ������\ps?�M�!V�FkW�1�ҩt�d�v 9z"��Y�$,����l�J:[C8����������|�΃�=�.<� 	���M�h���!�!����K��c+qȹ�Ь�6v[��6�翈�/܊�R���U���I��r ���&��L��
C�ƣZ�ہQ)>�gq��}��{�}\\��#z*0��c�o�c�D'���*��V�]���7���'W�a�eW�)c2ǨC�
��o�\�����G�dZk$$0�����}�Ԯp�}*cc`�(��O�1�&|8�5����'��Y`l�^!v��o��Q�Q}��c�;ӱK�s?y�L.��SGh%0���3�%0z���=�Dʄ�oC2F�(QNӢ�-���}����r~�!d�v���^�"5A��*��%�����*cl)0��І%o�������of=�]b���S��S��.���&Vn���-#�g�X���^�μ�F�ZLىs���$;�%,z�VL����ƈ�π�-�-����vu#.���{xc`���f<�X\	.�v�0|[`�;���E�?��x��r�hp���ܩ������Ģj�x�k<�\#�=��#�(Q`]���7����W�A�ƨ����/��ƚ��(r�ChO@��*���/+̐�f�(08����qS���?[|n���]"-�h�!����(����ͬ�%1眰?b�n�$ ���R���T��*O����ԂCϾ{��0�!���ƌq����I`DXN����5\|�r�	�"��� �U����c����jծ�WG��q�TsW���x�Q�nǏA͎Rn]�Ս6!d%����G��g����sc�*����yMܮFʽ�I4�����7�`���C���f��l\.�L8 �0w>�~9�A'AZ�vՐ�j�YƂ����g�boh��"x��U5�㢫H�.k�x���x��=�FlM��Kl�.]I-T`,~~n��<���;�!s	�j�F����hn*���f [����*��H��H�[�0�%wt0clu`���u˥���׮��
�D�@i���Φ
�@����	c�;��D��Q&G�z�Da���������̀p8�D���� �L����P���^8`��X��;aœ�������q�0�E����J5��X*:)�X(�}�tv��H�]a�`�� +�8u�,���ͺ(m��nQ�{8	"A��ϙ[9Qt=��8=!:�$o3؜@C����YX����(T f��m:x=��*��C�`uƐKF��[��U����&�Lc����P���1<�!���|�yԖV��)�����Ñ��Ќ�4�0D�����}�DJ1�`�̳Ǣ��Q��"<V�q��d>���.���OM��i7�*ge�,�]�����cq���LL������bu��0�sՈ�4b�<"�6`��5}�+Ǝ���%]�D%���2�MA4���<�����Ϯ�t�d�Ő/;���JҘ���(��Pn�n[���^@X���iZ�(�C�z'`�ð���G:��lR�}�cA�xi���c���&�8�%J|��.Ǽ�1X�eW$,�FW�>�N�]	Q�X_P,(����C����FW����/��'���iׇ�,S����1�D!���:�3�^��'\���{��ɹ,&wT�R�x+��WON���7���&Q�m|�Es������[31m�+8l��X�s���+�	��t�f��wr�?��7ހ�����7��6��$P٘��s�˜����[�5�����<�q�bէ/!\�
���2.��8
W[e��{ �F��W?���b�翇"���)nw	��׌`�{�������"�N����^�!���������и�<���06X=�JMXW�*2��i���d�E��[�]%����s-~w���>��0�O�N�-Sp��G^	?DU���`�IW��;�:���g���!��ފ���wb��7
�U��h2P	7��ƛo���z��=��t����Y6���d:�����B��R����:�nM�|Y��1L�Y��4��^��F�b�������ki4��+�_<�i׏j �°�
�Vf@9ЌLC�$�>�&^��{��9(�c�-M��@��_��z�VL��F$��rW"Z>r"I�$�S@��͝����C.{��9��_!��5�%�a�n(.���YcL��#r�[�J�x��
sf܌���$O'1���Җ��%��ō 邇sG^��']��n0�<i�-�Z�Q����]�}�nL�~���hW�5*�c���)+���x=��>���]ap�	��j��Q�7���h]��p�h$l�|^p����@��`Oa"``<�>X����^�f�q�\� �]#��x���9o�<�\{�Ŝ�tX1d�98���� �g������
{��TC�E�s%�"��E�1wL�Ն+�!&��`��D}J+-`���q��ǰ��I�$���hZ�0�Wծ�����gv�͗oY�sk�:�NF>��z��ȁ8���D�F7
��ȵ-�����$�<�Jl�eH���+��LS.\��
2(�x�w30�c��K��z��2�$*q�iZxc�'x�Y8�;�����?d��P����P���/x7����F�����`ծ�M�l���䳘��Z�s��h	����h��^��z��(~����r�6�P"�1���J98Ҷ�¾��ԛxc���q6�<e+!�L�N��O�[��>:�M�*��R�n�w����Z���/>����u�DdR��Xr�P�&�3c`H�U��]I4��Q�52��׺M��;��z�B�{��r�>��
�F�1�k��/F����(��7����OF;r+>��Oލߏ�f9#P>���� 
1z=��{}�'��9�;���e��� �8t��zvγhZ�.��L� �`(-�1p�LN�3�^���Vf1��ñ���G$��47���_�	w�L\s���͍�M��x2&�~>��GJ#q'	����xk~��rZ�*xvJ�	nbƬ
3pW���L���nAJ��&��h\��|���O>��w=�C/���ZvJ
Ve[�D�,,�EeC��H|�ٻƏ�ѹg������?P�ٚ� ��m�g�4/�P��\�7��*��h�����w�����"����5��kHy�W~��OL�,@9A�0�s�����
�ͦt�{�~9�5ZY���PS�;�e�9����y�)�
�z\�i*쳍>W��ό������3�E�������O��Âw_D~�Ӏ������Y#�+�wJ>k�w���Yhu�(�D��`��D�5_�GJ,>�AQ�d�.�]�l�M�����7!��A�>?$mG���䐋-�V���W�(��_�PfI1�*1']5"�Q �ݪ�!w�SP�����p�6X�Cw�$C+�JǮD�v��m��I&�Id�:x�S#=O�O��LCa���3(�����Př:��� $7��L:-w�'��������H��ڡ��dh&��� �K�X�{ ���q� cA�A��,�X��6Ӣ��+߈r�(礫���RS���&
�r��%��V�u������T8��3�>F�Av%�]ݚ�PMlK��s\�E�vQq��"G4?�c��Z93%�����dh�	�D:�t!��%�>DBHɂ��Z
�h,�(g����F�r�f4Zbmn�'{J\��4	�ȅ��
�h9+%�9&��X�j�S�G�\D�C�D�R�VY��5���j�*�[�(MPC�5��,^U1�4�*���G�Q��5=JF��O��K���HoDv����F����N�����KYT)Zn��ۡ��QZ���O��dq�)T�@���``�W�GR�\`ZaF�!'KD2�7�!��vI�óU<\I�*?4:-Ẁ%EYC��5��*Spefǉ!� �d
�� s��nW���Vv&JF��7C��L��>8�si���wM�2�4آ����
��+�X4VG&�Id�DEHyK��B_�B�b�A�N�&|<���qc�lή�a�8N��LJ�GE֖�O8J∁$fp*�q��񆋰�����	�;(F�h����E�1A?�5��Qe&U�(?CYw30x+6mJ���r+��H9Ϡ���d��qE��d@�x�"'�x�����H�Ӕh
	?�A�h�G?V>,q���SX�>W0��uTΚ�<�"j���=l�"J1�;"Pi��cgS`��K��e�q�O�9�w����羇r��^�p���E���+�n��7F��se,���QN�܍��<�B�r� ଟ�H\�g��cD�YX���� �y3U`��T�/t��&�b�RA+�e�j����<���Zo���yLX�|<.D[e�d�<�|���`�̈M�q�������J�F�|VTT�#Z���f��k,�~����U�%�kb���_��F�0�Y�D�v'�:Jd���?0$��jW���RW��M�'ʶ|���QGwm'���L))FUᤊS>J�J�C9�#�J��O�T]��U}Q+N��h��Ŧ��V���C*GG�1(���a�5��H��V��,<�� r��p�$yE�"_�~��<�f/Z�c_�1R	�cS��UQ-���QD}~n����/T楊�P��7�j5_��m�*>͍��%0�]��0o�|*K�
kL.Nt!7��Q�D\L�F��H-��,�<~ʏ����0��i���>E�x��,R�Qe����Ճ�o��0��]P*�D��v�v�8:�虁�T&=<�:\I&(}�YI%}Nf
�xx|H���[&��F+1:�YC*�Q�I�-�3k ��{��M���T���Mq7EƔ��*G�a�{D�I�ԋ�Ht�5�>�L��2~�k�i�fy���_���$z� Fda%$ y��gy�� WD@9R"־ �&�|�����B.x�RE���UlO�K��At�J9e>i��������.���{�*y�6�n\Ή�w���@��ZW܊����}��V�P}$�I^f&Փ�5��B6�Fbv$�������fS�j,�U sr��ḷ@�����"e�����ˢS�g�L�U�*���Z�!hפ���x�'���o"�m�#	��ƿ���N�W7����sjE�&�6�+ ��_Ԏ�8�����eJ��w!�	Ӷ�泈9Ԩ����F����rY%���!G��g.<7�H>�eU��p�u���:M��d�Q����S�CPwӎǐ)����e����ԓĖ��\����J�@��N"��Fw�جZc��0�(����%�^�Ϩے���Q�]�Q�ߩ ��3T'�^�����p��ZLJ�D�+����~��ˎ� Gn���:z	E������)�;��<0�4"����e�w��=�PB])�����/�p�У�gY	����ؘ+�q��P#E'���E*���2��)����Z?�[1�G�"�T��ȕJ(���;�QA���$� vٓ��O���,��*�b�Y������ి�WZ�ddN���rQ���ř��9Q��/X�Yp��y��ٕZf������k�����W
08�|)�):P<�|T�.�&l~��e,����}�y�:t�ɟw c�$�I���r��(zE��h��PcI��>)�Y ��E8�����l�[�s#6��b>+j8��EN�"pRhn/"��H�yT[�ީ�Y�n�RI�VR���� ��D�4��"h]���!i���e_d�S19��t�o%�C=z��rU�0Ljp� �����D|U�ln� �K�А��r������m�U��j������P����t+F�(q�e��P��ކOo?==����)�30�L�q�ЋT`�G��,ʬ���վeb������m�ߦ~����5��D��jt�H��֮Z�uO�n������) Ā ��/��^�\��;��mR3p�W���� ����ߧ�~���g����? ^���m	��~:����g'���=��hhk�@=�a���3b�Ӊ��bI����{�V�dQ(f�b�����؄��
�$ߑ?W6V;���S>����IU��to|�2 �!t�<ЬYX�q�������a�n�h�s�8��-�ŷ���wJ`���<�̟�}��?�;�E\s�0�n�I4���E�[����?c82f-��.C�����᧣*��!�=����m����Ћ�AZ�F,,�����нk�,�x\P��ؒ�0��I���@�'bz�O']�a瞈���F�Ǜ@�=��6�K�n�Cp�1Hl��}GIOS����X�(ss�|ci�r�Hؾ���~�Ѯ���Yx�F^ ��TZ�ʤwk����r:.��P󞲡8V&*�]TQ�4\ɦ�N}ae�0kҘ�)��w��n!0=r���7F,Z�t���q|�.~M�&c�u� ȳk�P`�Ӱ��9��F_�Ç_�l�;��E�;�q��Q*)�5�I���_���u9\5�&0�jd���i|t�Y���PW�I::'��J���>���$h�,���]�\w�Ht��M�b�]�_b��%�c�� �Ͼ�Z5���^JY�F��m����o<�`��$������b.�,�D��ǯ�АB3*Z��T��D���Qc\v-���<�Ja��F��^����)�H _n    IDAT��r`L��5���>A2�Fw*��qѡ4�,¦�X��͘���ÆǳMv:V�p��q8�?�9�-K���`�b2�v�w�"eؖ�ōy���Sq��k��o@����[~��:]z�Tn��}�]Ӏߎ��G��t��Pk����q���SC� di�(]�����.����D�Aڬ���E~ ��5���%T�!�~�6r+���N{��������R�t)�#E���������V�r!Tn��a5_2�ć@=M�\u�����-���F����愑�S�{�g�����.�7md��Hī��K��c���q����2� N��� vqc��D2�hKl��_�p��I��9���N,��0e�p�Tr�MXo�@�܌�������.]�t3��Db�,�4g��=~<���V����N�M�G�.�jmz�5�� ��8{�x:�7(��mV'��!�r¶��J
��KRp�9|3�֭��CQ"�?g7#�P����;	�������h��uߴ�Wˍ��7����۰��u(��%> l�"��D��a��/��g��]�O?f���>i�w%��y���G]��!�!��'5�$P�*���UBn�L�|�6<x��02=A���t��l��އ�-�Ѽ�+�߹��*O)�8+U�|����a�~�$6��	��[���ᦫ���[7�+(�H��bX1\x���w��ж��b��y6n�r(���	ߧ1�����A1���+nĮ�ׯ���j�2�L8�kg"�5U(b�ϡв;>.�n���Y�W��+���X<���+�Ҏ�,�Xl��L��r���"�Y�f��?F�b�YW2l����n���-v%*0���!N�zԉ���q]"A��0���oc��ɸ��+��-]�h�h)��e�q��p���b�����c�_oÌG���#�K%MGm"�EkҸ��;p�W�X�z~>��t�t݅���C2'��o���bI�2l�����:��bָ���G��s��� ��I�z�F\�}~zܮ��uF.�e6!$��إ5�c��O!�Ҍ��OKD��h�(��j�*���\���d
���o���h��� Q�r����2w&�\�O+�O�Ƞ}��h��)�I��w�<�}��1z���.>�}��]��z�A$��q�H�W��Ϟ�.*2J���N�c<�i�c�U7��F���B�j)>Ǐ��,Kj�`�r	�(����f�q�yi�q����O#ѩKW��p���i� �sɕr��ﳏ�-�<�R�r�p��7.#���������O|�Q0z�\�rNg���'��U�6�a��#�܂���	\����Z�݋�W�[�"��ʪ��q+�cK��nį�*"�c�U�SE��V8�72Ȭ���9�c��k7|�?���I���rƘ��މFԋ�,�Ǧ�"�r�x��JM�.��#��[P�P,p���C[��ܯ��?%��r�V|��A�vqF��[HB|��$v�y$7�(|��k�uie���+kh��;}���;�K������y��CUu��Q�.�:C<��y�=���Z]_R�������wV��'̰��ȥS]����E�����%�F��j,�\"��R�������޶�����T�&E�BU�wZ��d`�H��ȭ~k�|�A�ƉM��m��Ʊ�w�	�;�1�~75r:�|������ yq�!��2c�+^X��S� ��a`O��� ����^�h@f���*rT�*�����������Wym��y�op����g��9�Y��O��M:��[�Z���E�^��lK�r
z�,��U�R䏋�����Q��i��ŕt���
�韼8W�Qo@$u����|���H�iV����nD���ĳ�&�u���{�{��3G���>L�F���y|���(~�*Pj�11��!��Ӱi_�`#��T���-�~$��L8�ݨ�Z�ԱPR���M�'��'�X��^v���d_��~������y2�R�sz��w<���*4y5HF�'ї�3c00x����g(j��J`Tgj$��Ѱٗo�P��e��E����^S�6z�S0����QQ��MT�mȯ~Ec�97#n���1��1e�#�9���O��A��ڰ+ߞ�?[U,Tn�T=j��p��1Me�
Eo�����4��=A��Wc��z�	eSs$�V,�D�5V󏲌���B�ΫG�lu�������5?G�
:g��n:��Gl
��<���D_G}؎��@������V�By?ɵvEZR�6��Q[l�eC�yM�Q;r�ȕ�����A2�����&�FJ�^Ɗ/?��a��1C̾�ܶ;o}����E�����!QX���ߏ5��EP���iM��$�@��ʲ�B*7K	H�/b�*�XL���h���h-�D�1sk+.F�d�O�	������E�1�����U�4A����@��� �_�ɒ��A�09J*�d����5��ϐ�E5�ڕT��Y9"3G*Ҳ��M7D��:rR�����_�
C��b�QGö��$r<ʨF��D�I7=���hcq��j��ȶ���ӑ�[P\�*V~�)vv�pwgO�6��Qm�]�z�?;����s�9J�%袷c��w������J�<*�Y�������Xe���:z��#�n��Q2Q��+�o}��n�6
�Ejn������=O�f��@����y�}������������<
%t��a�p���"7�j|^q�L	��M�TA��(�@(��O�Q,{����d09�Y�T�������!(;ΐ+�2}1���.j�k�Q*����]Wl?.�X+;J�Q�GU��.i�"��-���s�~�8�u�(�)�F��vu�O�쬋�v�᷋!
U��X��d4}� _Ā~c���&����6\Q`D ���S�CJUc�������lt�AfxCd���lW��d�=���D w�C��r�(�[ø@�C%�O{��Eo܄���hZ�ɺ8R5�ZĬ�̅ׯ@�ϡK���)heq-@�m��M�Wա�~�~��W."nSۣ���Ĝ�VJ���!�������wb�"a�!��]	��î��������#�=�-0: ZDj&���.��$� LG��Am*���q�b�N]�u�V!$.��G6ׂ�_D�>}Pv������epةK7؉*�3��H!�H+�ǆ�b'KvB5�g��e̱���H`�}�Ň�s�o���Q��|[`t<c���bNc�%e�+-&Qd6t��$@�Z��������%�;%�HQ�\C�i���	͙ft���U-{�L����X5R��a�q�n ǈڬض��ص=`�ꐰ���,il��2ƶ����EdbQ�J,#0���D��Cw������"��:��>GU�ӱ�f�R�.Q�9��T�����k_J<��g�y�X��ֵrĕ2^�K<U��E�L9'lE`�O�e�!g�~ʗ�2��Vc��͔9��3�	����ۑ͵�h�[�ż7���K�h\���z����~{b�;!,瑬������,�[odJ@]�t0�^��b��ڶe�'�5�K�2�$ I[� � ]�t���X`L���qC/���m5FGj��<�E�̒#@!�Ќ\a�����n@��yX7�E��i��ð��H8:���!t��HR RH��X�f-&M��Oޞ�Ԡ�ѵ��j5XղN�
U��H�k�20ȋX����-0Tq�q��NWB7���(#�s��mhA3��%�
��ڴޒ/D���}1��Y��t�2��k�����r��q7�/~Hv�vA��.Ы�Qݝ;���Ȓs
>�f%�q����e�m�gǋO.����Lő˷�n��Bz����n��/�Ev���i���'�
z�ҥO?���Ԇ6<�G2a�-�ʮ��;'ބ��yI��v�%�k֖�������+Jb�ǀ�ʐ�FB��hJH��]|n��{��� ���|#�$��!��)�cݢYh�`�;dw|��,����pvۡ�?�ڮp�	����T�
�n��?�$vؾR�:|>ov�7�7����a��G�h�@10�1������Q񹱘�B`�5~���uҜm���T|���	
�X�~B��TM
u5lw=�~�~@[#׎�{�C*Y��m/u,Y�5vݥ?�|��;�X,�;n��=�,RH�-��yTW�b��ň�vG[����T�G��i}�X-��pI�)nޕ(��p�o��]��G�F��j�ge^�Ѻ�t�3�塃1�曰]����j`��siT�m̝?��&M��rp�mwcƣO���3�V�/+ee��_�#~zjz����?�����������I`P��(|%I��%0��ķ��ಋ�������V��^�����57��Q��in��ӧ��v���HC�|�,�f.~pȁ�a���6�A���V<7���\Ĭ �����W�m(���OD��' ^������D���@qy�T���1��Vo��X�+=�G"��^3kg?���<�r	5	wO������N�z������KX��B���ؿ� �KG�/�tt,\����wO��{�~�����p��GB�h"@Ae��E������Ə>d�5ƶ��x`��:a��Cqo=V}�:���b��W��n��X2Ҿs��x��ѣWOh�rՏ��4��B/�Ìk�X�p!v8wO�S���୆�_zS&>��G�����^#��[�%���m��q����U2��p�lW��liٴ]�pj�N�
��2Bz�S���Q��aeW`��᷿����XP��a� ��q�ģ�>���	a����!�l���F�f�B��q�u�4�$R(�6(�����e0�������Ъu������U'W�1�*�@b;h ��G����[F�ő�^�Px���j-��x��G"��.>�z^��L[+�f�&���r��FM����^���g��]+�懯�	R��*�m���ǟG���#��R��8�X�r%z����M'\����Q*�D�xyc�=�|�8�8��;�A,=�T���j�AJ�	P�N����0=jpu,0�L{�ء����H��fx��<�Za/DÇW.��ϡ�����FQhCJˢ�q��S��:)GC>O��j�	�x��'0a���ڥ'�H ���͵��@{.��+W��_��]�r��N�8�l3庐�}�I{8���Q��1�[���U�db�*h�B�3�-*G�1�߄��,����,0HhA�=~��Q����S��tX����CY��y�V$�~�N8nW;�(���P%aHc���3q��Qߩ�D|�t�@L)_D"V/��_-���O�F�w�L;H.��6Z�"�l����n�8�0�Bہ%��}�H��|Z��f0����m��OP���y-?��~��D�n��$v�bl���X>���]�{o���&��ke��ʛ���?^�xʑ����#�+#��(��T��r��`���8�����s��%?@��{�K�>�8����5B�jS���QW���1���a�؏'�߱��=�=v̙#�=��(Q��{�Rr�)W�����ĳ*$�:(�tۑ^�!�~����}��-$�$f�������Zt�^��rG�������跣�a�FOk�҅M8o�i8��(��$F\5�8�~����6<�23���ZEE``���u�l�`>�;c�8�h�P�\�IA`�!R�
}]
t8�!SJ����k��_��d�r9�{W|��,\~����E}������NҶc�U��k���w�{��B���I�
� �+�b����8���p��g`]&��:����{�r,�2�vĲd,`�HuY�%��m��]��� ��A�;Օ�S`N�V\��22�Pη�q]��6-��~�4���#q���ѥ�u��#T%Y5�<�����ѩ7.9
󾚋;@�/H+L%�l:�5+��1c��1�'~]�9�H%��RH:5���h�
泂���w	�=*>�e��g�
J��t%�(a`�e��u6�'i�C�
i���
��кA)��d'����2������Q@���I��!��a��F�iL{�>���&��=࢑���/�`��v�C�PSǒ���u�n?<Zjg�M�����������V�0�-��7^|���S�}��]��N��9}�Y�2���n��V�;�'X�Q*`��X��X�L$�<J�s���;�`=�î���Ʀh-��࣏��Gg�b1�Z2�IT�m��W'au�Zlק�N6��Wd��G�.G��.��d�D	1xAA)�TT���d&"
;¹�-0��v�bJFd��� ќ��G`�f�+ۈ;&� �}V�{������4����+��@�����|Q�3J���I����,D�.�L{�k�d/��o�E�a��M��(+oڍ\0����C�S.����Y�F��\!)�%EAS�#�+m�����(���ˮ�QhDz�B俞+,> �g܃~�C!�G�U�l[;�S4��3����1삑X�p`uj��ǀ��%�h�+��U���f�N�� �[�wQ�����dE8j�P���Z�m!0�T,v�k_�Ppې).B�!Z�Y[�̪�X�����y眂�T́S�P.`;:��툧��vsXٴ�~_�nB�� x8�2y��6���n��B���6�]��١��������1Ó��2n��u*�l�9�SB*GG�U|n�+��E�L�$	�U�as�ihI�E[q9KC�n;A+���䱦1�� \C^�0{����llhX�҂�\y�qe���>���]Q�Q�Kؐ��"i��.]�"�̒XT(�f����&��VsW+�Q�v<0�+��+��E[��h:ׂl�
;�e��)Z�#,� �~|/-���6�X�0ӪtA�����F�^�D����Э��ր����iȕ��PLCגH�I��d��|^��
G��#c���Z����
�o���f�^�����@;j{ht.2�۾ȱ�c¥�L�J��mH��D��Z��8VI<泅"z��߷�[6
���7ÉU!����T���D6���DcLi&�"_-v'�B`�9�#RKӨ|�K���۽=b�+�v�7�9���T���*�"U���
�S��x"���FÅM�����~j��6�AP2���O�B�?yM�v?�Z�Aw �MP���3��110Zڰ�?�*�Q)�"��)4/5�Q)�b#�klx����;���v�hȣ{��0�N(�<z���s}t��Kp§VƲ��E��o��Q(�g�$Cp�B������9�)�U_���}�U��\}��8tQ)bP{ID��D����E# �t�b/4iV�I�����X��Ac56l�H?e�U_�����A�9ƛ���Խ�����o�D*4�����pp��;>[�s���ɬd��=�|��aL������Z'�F
��gغ�Q|��@�$p��t@�Z������lJ{�$�o�`P�l��P�l��'�B/:&��2-2��kCiᣳD[AFGb��o9`E��=����M]T��),��;u���g_���>�=EjbP���o��j-�w��0�[r�9�L�Q],#J��-����!����4GQ ���b	��B�RSW+�B8g�l�Z��ܹ3L3%FB�%~��i�02)�LR(%�wa۴ќ/���R2��:\TY6�n1��(}��%���kW�8�8���o�Ըtᴣ�H2���>y��e؈��2�I���O���~�[Q�4O��	q�h�)�+ތ�C�,������$�P�QsT�D$�P\\�pMPuȐV���S�9�����C5/�s�-�'R9��I��0ۨ553v3bR뛰z�cF,�{��vJ�7�XDb%������5���u"�I3T�E-ơ�_q�B٘���Js�ZE����AnڼA���:����P��#�!)�lK�hD
���ɩ�}!Zr    IDATj"��ޅak(� ���ס�<�v����F�c/!����7p��kP�ұr�؆�g�G�ye�<|�2��4B=�<������'� ��,4r���ي�Fi�JH��b��%>Q�{�LD��\C{��Nhs��n��NQ��X�r�[��1�\V�%���ka�E�b�'�iH�%��d9�>Ǎ^�sRB.���dV�#4��x�韢����	��nC�bT����Cc;�,�:c2�XS+!0QR��c���Ii�567H~��f�/"b���J�4j�E}�!2T����F�q��Q	A�sX�z��'��ٹ�lh��Z��nM?�yZ�?�������n���x����\0���#.|��y�`�d~��76i�1<T?ŧ�����X��3�C�V\,�Z�J�J֜�[�3W`Ř{� H�UIO*��Q�$HH��,A�����4ũe���:�*�'�YʑV���,v�s���p�5ȥ�F�q�/�7��I�T�7�ݧI�ք�π���0���Ȕ�"� �7�2!������	�u�X�3YqJl��V����6��L���s���Qc��7�q�K�2�48�V�4n��:���S�d�l}g4�}	��~�.�]:����?jX>��^z����{9�ҩ~;x�
1.�v�6c��?��g)Z�L�l;����u"���w����X��I�.Z,L�b�Bj�^��d&I�`�F�4a����Z����\1���Dah�G����D�����%�6�>�c��3М��J��[�y��4s�&��_�Za�%D��8��r�bK��bPI�Ee�C]���X�'?�&�y?�kN8@���0	��g��(|�7����'����"�����~=�{`%:����7�v�[8�2
5c�	�o��g�P<��M�بu����h�[x���h��v���J?���PY�#q	��Ɯ�%E�J�j�>:�.�.c/@"!�R��"��1�o�y�B�R��\/'�=���>�y���͘N�3����<�*lF���N���n�ZcU�2�A߃�*��GEf�al�S��]�*�`1A�B�)wV��$���/f࣠�R<j�J�ÒԆ�S��N���b��	�ϛ��	Җ
U|[�m��`������q��}kW����@mFów�m�a,}������Ѝ2RQ��#���PD�[? 6��C���,d�<����%��5��kV�԰��.�?��E�+�NW�X,�6-4=|��&T�7�ȁN��G�c�^]PW�UR��:	]�g�a�+o �Wo�U]�IYBF������Z%�#�Ym����kk��� ��л�~'��f���	�p8 υ�j���EMW��|T�5_��";�:�ݫ�nb���@�$��*���B���$��T�(8� �9���C�ք�����3�ǡ�:I��n��,�nC���}�p��*�}�uq�lT�����x֞=Ʋ?�FOX���/_&��je�Z	�pa��3"�׿�w���͞�Դ$l%��i��E�dS#���f���S���5����a�U��0(�+�S�j�ç[��>uN�t5�tG�yr�T,Zp�w��iQZ�q]rz�6�N���}6����񻅓1�4�ثtS����*\�pp�sp�)g��r��.؊p���a�O��6��w��
[����S�#�D�DAY����P-V|�(?��
 ��nI>U(�5p�����bOĤ&,�P�0$f4�]e�%+_�߆N�Vl�`%��9�׌������6WF*��>��^_�A��$�}�s\������|��vH>������4��G_~���
^	Y;�XD3D�����_nŃ�_�BQ1�f,�b���m.��q3N�trF-�������Λ-(���g����?ؐ���ޅ�_~���T���E�1o�$t�I#�Pq�D�lW����&_�#�}>r]C�����K0�dt�Tˡ��&�ob��M���N85}��Mn�Q%��|"�闔G0,9���(�K|���1ĵK�h�Q0e���p���H�n�H�͗C�*dZBHk�XT�_W�=t�Aa�:h��H�p��Ǣs]=r�2�ٯP�:�G��g�J|��5�q2v��n۰t�{6��~��.7�_w�FI�D�M3��<�a�5���g���y�����Y[��r�J�̽�;�Z4uȯ���~�hDl�H#)%Ib���ֺm��{pԴ�تף�^ċ7]��7�E����x�#]�@Oa��Y�u�w��_J�X}�E�oҵ[g��s���=�U�Kf-�~������{Ҍ��+��bpfE&q�
���5O��-[��E�D'����+Sb�J�a�e��l]���b|�{�y�'2Vb���f��H ��BQ�yL����	6��'�|ad`�����ա���oF������8h�I�_����ƍ�8��Eبգ�
�vP�-�P�|��>�w�0�Q+ՉC�t���j����믽�\v��m��-�_�1n�5J�V6l�#�"����<���n3mևu�E3^�w���.���$&�R�t���ԫ�����A���Î�xc�EXx�t��M�C]��G"�9��%8�ĳ��<
[�l�c��Z�J}��N�#<�[֭E�#� ��3��Vj��<��	�+��V��Vd�w�w�{�%C���B�t��;�e=�7�c6M�m�nwjPpT�>y���M^$t�/�~y��ym�J����GO���._��Z�f&Fa�=�ϡ�����"}�X�a�)��]T(��[p���PHw�֏V#������	pY:<^)�k60c�8|�4��BU،Wg_��s�a�n�%���d?�UDhW�҉W���磴�I�Z^�sn�=�;�*��I��N-.�6O=ѾG�!L�$�I�Q
)��X� nhH.�a�Q�t-:�_���q��:��FIr�\�l���Y�ɍ�E!��0!���L�72r�U\�-�e�����'� �����+(~�	����v���>��1q�Ͽ>n	���a����&�{mڀ��e|��p��W��K��b��YC�N�'N���hX�.�=s��8yW��-#�P�t�R;e.6k�P�f�2�GX|�4�����R�F=8n��3.�<�>���Kxe�0,�?��v�N�&�އ ]���N<��ǠĘ��(Q3�J�LA�(Sn�LW�����~��ʭ��3ɮ4R�@�XϬu\�C��r��%��]�N��Ft��sa���"%)*�3�JDۃ�?;�,�>��g�dt����m��.nC����'~8z��=�ipI�5�Z*4�4���M|�?����Q*�15���i���<��'8a�Ll�jѼ�cl�ۃ�9f(���S����G���|ڈ{ߏc'^�u��m��6�_�����W���^���0�;������(d5/�5WL��{�iS�̇�a�Rȕ"\y�:��{�-A5"�J4\y���K�xv˚�Z��m�6��P��˔�Th,,ɧ.#�$)��)ZN2"߳��+��
nYVa:*��4��_�(xe2��]jhȗ����ݭ����t|�<�]<v�e��l��۱a����c�;o�h5v'5A�YB�¯���3u�ƈ�(T�5o����/l>`nLшJ��{�V5fp������BԼ	o, h�8���
�2`UZ=z����m�[�_��f.����ZD����W�=c:|�l�PҪ����3t�غ8�Bd�
Bt*7��\4Y�$�F`š$�J4�����.��G� jvg�3�f�r'K��L��<�"�4;+�)n��?�5<RY[��v7����5,]0��=NW���������Ġ	J�^&8�q(��P���?����,� �˴�NJ $,�z
�Z�����Z^�]#5|F/������k��B��b��.e���]�^N~����2uxF
MZ�T-�ЭC嵫�5}��r�8t����G&�$qR03u��Z(�5p� �\�ݨ��ƘGY	X�|BW��=�X�rv(�L&����Z��bq���L
㲶����cIӦăI����a,�n���Jsg5��R�� mZ������%N�a���m�7������?z֥��=>x�]j�J�P)V+ ��z�$��5$Q�y�� ����N6ZaR����
�/!��?�S�%�)Z��$�/�B��n�(�l=]*
��tRI]G�L�͗$�Ϧ�'w{��1E,C,Sig�Q�Z>|*7�z��H�$ϰ�h�[BZg>	P�N�B��������\�<ߚ�;�bi�x��}$������?��vJ������l�ǃ5zv�2��)�ѫ��)��B�h3�q[�1��ѳFL�����!1�x���u�,Q�T:��H���2�ZYk0����"�mnCJ�0*+v|��\��i��Ȯg I$���d��'�?G�ȫ�	��l�0�x
(D�{.��O�0� 6o���J>�˼Df3>0���h���|�L����K��tV�	D4��PG�v�4ĄuM[��wx�7�F	�
��l�K>���x��sQSi6�dh�Y脍b+�_1dԨ����;�Y�c�d�Q�[�j��6����6�%�i2I���>X���y�]J[�P���q:L�Z����BX)n)�n�˓��SKOk���؅GZ-�/c|�|/�&O�f������\ض	�+��<���m�ek�^��h������j���吧�x�>ue��}ʿ4]YT	�21�c���'^��_٭a�}�#g��<���x�3���5�a��C0c�.��.<�n����)W@d�ҭ�}urwuch�,�q�Γ��U�R�N����=Rv_=q�K�X�R�`,'�a��
����t�e��'�g�Zm|@��fg	� =m��c4���z7�C�b��7%���6e��R0p�$��SQX�+r�R˴�|^�x��7_q☑C_ޭa����3FM���6F���-jq����<{VTF�U���&|�H*a~�'�8�e,�[&�q,��-����8F�!-��	W�Q#���"��ƀ��7QCU��)i�/�I�
x�~�s:�*oD�zH���?�c�����<��3�ﬅNT�����P��7[�<hV�
Me�����Z\��E�b����|6/[8�ї���=�#?5e�/�j�"�a�mM��r�FP�4�ӷ�C�k@�cI^ �c�ſ��������?���RS��h�x$�Lx�\ghе3IV�Q�;D�h1&bw`�=�1M=8���֎���o�m��""����@I�3'#��.�� ���vu�c1<��lGr�b� ��ѱ��p�K���!{3�2�7�+	��BI�1b��-[8��=�RQ������d_�Ca�f?����x��@����m�k�3�J�.����s *��{��VW���{�L�N	������x_>V��P֫��G��ʆeo����R񝯖������\8Z�oy����,r0�&�RA�mNUʛ	��cP��=����8�(J%��f5M1�7W���Ο{��R	1�1�'Ti�&��r8b��Cy�����,���*!P�,F�W@my^�c-�=��0�+��R�mj،��M�&O^e���a5�C��5S�'�T�?�\d�U(�K0���،�/���D)�/�����|�7^!�iIN�XLOb���n X{�� �I �A/lDgm+�����=������ҵ��0�/b�[����,�vVD�c����������{$��'ޗ�O�>Co��ϡ0m��C'�u�-�j���0���%m���w[C؆#WV��8�d�E�]dc՝�p���ثc��^� L�����T�|�t���2�F��'(c�c�<b��8z�5�g����!й�A�+&�1��b	l��3)W�򐽗�߈��F<s�L���Km���`��X����`R,�*���롇��F���;>r:�:�ރ�/�OY���%�jh1��;X�%��b���F������=��Q��������0BW��$�e�ni�q�=w"�u�W#h�{7P\>b�T4��Wk�P�� �7�6u���:�z!o�IBC҈S��\5��H|�Y�Ӵ�����0d�	�]���ų0n��8f`/^I��P�X8w>V����D�����a�3X�a�~ElT�qg�!L�@�h^�}\~��i'��0*�mhp�f[ҍ�i���7���5����a��I�֩C�W�E%��KF�P�9�N�����u���p264E�b��8b̵�W퍂Q�*$��\��R�������q��&���M!�`v�C�h3�_2cƟ�c�F�g#O���ebѼ�X��[r�bt����܇|DF�N 5���GLG�����`i���=��%܄�w��0dEqʜ'��1�&�0D��E���T�(,�3];w��^K��p���O��N���=dȉ�B	�����3�.�c���Y�����z�l�1�I�]�<ŗ5A���v�n����DegK(�d7�&�ml����7b�*���T��[��v��y�Gv%����2��l��X��s���1i���dInO���<�J����U���ѹs�j���	�K1BF{^C�R�95e��,��]�|�^(Y�`�Q��	A`�K*1-���~��8W%���zzVP����%31n�98f`_�0�"<±M,�{V�Z�89��'�{�=��c؈��}����,�P2
s���u�s(I<F�c�}}k���h�a��C	�1�4��蓙kT>���Fa�܉�Թ{�����/�a�㹫��x���t��]�u��rfM^��hJ��	�gF�d��c:"����� {Z��C�a�2�����lØ0�,;��pl�*��[�Pr�\�JA[ƞ��#>$a���
�_(�q=�8�������+���y���2rҼ?��0T��鞮sa9�,K)"������F`��ɨ��M<���ɰ)�#GUB	�4�{����O��KGHKPTL>s�O^�c/��l/�*��M�����KbY	��'&�_�0,;�\-;(���9�_<��� ��%M)��0eo���j�W�{��|.��JP��a#����ֆa��v{�6Ɗ�;y���j�a�a�^=�1T��:�1�\��2̝;]:u�K�{��#b�h�+WUɨxs��Æf�'-��/��L/A��&��$S@B$�e�QC��;��v�-ư��w� H�)2�j�~�B��w��/����$��m,�V�z'|U�=��r5f
����/��.إa�Y��QUI�p3V�qyn���C�8D��G�9b�ܧ�b��P���Y$WFd6�mF��1��l:�q:�Lnd���0��F��tT<���Y'�de�7��s�i8��d�@� �|��}L��z�8��ӽШU#G!�te�k�#LH�T�S�J8�a�T6���vu}��q'�9���L&��،��zl�3fa��q��_���EQ9�O�馛��悔ޝR(����~�1�8�7l�5t�$t?�:�z&FW*��8�!��k���RU$��p�%��vø���O9yޟ�j:�N@.��%�!�/n��gxeŵ����9EN�"L8p�Uh�7�?<�1Zݡ�^E�E�
A�AK�n��à��(,���	��&V��o8�G���(�(h\Z,�{5z�$�P���k��P�ʎ��ŋ)#QH+5ZQ�$��8�r#:�#8�6�����e@o�ۧ^PhZ��]�^�����o���JV~�μ&O�����=G �+W(��?��ngM��� ��p]�7$���{�kk�1�m���؉�L�����$� �M�8V��	�x��o��A�l����2'�B(�Co}:c�
�o�M��\����gJ��􀓿-]��⺃	�
ƺj�1QT����I�P#���![�c���H`}
�����l՛aI �Qqh�z�    IDAT���_��@�d�-\�����m~�GT���.D�Yu�Bz[��T[ �:�u��0k���|$�&���0�$�4/_4��=��v���q@�d�+`��}#ȣC*@��`��HBƜ���t��bHJevo�sۊM���Bj��mo���Dx�03Uȗ�l��I�0��I�������A'���+��Z��L����U�CgF���/�1#�V�^!}�+P��x�3�*q�2�
~��c�^��A��Q$a��g	L��6�hv&n��}XE+�Ð�Wo"M�,�f���<�F"x��͟�,�ui�E)��ga!�D���#��,7�\��!�/�LjP�CGI))<]�O!?�0��&1 ������)gU���9�{镴r+���*A�:4M�\�҈i�g�[H�j�c|��j�ؾ��g�,����6?=!#W��Ie�FI<I��\i�q�;k�|��}��F�rAC�)� Nt�Q#Ur,ͤ��y��l��(��%7���![�fkP���?K�6�} �t�pG���2'�݌�܎������??	I�)����"�|aK�Q��G�c;!�8A�DȈ6;�b�x���R�>����+8"��{��q+v����x�$4
�z�X��uJm�6@������0ڄ�jWUR1{Ob�Z�Qw��{&�+�2d�c��I���Q.Tx���(V�� ?R	�Z�yTF�����.�X�����_p����l|4��7�#Ij�O;i�I�T1�ib�\�?5*{�X��%����0	K���(r΂iā��(�[b;3�؃%�n4.A��Z��\v�lE�m0�ۨ0���+�xbl�c(�yk��&�h_�+nq��i��#n)#����f�Ҫ%��!��̡x�=�:�L�S����Gy �V�^*���X̋k%��l�k�ZO��c=*wGMg����Crbe�!�8�I�+�Y�0i�'����sɼDȢ��Ğ�>1lz	~�xO��U��k�O�?!k���%��Da ^)`4y��z��%$w��hLP�x����7Oo�-q��J�t�+Hnl�	�I����O�ѿH-�<�J�8�����[��s���-�S~�1���l9^Ib���mx���-�ɱXFȄQ���v9ȚG쩨%ƽ?R�
���q�{'�xw�bj�4}al��"U����h|��]�֯����cH����ю骂ޫ�͆��bɆ$�'#n�8����$i����\kI�*�H������_�Ժ�3$V�5�0�¸�&�^�k8DV��	h4�c�v%�xr���Q8��p�̟a�+y�R��^J����7Y�ja:n�����!���M����r��GM�G|�$�k���oF{��u�j��Ee�-E� �zc���B0�`�Eۑ}ng�۟���M$y�� �a�?B���a�aҕ���G��� �Cl��&qd퉇��J��1q��i��ai�����~\�R�Dr8Z_�T9�G%{}�o��j �S���{�>Lؾ%�r��x�v ��tQ����j�I=%� C69 |H���sw������#_�8f2]�ױBH�[�Z�&�=.��	��!���7��"Yud���?�*�/���]hh�5�RQ8�T*\1�������D�5)��sԿT�Ί-��Q��ѹ�����i���%� Kj�4��%=^DR��� �Klb:�|���x�<I�J�h�{��H�2C��[��S1h��e�P��k@]M��7�(l�WjĖmM��J�lMg�k:	�g!�����0"�?[]]YH�]=$Uٴb⑊C}�@�Z!�X�������
ٶ}v����[�ў����D�/u3x
�z��E���!���FO�|�r��b-yF[�dL/�=���Q���lpe�r��|Ԛ6�}�W>|���V:=�b���PW��|�lY��"��s �p:����EIKAKנ�(p�>�5�@k�QM҇V}�=>�V_�ŃQ����`_��a���}G���2��˜C@0��|+�B�$S��M0��	>���J�RNO뤬-��g�B�LF#iH��뜩�ѻS5>~�oX� o�N�C�9��?2�(����T��o���<�L�|*`T��w�G�����ed����2wQ��˅�(UM���V���*��dUA	ͨ܄��%�b�P@�<�����ٴ��5�$g��)�+w�U����ln�)UwT>/G��IC�|�q���m�z
��ADb��ql�?��*-,�n8�����r�=��A/�?������Ko��OEV��hI`��#n�y�o��\���y	g�v.��0q��[���g`ejĚ*�q�h��jy�Ʉ6A�WtYHRO]��=(
�?�+Ir��*+I�e�̕�Lg�/���wa)�9�P�V���/.��'P���z�s�L�, �ƢIĮ���� r|R�U���^�f�\�V�JbFd�7�ؖN0INI*�5�%��n	�TVi#��>���/�A�{��A�^��|�����8J*���x�u��w�Mx��_��3�g�ES�F٠�ԅz�Xצ��LZh��*7��L̻U���DtԷ�[��͊m�u� s��?�.S�(f ������Yp�(e�~��$6%gUj��G�l��앴u���7Q��B�D����	�1�����q�_�~{w�
#Ij �8VUa�B|�������Kg!_u0rf�����_�� w�L�M9!ZT�_:��D���t�6���3p�����?�S@A�n
��KQ�����c��]�#�&��Il�\ ���ab������p�����썜Ü�BT,�4�� i���B"q&$ơ2 �2��HS��o~���z��z1��W�荰�֌4��`�y����t���+f.�~ρֽ?"�k�1H�Cq������q�=YjnSK�=9F�㎉X2
:v�(�x�iȌ�;���ΤMB��0k�|{��(��-A*��ܹaȅ�E<�� �����b���~�c�d�_.��tQ�	��U|�e�Ðe|�ylj`�S ��H�	�-Ǐ��)�6��}�L�N�)���mt��*aAP��(��sE�.�QS��m�]3V��!Io��~G+,�y��T-�����a�x����w�1Sh����v���6�q���׈I�~�6�N�<�mKf�W�[#5�	���J薘`q&@��isp�%W��?Mz�"\߅ǐ��������۫�����_݃O��A�=�8,�,�>R�'�$7R{a��#�SÓ�2��m�p��9_�*{�t.���vE�PVd�%�?(+��D4QRV���e;C�� j^��<��*��x!�8pX~$�y�XK�Ca�:���F��}4W<Fblʩ�u`��6������NB�q9	�j9s��@o��L-�{
���l�b��K���>�2Y�yD����qV�9���c8���Qs�D��hLt�<aq���0�fv�K�{%1U(O������б8�F�kz��;�H�J�TX�e)Q)x�,qE�<�����̒i�l�0֯�0�����.���Tʉ
�����𑳰߰���u���a���ѦPr�̾n��o?�I��� U�lI,�t���\u�m8���1�r��̮B	2��rR6B7��Q�������{�ۯ/�(�u\��\�����4�*M6��(�"Xr��u��1@fç܀��y�8l���,n�U��T�Y�HJ,)�w�Ie��ft
?�P2��0�O��&��S���)�:m[�����=�&�z�TӐ�_B �r�Ģ��S�Ю�+7�[�ᔓ���C����7Pg����&+_x���	��`l�2�T��0X	��rK�2<8����W���'7@��,�=ߓ0��_@�i��f�3[��q�R�_�#���z���[ߌ��"��Z��\K��e�Qs�Ua��a$ɧ��Y6P���Uۀ�,��C�; ]�j,E�O�!S]+B����1��_��E���F1Jn����F���Sy�Sǎ� �5-�(���i��
��f�N9Jw�c����CGLG�n����W%1�"˴z� �ӗ����!,}("�"qMv?�u��P�Jܔ�&Y�.RQE [�Im�F.q�X����<#�����G��'�1�J�T�'�妆p�;�p�1����UF\�)Ɩ7��7b��a���0�PE�43�|��!o�*��e4�������a�=PH�:@�!�_���ʫ�[�y��)�^[^v����&iZ��%�T��(Wc�3;�Aя�1چ�K�`@]�~��iP`�/5�Pq]�S�'��G�N����W�Jꪥ靌��G���[~���?���3�e���mT������d+�&&9Cd�&����ܭ�����!����o������,2��`��iZ	f���9Wi��%9��~��_�EU�e�%mB��}��?9i�Ͽªą�N����j�ap4E"�,t��`�/�䳇�ic+({�M���b�Hش8�-���dd�IL�֪z\T�4��o��������a�ᆊ[���2�ފ"�H�iőE�7	��7�9�R��V�4�?j�a�kS����14H�[p}�:d�?�'?�+������:eɾ�<IO�j�f���_�lF,�IB��k$i\k��˯��y�>�n|�Պx�n�BtO��+ K����&�G�v�fcG����X��4[�ߘ=���\�����E�2np%-��z���rو�^m}nw���� ��Ð:ݴ��`�l��>O,�	�;���I
�x��vx�U٨"_M��yղt˸[��Tǵ2���~��50�3�^�Ԑ"�Ꮠ@6�uGu8��jng��Ƕ�"Z��a��0�bzU�#+�j�P�/iKc��+��#3���=r���s�
C���l˫�D+�|H1�[�����n���Gc���W9��1�V=�u�\W�h�]��n
��P�\��X��/}�����C���Iw�!�C؄�%/��NƆ�ȑ�Q����+���!�ǿ��[����a4-[8��ї\��<�#珘4����0��Z�.�d�2����F��a������.?�/=Oe�0 �yp�G��8�`I��ۣW�mC��r�/n�Wf+��x
�?gMX��A��+�r���sD�p�:�Q&�9CSp�v��4�� �M#w����WV��/��6z���7O�Ƙ��ڭa�}����<�_�aD�ZG��-�v�����f6��o���ϱ�+`�]�d�Z&�n<�2)�^��*Q�&NB���H]���O��VǼ�Kqǯ^�ާO�'�j����/_����<M�`�(i��cH�о䳨A{0fh���?k�>z��)s~�V��4X���p^)�
�9E�����1�����ֽ{�Mm��}MҢnG��&Q�t��X
l�� ƥa8�٩m�H��6����Ŧ��Dyh��R�D=t[2���QU�s[r�{�8U�+��@��媅����A��4����C�Ƚ��%�S�*Q�A����
�����'x��Yx����l{�9=&�� �l��{k���Dmߣd���웴�iKF��n5lT�w�s(���헷�c����ᣦ̽�m�����M6V��i�BP�����;�G������o��x$wi$��ÃκL��>e���,9�⍕�t�yʓ�G���-˔�J+�����r5~�ԣ�α��� K�jx&s3�+Q	�a�Vj�$��S���;��:<Ɋ�����}�ހ��	������ݐ��M�jn���H��՚QW��,����z'5Pn�TO\�;J4��ka��n֜}���5U�W�}�7�]8]eK\�z���a�(�勧}�ҋ/X��P���#'Ϲ�-�����DÐ-3f|&4K�Ϸ��Ƨk^�|�����X��r��ϛ�a�Ð�;��Q�Tqf	�o� ���v�� Ҝ��O�W��7?^�,��5ٕ����H�u��Đ��7������rr{&I�QW/�}\���s���Ƀ$S���-�TrT���
!��(7�R�6t�>�SKf⅗�/��Z�Y��0"2*aek��{��Y3Q���C�J�b��!�S1S������\y����ڔc��0����`�.�*ӸBHè-|�ՋG���b٪�z�soCS�Y�q�z���o�3�^,au��Qml�y��t�Xh{����T,9Q��]�J���t²ZLՠ�i+:�BT����f�/�_�G�2KpP�c�	���G�1z����W	�����Z���ۊ~}���.�N��2��9��ٚ� �S�D�V�!�C3`�[ѱ�!^�g6�!��5a�|�x+np��#�$�d_�P���OB�3f���a���V���=ޤ(�O�Z��T���e"DI'B]�#��e�؈����B�Th�a���������/���� l
�����ceR�Ls�!��-"]���et��	����Q~�Y������j��: 5CH>Bq�
dGa˓W�*�/D�� �H�N�JRړ�=����3�l	2��!j�D��8�op��*�@���FM��ن?�t9�"˸(�}|��L
�|c�Ks���g�B�ϑ�.׸-�V&x��R�hO���,���2s�'+/����:�Z<�&����K��,)S��GU��l��Tl��<�F~��#�ڧd.�1NL���������SK�3���F���c8吽���"<Q�Z��
����Pf!RnqoCT�X��/gl'{ �����w����q�������1&�b(~�,��Pq~{sk
gz>JhTkE�4���V\�	��1��E� ꔃP#q��b���Y��9��Q�x��Ͽ�^�Ǥ�VL�~�b�I�<�%�����^à��*�(q���,���닆a�3q�atw6��Z&.�[�a)/�O�Ic�W_��OE��`4���g�aPK��t��R���Mq�|3�j��{y����?�+w/�/<�/���g>{�Vӱ$�y���J
 j���Kzs�҇0�y8f�upS]QD5�	�m	�!ق�y��D����Q�����fb���qD��Đ�+���(K�Ͳ8�[:硗LG���
�g  XՈ���0V��M��6b�ڒ|��ÈҒ ꑇN�:���"\5c����2�l8i�\�@ΦӢqFؘ�0sҍ8l��(���?%�Z��� �� S-g�<�n�kR+,*��N	G��1���Y��[��G���	�(R*�H�cW[����\5����W�u`ظk���?ǠS`v�m��HO�H|��4�H�����������:� Kⅻ����g��=��q�� _R6:�Ӗ
9X)�G�Dߋo��c |�D0�����	o�R��*�l�a�ݎ>���TʄdV4hiA*Q��s�+]�i���!��E��B l8���{�42Ӭ����+P�P�b>c�Sº��wPnB~u[})�z&�&��CD�Y�&X����ۯ��?�í+c���@$��ċ(�:�PP���~Ç�:��#�Uݱ>�ê� b}��x�����"nC�e��<^h80�[�����2�ǜ�c�)�O��f�N5B.NŬB4,'e���	�N���X�kx�����H��ٽa�Rs�]f���!Z�:��8�'U��y#q�vXF'�_<
�ǝ���<����OJfˠ�L!W��W56t�C�,�����[���V�|4�q�3�D&�Ze�N�@JREt�����+����2#'\��:�uA�\[��:��/���}�u\q�B`�����#N��&_�Nu�rQ���0����h��C�dJ������e�L��1p?�,�Ejy?R���pH�����G�B��C�1PV�Rg�$�D�uC�-I��-����&�Xq�CGM��`[BI��j�ֆ�	ʨ�c��1�t��8f� ��BK�p��zI���L����s�V�~��<|��}���ʴl�'$�����Q��/���c��*��	��6`�'�b���QX������_��i+���y�>�Px8�>��C���5hU��T�@L�    IDATv��/j[�|YÐ�'ӗR�ݍx�q���#���n�t��?�I�R�%�w���Y���л��KY5v�cm�|2�n��ضy�{�o�-�6@e��j��*܌�n�p�@�Iy5�F��җ�q�&���b�������y�NZ����M�v�N���d�@�i1ތ�����(5"��r���I+�a�6��W*ɺa�_
������ �,�"85]��)4�
"����YxLwiINQ�!�6�e��uQ���f���f��yU��'���
b��oy�3�j��+<�I�#�DS�uh�-ø����9y��m�I#�$�$�gV�#P��6j-]䤂����#���k:�.қ����0�ڽ��7kD��8M���1��*E�|~���.I�uN�q5���eW���Dl*�(-�2[�wcU�2�l;KXI�H�6f*��\�L鴃b!�T�VDg�b�Ȏ4K�)x�D�7 y�������G��v^A���0SҊ�����Q���l����Ɗ͒����7���8a�x��?z�Isi�aHqse�9�/]I��V/�aK�wQv}�p�TZ��n�Uf��e����7��s)�M^�@�	U+\���0ĿDj��xϗ)-x�Z�a�@x�Iƚ�����2%"|#�J�*��jh*9qY�����%�({�+.SC(�)�B"��i������^]�2T�`"���҆�D_����0�4%�,J�}��P����/H��F������E��l���\*�o\�p�=�1����Dn`+* �x%�)���[�JV��(���I-#�c�z�W-%��7�+aS�J@��@�`�l�/��YJ\���c�8�Ed�iY�XM�1����lPF�hq]�G7
�!��s�َ��[P�'�<d3�_c��-��n�3��=��T]VAɲ��	˟���YK6��G(�x��j�RN��H��*�P��(��0V���٣��{�����"�3,)����Q��R�,d�Q�U�M+Q+Hq	�j�t�|p�4t�!�����K�-���*�)T�.%���ϝ<��|��z�ghJc]QI2�(�6��&�@,+��Mtۅ��W'7�"6a�)�*'o����s�PQ����w��~.{8�c�ՠt�(OxL���*I���>��-9���B��)U򲖮g�c��0��<��6 uڮ�|�����yLɖᯠ<]�Cn %���{�*�bY����IOD*'5�J����I�9�O���I
���~�����8�I�TU�A�'��.zn����JA��Ϲ���8�5uSI>p_�]NI�ZA�c2:E���U6��A��[11q'��/:|�ra��Y�}YT���vF	;�dُ�eΐ�0�ސLSe�[�S�>�T�J�/���=��ۃ.��$TJ�"P8Q-���"5�u2�(�p]��Д˫�C�k��#�
!��Qln�ϕ8 �R���U�r�I}c)���u't��l�5!���GVg�Z:V�_DZK����;#W�s�0*
קw��`%
�+wI�It�p�M��JjE'�	p�����P��KlYS�_��JO�PjY�đ!��,�[U�7׀�AI1Ű^P�l��Q��N#�z�����qJ���W|��A�("��bI�%���dm���TTjB�Y��aC`��pR5ꁺEX��M�$E������VXB�a�{�Fs���	���<)���q_Z��Q�b�,-M��*�JY�dYF^N��ٍ�A�.��r	�Cɍ&ľ��d�#>������_B�LŇC-.�������+�oǥ� ��j���-t���lM5�%5��$��D�v)�3�BP'�7cl+�<�n I�%�r�H��������D�c!�J�c��X� D���*�8��\��ݺ�Cڑ!N�4:o�/b��*E�y(�s�i*GH�����|^Z	ZA<�DV+N�K�	�S\��+�2]�d��=w�l��x^#,ǂg����&�i��\��|N
�b���t�A)�jH-V�|G�%a��'�����Z:h��fb(���$r6+��0@���s#hl����,XF���Q���"��(A�oy���k{��C��*}S��ɤ��,&�erZ;B���6C3#)b"�M9�BH�g�34�]��r*�R2m��!� ��u�䉬�,j���؉T@6A.�T��G(����t��ư#zL�y�"�� n䢙���� �T-rVHY)��y���#��p�ɕD����p�+8_ �+�'*[�Ԭ1|��,Sl'R<;L��������\��Y(�Bx�S�\�衐;��P,Y����0ڷp�2k�!koE���L`*3-�F�F9����7���	U�#d�.̭nIT!&#���pɱ)�<ܮʺi�2Bu�٢���"���	�R)�~lp	P,�^��Z�\>&�
q����p#���b�ơ�eSY���c��)4E1�t�B�P��R7�Ur��*�&هm[s�4�L#Dѣa8r8��Ӏjzٲ���PE"�#�@���K�BB}i�E�?�&���P�&�ؕ�X�p�W��P7 ���F������&��0��'aӨ��oF��	���i�:��YzU��CN�#t���e��\C���
��ѳX�M�Ig�d��r&2`���.�ha��e갵"
�m��nظU��u���T�[���5Ǉ����a�a���(����1�����Q<�L�Z���zҠl�% a�C�ə�B�sa��<�xՖ���|��W�P(QۡNr(�����\tѣ�^H�r��l]�X[_�2����پ���|*:B���b�Qx"��͓��B�ۄ���ǡ�Bm�Z�������+��ߗ��G(4n·���y��?�U.oP3��zϬ^O�@��p��4��طe�ې��r���W=�[��;��ף�Cg�|�x�w�A��M]R.z�쁗�[����c�늌��J���{���O�0�����*ui�������L�]Y���]�RN�����s͠���c��zⵕ���ǀ��q��A��^��	��� �WF��0��1x`?4or��k�fK[K��/ۣ�ve(��1M;i��h흮�
��*�4�f��_@��Ƀ:�_o�<�V�
|��s��n�� �Y�a�]t�i�k�:|��'0�4�[?��}7\�����!���%Nxc}�B�湗�i<�*�IT�KRjVa�bȡ}1qTo��%��Qk��o�����⋿���	=�6�TzX{�!�p�/q�Q�b�y=�֫e��� �����;؝��h0P�\��ȕ!"jϬ��pr������G3�E��
Qӧ9�����{�O1�GCq�`/�=Ė���l�r˳���p���!p��/oA���e���^�V"����Si�k�1�i��3NڳRs;�:I��ت�Oվ�����}�&e"�o�ms��+n~~�%�Aˮ=/<�1~���y�yx�X��x�ݷ�ǣ�OŲe/���`�Kw����7�?��&�u�,�Q�A�.�uK03���������O���4�P�fk��z�zv��o�}�æ='?�� �&���&�C���ptg�x����p�����b՛y���ߠ��P�!ym���zbA�"M덫���s0e΋�|�m�+��߽Z��F��� ��|�࡬G��s����Q_���?���A)@�J�>[�T�!�7c��Y�}�y�hm[;@Lڃ��a�a(JQ<>����5�,7c`�z\x� �h��t�B���ۀ)�5�t0k�Op弋���>��~�Щ�߼?�w��7�ޔHےK��-f��t�s�˿�՛�j$��������]0��>�A�k?l+z�ׄ*�N�����o��Go�����ƕW��{�1v�i�h�8��#q�{bܔ���v(P��C��o���������0�(����t���Ȕ�a��`d��Kđ}�a⸓1z�C8��� �ࣿz
MZ/�4�L��'��ϋ��{��#��R���Y�w����� U�EDε�+��b���G��`����� <����۶YI���Y�ڔJ�*�GCC�p�)��ē:�򫟄�aXv=����N�|����Y+p�Q��ck�v�68���#�����^�S�d4~��!X�6��~�
�N7ԊDX���Ȱ
�n�)͍ͮ�p�1�����p�#(:�6�[ؿ�<_�z�s8x�!��I��}�r�y�x���b��0tԷ1�ʟ�SO��'�b�5� �=K����8��#pѕ�0LQ8����4�SZAHIM�oވ>=:b¨��r�
�6T&���ߏ��Fc��?}���3�����em �~7�$̜r/>3{!��yW��,Æ�!#����c4ߵ`�ɗ���n=���>r��)s�i�a(�E����I����3~	��	��Maܘ�8��G����M�*�0컇�G�,��	L��,<�Л����ix�mx`��~��V��-�p�����5�g/�OwGFKJ2͊��`�-s��T��{�`�E=1}��0;tG��ѷC��c��ᓟD���q�=qͬп�>�1���ﮧp�ȓ1lگ��O��N��u7��:[7�ǹ������a3�v_�Q;�Twdc�8� ��G@=ִ-�qż�q�-´I�`�m�����̪�Z����93��PFA�!16�r��(j�I~#�Ad�� )6�WQA�A��$�2 خb	2���9gN��f�ooa�k�y<O���o�o���U�������ˮ�h�_��폂�C���hށUs/������� ,�#P�H"Ef�^R�j��|�;��,
=4�_'�|��lF5��&^��lĶ5�u�ނYS���;_⩗_�-�]���X���֡.�桤���؉��(�ɜ1���h㞧6�t�f��D�T�7�@�9b*sp߄JQ����s���*6�F$�Y�%[8nZ��8	���7O{��è���
\��Ӟƙ��E��;`���?�d465`�X���Wo�)d���Ty�H����$R�Ԝ<�&����8��/ ��|��qr�1�:|!�pg$lb!���fa�Ⱦ��ۘ��i4
:uA}���i����w�+Y5��T���dT&$;I�q��ۋ/����w�植�N��l��]9�3z�聑����{@m��~��x�=��e/B���j�6�\$����/C	���5@���WS�:�.+M�.��^��/���kZ�9�ǅ��":�U�:�L��7���=�`~'��v���D�;�9�~֯q]���C aǝl�R�c �,����&�M�g�'�OC�)1�@N�[��_����_�� ���8n�Gu������/�@���]w\�ʝ��-@^PCYɚ��G,�h[��A�h�b������?���x�<J��F�����>5�t&o7�P,��%e"VW�ӎ;'��S�s�lM��w߆�`j9��4qF��(������a��g~->(V
�W���슛H��P:�+�Ӊ��M=I�yU�����il7"!�\t�! Yc`��j|�����'�_|�vN�]���rQTt$_�ݏ��~�Aꯨ>���d{�
�
EE��A�� %>oBN���\��t����2�G�>��O?a�?I�L�`%�����X��Zl���d�p'��D��g$-��u[�O�.֌PN������V��c��C�0���=sU)Ȑ�=��a#�#��S7�7Z�P��H.o����Ò0R-h'�nG�D
��|dH�D�3
�$d��*�����,�]e���P�ށi���g"9~�$�k�!H��$� O�Y��h���:k2�0-)�x��.|2R��P��Ɍ�K�$�3$�C�ɢHc�g/�t$`D���#�!��`�a�`F"[63�8`��z:Ú(�t>Ӏ�hJ�hױ�Ob-[��Z\͖���,�WXۢ��j@E'������I,����S�1�%f�4$�..�O� KBʰ�H�Y��:dL��.)YZ������=A�I��_h����Q$�Is�n�M���1H���a�SU0�Լ�?�d�ivj�z���_VGtU�\�J8Sj�;
�J�+����룣��b�ϝ���$��}�D"P�xV�	^�t�NӤ_J�K�=�ᙓ.1��~��č��L�#E�J�%�_P\�I�E�uN�3`mr�9V��S��G �hD�~^i�����iK�(E\�J|�t��n=��A�Fe�!�q�Rw�J1D�#{�l�4���N��7��*�ihhDT5� �GR�<$�s�1�p�Ej��bP��$b!��4!�#��ޑ���Sy�&��V~��AR��X:}!�u/DP�{���1�5����o����͒2T��Fm!��4L�:�&�i@*�+t)H1UN	�)�����P;:'Ľ��� �cW4fd�dd.���E�r���
� ���A��X�6��,�6Gy"�VEgԃ�y�Ds-l"f�izNw(�����<�"��$�!��7�0�X���Cد ������)��Mք���@���}P5���BGSFB�{o4e迉��f|��+p��/�q�o���q@�X�xŐ!��~��u���<ڣ&b>K�M�r�B�I2����&Rk�L�KuDVO%qŁx�|�D���PvҁBH�KLx�� ���[f�F�IO h5��s�t����"<j6����oݠ
�C9��~�<xD�<��A����뽨�	(��P�l&Q�y=��z�A�
�����T>�z<*)�O�r��i� �
���#1�I�>��4�KV-wׂ���]�8��/�:�;_Bp>��f`��AX����hx���EZɛ�"�[�E��ۣ- a;�G���+��I�?�I�a,���&�@��rX|:�:7㍹� f=��`n$�H�o����Ť��Fd@m��Jq�)��QKF�ʢ-�w�s/n�!�(��D�R��jT���J���Sg<�rIz󎞡��AHw�^�g#�+�e��&�q?�W�+1֔��E�7�c2��G�n�@a�
}t�/q7L����B��F����z�|�r��@��:�o*���/�Y��v�/�NG��)���v�N��=Q:�UR�%oefP�Ϡ�ڃWg�dvv�}#�-qc9�<�n��K�N���'��[�#����x��;Pc�:͊
_��M/a�ߖ��i1��j���9�����<�j�1�aĔ#��d��1�Ɣ�]�{&_rݐ���1���l�]��j�=����G
���$��AnN�H"�I�����������V�G�hE�\(�&�i�Y�G��Q����
ӟ� w���Q��4m/e�\��#�nDAf'�?8�l����+�-"F➠6W���Px�(��	;��,(�R>z?ϣ��qB5bϣ��ֲ槫Q�z)T���\2��E�m�SN��~���Dq�	�OX�z���l/�^�Ѳ`��K�J��,��~脻l�a����]���*d��i�J�Sȓh��2v�0�ټW}�{@"#�%T���$��΁T����v3)�������8��(�[[!��2��jtqvc��I�̯�'Jw[���d�Fb2J)�.��ec��� ��c8v�M�����yXWI��9zқ����j�3��l�db�Q�~�M�DW���^�}&,D����L<�����y3'^:|蠊{�%+F�������`��#���?�\�d�t�eu�[
|��1����^5���9��AWE"o4�A�:�R�T\� }�Z7�=�nԨG0��x�i @d#���$�G�N9v3
t"Z���=q`� �m��N]q^RC��G���Ǣ�	�!-�p�U���*Hd��<B�6ȨLGF;�{�il_�?P�Z��G
�b���)
t+-T=�b6�|��a1���,���<y��g�gM�lXt�ڃ��c���y�bh�����2���
6��Q����C�l��b�s  �IDATFِͪL�9̫�O����nGn��ۓ,��	c���+� �H�=�N�)G I�*�]�(���3]�`q�a�|,-C3�_a��ɀ���d .}��%�qR��ИHs
H���=��-_����j'^6��)9����<N�x�]�tw�����齿b��_Q��4���i��B$'i��k�][��̀e�^��L-DѠv�ek<}�*���0��gM�����p��qC��5���Ὕ�C�C�TB^sg��BQ������nA��5�[u/?�{��*�s=��B�"���9���$ʮ��
���l}�ށ:�I9��*�àݤ�M��J�Ŵ����x�̀�`6{�7L�������$��h2&���;����|��)9���^,A�S����a����"D�8��]�]/-㬈��4HE5��KW�b[&��(�q�5�����7,F��6Iw1-D[�.?Ʒ�h�y3�\6|h�k���ax4C%Z1u�N��o.it�g Ό�ͯ�n�}�Y�����N3f݋�Y��F���rc3�=J:����W;!)繴��+ܹ P�u\�#�k�l��x�-�U��l�d�c&��/N�	���-U������/�~�0.����EF��`(٘���<��l1F.ZP��*�~���HN��^��=�P(���pn��FL�2ŕ�d J�:i�#�X2$��ګ�������ߑ���c<�h�ء����m��
�8�:/t��n�+��v`�Q��g��(<:T����.��nhsH'���Q7s f_�d��^툤�+��jyj͕�o����i �đkVc��[������N�8}N;����"5�n��TTn�r5MX����@���c�:�^AM̮�0���[B�(Ix�����a5p�̌�2p����ɇ����ݜ60��1"���.��	}&>�_� 4��<]�	��e�fN���磋W�:����b��9=e�m�l�@P���IL����"���M�~�Hv�p�6�{/��LI�SX�2"8��<u��q��Q鈔,x@|^̊~���M��l�#Ϩ��{ou=F���ɓ�3�N�͚�A�f�uL��fl۾�5�L�.���aPZ*�ἴA���D�{A���%a�?�]lM�㟞t��#77Eg���`��񮖊�j��c,A��H7@���U~ �.�X0{��MW�Y	Sr�H��/	������p����QQ0i h��a�z�(N����F����E^$��:{i�h���PF�낳�ގ�0Zȭ�}o*g*��pD~b�a4�Q��>2�� US1f�H�:�'�3ҀM�O�6_T��j!
.��ǟ���m��6E�Dɉ����.�,�� d�a���M��B�F����9�AD�~�-��il�1��[�j��`��`*]�{�c�����h�oo�2��0�g�E-p-\�l��3�5�Ԡ��y>x��H}�(��"���3j����>�OйK�)��2"]ݼ;V- �Q��������Da~G��I9��Dݣ��Z�;�N��af����
���^����yX'��݌\���a�vL�q��ĉpꩽВLs5����4m**+w����^� �/��O�+uk!��%�'�*hH��->Z�J1�~�<����0��н�C��8�&��Q݀&L� �|u���LZ�G	���[ܶT�@G��3'�f��A�������1d���:f1��B� �"[%4�jc�H)�$2v�8���EB��x�ILA�C��+��o+�[#���m��~��ܾ��& J�R!?JXr����Q� f��#�[�`��k`�<ͮ�1����(YM�:��D�8F7�pN<�R���ɓ��˯��Ћ!��oJP���#��ʫ�z�5�����a!�ɼ~��_���|���WCs��~����׎'ۉ�1na܈�P�[���,��g�{�Z$-���j*�-�د�x`L˼{n�p��?���hђ��f�;u�b�!�!���t�N.�D��# 9̚Gmwj_s���W��p4��+��ހʏ6��:���D�@e�4f�1y9y��Q	9e��~�.|qT.k@�N�f4�"X�|����KɃ�^��8��g0:-��[K�si�L#�"��O�N�{�Yl7�<���?�v�r�(:�/�\�L�EMTQy���� 4�]i�(�L7 d7a���hx�9 ���W��W%̝>EyH;Ҏ��Ҙ~�T&���A��:f�+��˹/��5r'�����W��X��RR!`G�<<��~#�^u`������J��=��腨��9�XA�H�
zE	zBUO:k�<%w)PGn���72�US'����4�15ۑ�݁�_�q�m��|�C3|Mq�hV0�ɷ�)
����t?�$�I��a6\qxyi���T�aI�B��V-��ћ�h�4�4An�`����[;���)��ၥϠNꈌ�"��1m���w�*h+A8�#�bQ<INQ^�c#�qXB��d�64�4+�;*�D�ބ���F��iX�j�<,{�%Ȏ���g\
�[�~hQ0����b�i�6\�+y^nⲼ7Q-Ւa$�Ϟ��`����2��G��^�Z�0�����|��xR\�	�G�ܗ�Ӄ!"[p�A@��Y�rXݝ���P�8|�ǥ�uC'gBH!c+h��o6�l,[� �a�*�Ĕ�� �i*�*n��%ua�rFES�=̀^�j��'�x��_��_DpT ���3о+V��5��Ѣ��&+H�M�ׂ|}2�Z�Ȫ���b�7��N�L`!��Q��Lq�T�z9?B�j�?%cd$ah��Fg��h't҅�#�|4�R�\�LT��V��X[>�c�wЁ�K�K���Xt�臱G��L9��vQ�d��K`[����e9�V�!PR:쾴9DWd��Aq�����?V����n�nD�҆�X�h�Y_��Dn�%aD�C�0!�e'Y��[{o�%u!yo��\U�M#�To���A�b@�؃�����SKӬp"�k>m�6�H4�aPe�1�d�Z-n|�``�;:Fż,W��`��~��A<]�%�"�AH#nA�@?Y�Z\�S]�j` !��Y�7+chrr��Tj����ԓ|?���N����?��X0s�Q\��ɒ�	w,9cԃ�E���Jf�u=�bN�Ĭޔ�w��kx�"3/$��QUQ�1B�0�ڨ'��[m����%�B�ӄ��BS�x+�Ӊ̎��6��@wJ{Ncm�Hg�P뷇���!��OT@ɿ��,�X��HT�z��Ԃ�0�p� �C���1lu�Y��LC#V<j���%X��� �hT�1�n��qPA&4oBG�_��'<'�nu�j�n-8©F�6�R��:� w�V����P�v2L�B�Qj��Ϸ�4�F��ϙ���4�=;p�����9u����kR:J�!i�� ��y4�ď3� VR&W+��(7\)
⤢a^����
�=�Xa�@�"�m���q��հ:�Emb�ԋ!��R���0�.tq!�(�%�����ꋄ�th�@q^�$��MBK7C�P�/�+��?2a�
2@�.�uT2E�)��OZ�:�G"�h���O�.���,���	K��Q���I�Ȯ�߲A��NG�zo;��G#)E����� 	��j$b����"Ø;鬃�9�[�������s���!%^|"��>Z+�)�oA�����`0h�T�����+����l"S[����'�ev!OR��R��v��]ð�f���ԗ�!g�2�K܂�[�̟H[lK��k$���'霐�[Nz�.2qR'N��ĔBT|^�]Ng؁�0b��]�k��\��Y��(��@1�"�3�9�KA"���Y|>������F{�Ჟ+��ԃ�S,_>vJ�x���P{ �(6���H6��Ȥ{&�Q������;MX���g�|����[{�o�1�_�X��7�|���	r�׎)���G]R�GG���������X��"��@�K%=�MkIЬ"j
����}I�p$��=)}�v�|��7D��,�a����baL�����a���� E)����4�:+�I{����"n���g�Qk	�.�a�U7p�K�C�Ik�R6E�����D�d}��m���]����6h��io�)���AȖ�%�������:́h�[<��j�	[1�8���G�~�u��r@Ø����aCG�_���Upu�!�^7���&:>F@yT�8$�I���k?%@p�t���J��>���fh9[�E'� ��Uu8���p��I��Y��ɓ1��
�Ket�# �����1����Ҙ�S{��h����ѓ����θ��*B���+���D�{\�s��Һ�b^��E�Y* V�<cέR�<��dd,q9�I�ǘ���縮Q��������m����_��;������>x���_NsD�ḧhɧ��>��J�O<x�Fh��l����8���{�Et]W>�l�d�Q'��*�5ɤ��q'�0�w�ޱj��W�8�T��'a�R��;/���^�2�(��<�k�C���IP��C��q��a���85�����"[��������K;��Uv��=���Ϸ���_A��Y�耴�-��{03���8tȈl\�ڗ�;�zϞ�[2FWJ�e+u��訩�X��X��c��9cq�#Ѐt0(4�dI����:��a�u�i�C���2i=S>hH������믽�s�����G��T�u��*6�ߺh�/��gg4�j'�B�#� ʝ2�ʁ3���am�/���)SK��A�*�x�����������Vm��9�8�	��oWvq6֦5�/\�(RJ%�|����3h`tB��?�cٲe/�'��;w.B����ß������y��WJ?���Ej0�I_S��MCˆ����i��O<�L�/oQ�J��}���A%�Z��6������-����X���������yc����غm�i�T���%%W����c,_�ڱ�I�I#��+���?[�ֆQ^^�aƲ{R�K��۟�����ͩ�xm|e��\��ҷiVF�����]�x�0���RD�����0p������4���P<�h���'g��TTT������+��vdn�F�?��ڴƊ+��u���{6�yqq���Z�p�����k�0 �[RR�'��v��몪��2�O��hV��k+u]���a,)...�ƽ�o��*]-//�4�KZ�[%%%gfcs֭[W�u����cS4�Z�bŊe����p=�����ٸ���x�4�K[ƛ%%%����ُ���FO���n���0�b�0��������QB�eY"�YUU�@+��m�x�0�?�������o�ˆa��*�|cp�
\�	>?�F�=��ƮX��)]���c�_�|��0�m�16�������SQQ1����V�h4�+k�+W��K&���ceqq1-��s��kM�����8뮽�ھ�ؘ�k׎������0ލF�YɈܬ�]���0/..��{�O>י�yN+�������llNEE�����٭�h4zz6�v�Y]�/����=1p�@N_���˖-��,�W�b��|^66���bRee�V��v4=#k���뗴�Os0z(>��a����(�5��nݺ��n�z�g�e�UZZ���k�u]��3�@ �Ԁ?����(//�4��Z%�KJJ~��7f�ڵӪ���t�]����...�2���c�d���"]]�n��[�n��%kt]�x��?<=`��+~4�1�Y�Z峢�bzee�M�0�\��:g`nI����bN_��p�1�5M��CT���������0V��P�yXƲe˞�,����&�V����5�\��^Ɇn۴i��P(�m�T*�NYYY6�յ�a��y^E!��篺��~4�Ix¶��4z�r������|޲e˖�Y��DjL����Ҭ����� �G��~���k��u(>���X�d�R ��(�|��ʊalذa��͛gAZ:�&5�#G��e�ʲe�^�m�"�G\�OF���� V�\9'�J]o���ܹm�ϖ��e�Y�f͠>�����;��pgհa�f�0V�XQ��'I4k�����,���+'fk�o�sXy����Ζe��i�i���e��nݺm����ܹ�g�i�h��b�f�QG՘��w��A����$Ɇa4���U�=b�Z��6���Q%�H~��8�<�!ڃ�����92f,    IEND�B`�PK
     $s�[��/F��  ��  /   images/0c7fd013-2f4e-47d0-a46e-2d19cc1fd6f6.png�PNG

   IHDR   �  w   `�3�   	pHYs  �  ��+  �RIDATx��}��U����קd2)$@� �����T\�����b�����E,��P�� ���R$"���H�(� 	I������=��޼d2d&�̲^>a޼y����{�=�{α�o�oc�o����7������a�mlpL�X�h�2{���;��C����vuwT������M_r�G.3#�7���{r����S�ryJ:��l6���^:���4	�V%�;���+����_��W:�݇�xo��<^�̬Y�h͚5�������|�~t�Yg^~�Qx�����n�i�뮻��<����Ţy�G�iQ��8��>��J����EG}����z�U'�x�[c�[�0^xᅶK.��w/���S>t�G���_h~�c��ܹs�������2���$��r��U�VA$�ʕ+m>mg���=����}���a�4I�y�w�%�\�N8�����{  �"���ðx���Xx�]w-�߃/�˟�袋�ݒsߢ���/~����2�K�~�s睷��OAX�z�J�P:cӚ��3[M�eT��aX�:�Y�g��]�����y_Zh>��C�O���3�������y�{i�������ۿ��M��ַF�oB,�H�;�:����x͟����o^�/|�7�cKq�-B�?��>����[n���V�s�=ȶ]�
E�811�T�O�G�kS�=�����p���}��ߵ�#�M�_Yb��GWg�(֞w�9�����O[y�������%�a���i&�7����'���3�8�ܟ��'ߦ�<6;a������΃~~�y�O}����I�_���~�dSG�'�Q�t��~�_�۟�̙���t�9��KO<���7�p�?�V?�p���[�x��)8���8���E���i^s�5�~��o����1ڌc���W_�3>��;������~����W�d�!C��Ü�cvj��5Qlx�4�+Ez׻��'�x��k���eq��%�\�Cڂ�Gi�o��z���;�^���(0p�DI���QVL_��O�����f#�~`���8���{���ݱ�ڊW����5oGDF*���6zF�^W�"zz���6���S��<������k�|���?�����Rɣ�O���F+8��Htp&�f]�7,�~C�al�`�#�J柿��������AJ��S�d��XB��@N������<�0`"��R����@L����4m�1gΜ%�C�b}Bh�H��燿�c�l�6�(�_�hQ�����	��,�q�Y�����6�=���a%�f�����,�u(m��^k4�H��T��(�ʊb
����>�Z����~��G?N�q���o�Ή�MK,���Ot$Ću��j��q?&볟��������r�`y��~��w���[y ,�G����dR�_�@��,�I�:�@8I �bq����s�Y�r�i��}������?!4/��%N�f�)k(\����?8� ��9�y晃|����r�2j�h9a�t�qןq�)4oގ"B�@��⹖-?+�
i70mlݒEM	a$��d�w���ݎ>��c���_/ᏜH�a|�+_9��/���KNwB%��"�5A x�������κ�?�j�h)a<��s����{|���Z��+5�>��w�5�	b#�⍬�t�^���H@H���t��O��s��i3&�����4��$����L^��%K����vۭ5f��0.���?����B���j��ƺ%+b0Z�p��'�e2._���}�s�Y_����Q���_��'�l�$�h�����-3�[JW]}�	7�t��=�V�9E�w$���R�U)Z�`[)ל�j)a\y���$W_}��4	㩧����=�n���;f)ŴYG�)�3QA����}��ٳ��|��ߟ�{k���Yok�!o��④���Θ={6������6��ʛ�c$�����s��丆u��w���~���������`%&���"�E�'�x�Zqݖ��z�#|�p�χ��(�ٸ�b��9�ݬ�a�
�,�ŋ�e��`%o�scJ��\��w��ElOO���'''�Q�eaX��b��R܈^t�A��CصU���|;��ΫV��@<��cq�i�5[FO�����9waÆ�o!=1O7���''X�Cs�8�9s���gvn��V�X�GBo��Römѩ@�K�.ݱeץ�cƌr��`��6E�Y��&n�vp9@<��N��ݴz��Zu��^{mF��zk�D���\�r����n�k4����n���v�A	�ʳ���Y8�r�I�1���3Zu���y���	CɾM��L|D���I�ܻ����fx��&�fs�&+a ����m���B�44�u<I�8u"RxN&�����e����(��0h+�u����M���{����I<ĘDb$��y��f�ey���,:F�Di+G�y��l&�ɇ��,�Z5ZnK&hnِI�~ɢ�� ]C������G�\t8�@��c$��pQS(�b���dA��fc��|f�@�1"[[�4�AFK&�RQyE1��5���
����300H��J̈́*�O �	W�8��H�����?1<����Ds�K���2+-�}�hp����f�ϙ8��3o}c}����\=�붌0���Z�!#�-8�4���A�@8q�v�����^.��.gC���9���r��	�ɐ�$�0 =��,˥B�P�c�%�#�$
�h#��l�ha�p�+��P)�d�-�n���E��b�,�q,�cK/p�;OVrVK��q ���4�<�!�`n!��rU�pŃh'1�To�s&9��$�J����i�ò��G�iG���pY��J%l�ǜ�䵵A0�6���@�=��N�)�O���;;��B��){Z�D��g����9xUIIĕ���ʥ���N�9'��9ژt���D,�)r�J@:�E]
1�F�o ���c�Kϟo��_��;�h�5�6�`D3�T��{"�p�iӧ�?��:�5%�ϻa=�S�d��-�-�1�'@�mSM$.rȾ�����|;��|��fϞ]?��w]s���9q��xԑ�w�GN���;�8ꨣ*,\^p[�nV�8X�/��ne�F��D2�ň�Mx��t�mw�׾��2�����p���W�"	H[s`���[r Z�c���ğjU�=t�O��m7�U�t3��4>�K?vʩ���k�������~�/���}h���{�;��v?&�4+���=������7�y��@���ض#�H�8o:�pL6'W2Z�i���&k�*qpHM�G��_͋��,:v��W�.~����¯��7��v=�����8�?�o��Ƅq�㤎�5�/)�9L�n`?�tJ�D�����f�6)ul@rj�i;�/��8��aۺp�O�-�e�Ϋo�麅�v���+���/���1������ʆa�`�$u4p'�d�Ԣ�-�N�g2�|	��d���c��W	.b�h��~3�h�X��������q��_[�^��/ް�N;�:��!-�Gn�V����c`4ńZr�͇��)�dd������;�v�u?y�G?vƒ���g}�/�4o���Oc�������;bƮ�5�p�U�!�}$���%`�W�a�7w�r�/��r��xξw�}��]��/��?劯~��Oo��дz��L(��BVV�M<�8Fw+���	#����s���=������Ww���;��e��Ѭ*\��u;I8���u����%�`����1��m�}�{�\r޹�]��.�={�eW���oY������1�b���%~�@�*�?0&��1}C��'?��3>�i��?�J�6
,>v�����u�ǎ�N(����ئ�@���ͦ�~=I9��������0�/�����s�����Cl��L���PTA|�u0�ZEbu-�7%a4ڙ|�!�F�W,�0ů0�~��#�f��a��'�p��Sn���w.\x����ͯ��l֚l�)��?���%�.�a[0�:�rW�S'{M>��5y��?9s��#�Ng�V�Z��o~�۷^x�E�IE��
s��խ��shp�֪�1�6Y1��x'��~�����A����.��9p�8�1��JW�Y��c�r4��&�X�=�9F���Oj��s����s���=�<󌫘����ȡ�������<�OB���9��0��D���G�͜9s���5�;����n9s������)V3��M��F�_$DӼc3r]�b�i����}���p]�*����n{<��7�Xr�Fͮ�̥E#^7�n��[9ZKʌ%
�y�<O��bq�����M�z�u��l�o���F�VϘ��dN��m��ZB9E�1Ls�V�PEl�g��9�m��.L,@�nR�'��ko�w�̖��d�$Y��N��Y�2�2��);_�1Fw�01���Z�㴮�ũ���e˖e�I��~�'�R6��Ea�:�C��δS�7��sX�R)�OW�ߣ��[������3�<=�Ѓ�����a��0�D$�E�b�?�R�Bm��F��ߴ�%
UK��8����������k��RƧ>��k_��SN���SNy��]���o������D�*���Ȓ��0&��3�o��V��R��^uC����oe���対��Q�}�����NZ�ti��;�8nqk`j"�)s.I<�5�MǞm+[=6��e�qI�]�,tH�Q������E�_�S�Rؘ*oZ��0Y�S�_�٥���?w���y�G�������s�����b��re�` Ҕ�S��M�M�16��L.� �@nj&���d��"a跿}d��~��Z;�BVG#����Bt�i��p�����?�~�d|���G��bT�������1g�Li�500 �o�m���Z��e�]�p�%�Ă}cS��x�)���'�J��A��f�1T�WZk"������\�믿
�DU���@.{���HED5�u�*�EIh�������ъ�C�}��-�@�R���䮩�b�������A��
�a{{A��_
,&�䁠�	~?����z�>2�E�d�7e��IŜ���*��ۻV�%%�@���(��fh`܊봮p
�$/��v�$�K�'���Hg$ҟ1�j�ƍ���˚��(�0�p���5�؍��0WenL$�\���	�8��c4�1�S��jPK��~;Q�uO8�1�J���h����8���8~����`&�k�U�u�!�>�ĸ)R��c�j���)x=���uK��Vr���I1`";���̶'Al�oܦ���ٔ�k�o$z�By�ιNKJ�LF�h�WM���uG�Ҟg�>��0l�YՊ+�-���O"<�~=��U�o��#�h�Z^�>�c��Sa���cL�X�dQļ�-9�X�x���-�Veܵ� l�^����L���X��Y��Wl�h���s�d�+Y�¤s�� �N;�v2I�Os��78����
è%�d2�f����i{{�@+�;a¸������ř�>��<�(�j2Yq�o)te�\Τ�����~��ex`�6a\|��Z�j���^{�<<[���':����UW]u��>���o_�`��M��	�#�Xj;Ԩ=��pR�@d󛬣ӦN�J���B8�?����p��_�c�׹�;N`>�T$?��{<��*�-�܃|{��C���#���?���i��0C	���8�t&�/7��,�>Dzz�!�7�8�+��leSn�H�:a��$��$:���P(��Ƅ	�Z��(�b�{'�K��
�o�N o8�Ht��cpp�mS��Nr:'�� �JUBMz^�D��&`C�rH�q�R�\.	xk�4@�X��k�x���r�f�Y�(�[�2I��V��'LȎ0:�<��@:)�R�,S�M@�^_�]�1i��Ġ�F��[�ӗFI&%�L�HI��tOE��e���D�1h��1�@�J������iH�#Al ]g$����0��O�t�ϲ�U�'��1,��@L�EO�\�%����	�sM����w7����,@ {ǟ�ST�BJ���}J��3?�,N�s������HH����wS9�����\�s�ąw�YoX���&�a����&?K����D���g����#���)ND?�*�)Su��b�'�3��L�;�ǡW�S����:H���xA�`�a}B��'L�m�N�u�������2i2� ��g��d6�c��	�f�!ʘ)�{ȟ�MaP�Uf��R�n���ɷl�XS�w.��_�f�đ"�Q8F�"z,e��'�I�Q(VM����G����uV��V�R|6Bз
���xD)��a��cC��M��Z���.�X�0�`���Pd?�C��a�:���EB�O�0�8�>����l~J*��j�Sh��3x�[)?��v�ƺ��N	�gx�"^�J�L�c�x`��0�+�O\��:,�׷�I�*Lm��̘�*��e&�����:>�`̵����Z1��e��aa`x�n��i�j���<0$��P��q�S�x�@��d���ab�ۓW�2��	�e�vT�Lc�p�g�͟*g̺�W�L�$�0a\�݋�����|�s)'���Z���d���~z������_�P�^ه�"k!4�����e�[��^`���:`�[5��&ˈ�}�&Fd�S����a��hC�D�k9�m��n�F�U��2�D��,�4��BoQ�^����C_���ڔ�|���O��''c�3V�Cx�s�]{-}����ț+�`����\8���+�h=����++���������|����Ь^�����+_U�}&5^��yU�_8�4�1a�8���y|�������rՊ���N�M}���'?��<�����[�CF�Ȼ�������p/M��5cƋ/�Y]�-E:��(���ul���,5$7cF[��[4���#�X�ݫ�Z�:��k>1����V�~Xd!Ϝ!8��&Q`T*7�s*�T'����a8�N[:AնxU�-vg�R���g	1�ޠ9'��y�rW�^K�Лc��k���J�8�2���yQ*��avEp[~���o��Lyh��2�N+��]��SO>��1���ʹ"/m�N:��N��u���o���z#������&<�|⫞�5��a6���i���cPkPF�[�0l;��e�2�Y���E����~߈�]���Ӱ��(2*�遨�S,v��I��������l�a�2���A4�e�6&[6�Ҵgm�1�0n��?�;�����:u�df���%N��<6��5����AZe�������wڐ�E5��c*�����Yfª8*6�{�:n"#e�3FD���15�f��K���Ղm
�TM}������B���H%Ū�;N��xm�>V�q<�Ib��f�v=2~z��~��j�H{��^s��7�ڊ�������]uH͇�{vY��ӴE^Y<Ł�=�Rۜ ��+�� �5n�7z�7F��l�1�]z�7?������O#�/N��q[��'��s3��&��1���t�)�GFF�����(ӂɏQǣ�l����:r���L;��^s��6yٖ�ڎ���sh��������>Y��Q��m�o��T(l�m�{��]�2�,�a�ෞ�e���J`K�cID7
׍!P뇬��\ެ�N����j��/��y�5p4��>�v=��΁0GE�c�v�1-�@����۳���(�e��ݨ�{�r�Ƌ<�۴׉;0��]��H!��M{6	,����
�A�ӑ����y�в!�R�y
����:'�`k�0e�qVN�6��z8���1���9�C�
a](d�Q�Lo�V*9��08p$3Q��4����<~�i��R���*Q���M�ԫ�O�;�����l+�E��0����5>-q�����.��h�.;�`��`e�ژ[�\�VU�{��S��R�����G$�v�ܝ2�IAy��R/Q���Y�y����e�yU�8�E�De��jmE�&F.\��ڱ���pb'O|�뼉v��7�9���Z��z��[��$�a	�p���K+�Ӯs����p�������P�_O��/�ܗ�A�]Z��E��TIt6�l��l��LhU������������p㭉������yÝ�M%6��TF����ub�H��z�H5w6Kܜx8�z������,����A}�=�LEU*�j��6�9M�"�?���akǕ.�&��}l(�APhR/�G�bA��iȿR�'�=��I�=���UQ�$�A⼍A�!��x�^�F�+ejgkg��D�gH&?�K�O��(*Ih��>?�_���PY�V��o�� N]lɬ��aȵ���R��<d��L�� ������FיS֘`�8>��e
m����2��^�~�}y�u�oh�,�01��L�Q*����ג��S?�bŘC��f�cJ�0���Iq�d�m�R�F��ވ�e���(�����"�%?m���]B�(G :�	�4��g�-O�R?�%B�� �hC�7��,�l҈=F���ұ@�G�
�#0a�g�̚󹙔�����	i�0�6"��X��ux��������ƈ�2F��U=1�R��O]v̧Y�P�;�?�A�d]b5مN&��{;��NN6Es+K�PVd�V��m�_��=�}�T	ҁ\+`�� b6�z����� .'��  T?+=�g�������r)
�a&eD�j��`q�C��D���qX��+�Y`�e�XD8F�O�"-��wl�~Z�6D�2�E��&/�̈́P���N�ya��!6f:�(��Ї�7̒�`H(*�f�XBw- �d�� L�ejc%���b��/%<^�E�����KT��M7vRi96�P����ׂ�����%�ʴ��R�t
�R�qP.�F�؇�7�y&e�GT4�� JF �G�����`����+��,X4~�]���l�͗0M��K�h�&�v��)�����x��L*��>X4C�
;)�^#r�<_���o?��h`�� AVȊZ�#VH����5h"����w"�G�χK�]�Akʒ�p�y,F|�T,f�>��1���+zP�D�C�d��"�L� ���L���X;,ZB_�"�!�m���3��I��2�tA��D�
0�V�b��9EԄA25GQ8sɄ�BJG�� ��e�?�)�J�]�����X"�J��|QF-��.�j���0D$�S>/�
>�7d!Գ(U�l,�0�J�r@��<bšDgRt3�����q�r�M�F�T����[�S��V��;�&%n���6���Ĉ���G��^4yc�Ԉ��6�$���(�6-�\H'�p��P�
�MWēMUb ����WFT$��m=m6>D_/䟞(%���D�Hq9C�|%>#э�rMj��P�91�y���#���{C�Ew
c��"�_���ޘ��|���3R8E�(�.�Cs:\_�|Yej��cXcG
3�5�Dk��^djq����;�R%��0�ݑ(�"!��9��P���'�D�C��W�/�J_��{$�(9���,�G$,�l&�	W?T�b�sX��
y�9e�B�
�iQB��}�ܲ��`��1��Q}O��8�|���(�0�c�F��(W��:5�Zdَbq��WT�v�T}�g��}@/*`G�՛Ĳ4ʊ��Uiu�;p��5C�e��D�	X�����	&��(9��f��p�^�H+�X�HqAc��J��4��v��H�[�8�1��>�d�����G�m�,�S�u'�>b�����BP�q}�R�5SDф�|V���x�.j�#6�M-�#q�Í��F��5�U�]�+�M�/L&(1g�������������X�bs.L)	����(�b7�[�2��B�ն�;��w�S$�Ѱ��~�h�T�,��<�Ta�_�
�{SX����8 n~����7#�,d(�4�h�4ŬS;
[�����xN3���"�E��j�ǉ�9�a��8Ƹn�(pvf��7�T�b���Q�Y�ld)U�PրUi�Y���bd�1��8���x��q�k(=A�%W�.N�9@鸇��6��6�H�~"1_�=\���&�и6a@y��3�\l��&��GyT%42��`�q0ڢ!�`]�b�ITi��xp�0O%�n��[X��Ӵ�G8m�1��q��NciKqb����	c\#VR���@�66��g�����O�� ea�D�(d��q�dL�K�&����/>���b�6s��J�T��UWe #��w�*�v�4d�4e%4N�F��L	���XU뺎��*:1�� g���i�h�9Hy��sfQ��$`�cS��aJ<@�a�邖���%bK�h�ڃ5��5��X�-�s�����#�g�Y�0aq7�{&0 I6N�8�bļ�,Y �f�E�B৞�z�Q��t�OJ�Mg�Ao`����Y��<�ê� ���������Ar��^��!�� ��'mJ����2q���sT�2�@��K����(�-��9�	,,�D��4k�:�<�2�4��I��< �: 8sr���T3�;�c����fnQ���i�[}�e����"B�j���w�b��mJ,V=;�&{�Z�Mִ�@F8�R=�aċ��J�.S�]y~�6f�i������W'7��)S�O��DQ���m�PDQ���xd;���xK��d��A?�d�����+N$J_�(Fù���P��fã;�!q!'��������H�O�Kވ��"T=�JL����
|_&p+�'+,�����aQY��?��3���+�e��,X���O4�ﻶ8�&:�h�$��W�'ɤ���9�M�ޫ�rh�e�c�H��H$�XIq�b#��0qYQo LS+ ߫0����+�H�Xs'^�����e�\Wi9��i���I�E���$M��	8�T�8���F��� �jHWg��Qۜ�C���"��:�ق�Ļ�(mz���ɅŐ%J9��L��e+/0�ϊ<b����	�X(s�1R�g���$FICX1���@�c��,�W���=}T(��*�F�
��,o��� �j�)�0��1�ɫiժ�|BJb� �������R���7�o��Z{� �IT���$�u!6I���Sy�^[��A4��K��1qx�:�9C/K��	ϟbQ�fh�LY�2_�.��:�N���(�#�f�N3����>�Hq�!Kt�(gieSG*C�ę���@,�b�����,�"�&�cK��F����UQe��㇅�Jj-���;�#�Y����W(�1A�9*ȸ)����;h(J�uR��X_�q����wS;�D�h$!oڀs*`�XW�5����l����O��sur&���Rm4�{��,�||��2hwQ��x>X�j��!�'�A��J�T*�y&�
�_�bT�c6�� J��1�'Fb�Xm�#*� /@�����4C^,�x9,V:�[%yRBA��X����	��Z�,k�a�5r�a����]1a���ڌ�tl'A<���iPܘ��}��t"Oղi0.(���q���!$y�E&�
s7q剗��P�]��\�N�_�����N��>d��C�X�*���� �o��&�Ԭ=���YN�<v�I"ǋ�:ZL.�j7j��m1�P��7S�6�S���r9��g&d���Krt�z�-`B>M��i����/1q�
��f��9֮s�Q�aa��FcP�L�����s<ǩ"&�&]�V�C�R3i��Aui�w��$��_�TYl�G�%L��c�e�N�)����}�,> �)��0��z!RO��56QbF�V@��i�1'OE֜ײ������s���ryuX��]_��ꄋ���^���*�;�l۲��>E=QAN[��XD �v����(�ǒ9��9��N	H�CQJ��<���F���	Ew	"�1aDl��R���Y�xc#�Zz�.�]L�Y����{2W�dR��fѐ�c������k�#�ֳh�W��Úc��G��D�&쨋��h=ǈt��j��)��Yc��'ކYa��~����L�U���@S��.3G���8iz%��o�	Wx+QM�O�9��Ma�s! }"�P���	#�,[��\
�T��"�Ֆ���32$Fo����x7S:��f"B#��b���u��>�F�:EA�0 ��u� )����(����U�_N�oX�QJ+��j=d��#��ۈ*�ߘ��U51��ŏ���2J�K�������ʬj��M�I�\�I���F .���zVEW��H]�H�F1��]��j�Ni��u�GM!�
b�/	T�U棸J,
ewF�x/Ԡg�pr�MQ�~���§��8u�W>�H=h(1I�B2��b�a�U�C!���0�8��L��= L=��5��&J�5��G	�N���t�ر������2���c
�K��]�K%)����^���rRH.S�bI��aE�"��Dj�L|�����Ig�ћ$M"V�6��� 55Ľ�Xob<B���3�1�B�u��g�5R�	_j��G#3���&!*xK��c�J4�h����$�@�{_��u���RJD�<�OLlDԌAR�K�B��j#"Smr�)4~.�HGx�i�@L�d�k�i����e����hXE�Òg�@#��"3�֐�`���¶N۰5��z�T>73�HF�s$�������J94����������a�a�cWU�� CgV�-�G�hK����6�c��9'��ǖ�M𼂫h�7�Ok�(C�.�M�Ex�r�)`��TF�4D!A���Ñ2UVL���%�BHEmC�)�J$vMPǰ���ݫج��vA`�á"- Ԃ�fɡV��u�-Pe>�B�x�n.�xf��@e�+(P�;��fJ`"B*��RJ���R�l�&z���@����:J�]�~}E4��E�w��|&U�-��s�Ɏ96D۬�$6��]�la�n��%2U��V��g�d��H��,Ca.BC��f�'p���@R��Vk5�]^ac�K�/�7��4C��" �%b�R1QD.��&���r=��|�8#�l��gR>[sE�Fl���:�9��G�ceu�C�� b-zH�*F���'��6	�3��6��uٮ���H>����QO����OB�tq�H@>��T|�]b�=��Q�[��K	�R���~C�Vt�0)3I�Y���ua+.c4�9��G��H/�Dt$�*��<�5	?�!bn���5��'�X�0�cC�������_]��U]JB��Pu*��'�~�ծ�C���C%*2���i�s�CQ�Ė��W of
KV-Q\-����g��p��@��P5�ee��بD#h`*c��K��Td�P"I<��b��\���馩ce(���U��YA��6�Y�9Y������r�� ��^�\�@�rI�c]Х�����t���|��m�i�	�75�GV<"�m��)R#3�K�xQw�;�-��������L�Hsg̢:9�3R�R�����ry�"��T;��p'^NW)���i�c�!{���w��uk������U��Ux�r�i�P7��c�)��ԙs9)�x��ixs��>�r�5��|�,���bţ0�Pn.[ ��VA
e�Y�dޥ��\�t�]\�N&+DЖM���NTJdY���Di�ζv���g�à��6�_ˇ���*���`�*�%�I�����ja�	cc�.I�x�b�Lg|?z�e�'�7P
������Y9{�fP��3�|ǟ��/�P��)���R�r�H��}팝��K3�6+ǚŮ���]������3�U�pTS�\*נx����R.��b�`�S:;��,xa8|��^@պ'Չ�s�Z�*��(�L�" �2b�gsm�;��5R���4���V���LA���v*R.D晋Ʈ4P*Q���JuO�7��2�<g�#�B*b��զ&��h=�����% `�o�#́�/jh.��57<G�y�L~o��3��3OڃY:@�W=A5�sYތH�Oc�&��A����e�Sɢ�5͞Ӭ��i��i4��#�u��D��5��L�u��a�`������6�������I�:�;�8T��y��������=��C]S
⓱b��������S-ɯ�T��ďA�j�ژ�Qq-�S̩�}�N>VS��w����+��)�E�P�Z�klvQҌ��U���T(�,>P�J�b�O@%v�hM�F��<
m�=����]��󎦽:��������Oh�L�����f*�]s�3��&N���g�C���V3[�@�4�4E�_�5����7���1�{��Ī�ۦS�u�����wҒ����;�F�z����^�ǖ,�߬�:+�(�]G@�Jo{�|�6�[�R���2�˫=��s���A����6��޵�n4�};Z��rzt�2ZSdn6c��F:�s�Ϗ>H��:�FE#Cw?��E^A��b�*9�/eM���;�=�@��	c>�2��$�2LV���cy�tC˱� wb�O5!Y�ev�V��%ϧ.6W�t,q���{�dyfO�z����TH���נR��U����B�$z�L��^��v���o{����_,"�0��2��3��ϡ}�a�Δ��Υ��w.�{�誟�KSXtt�N�s�NL5W�m>辍n[���0K�t�>�h�;�q��4�Ŝ飴]t�r���%T��m;��>w�,�ޟK'��?���h{�]�ɺ��}�mM�DԢ��K��C�jLS�X�o��u1�sR��xuCխ�ݩ��P����Þ����O=K�f�@eF
��TDَ<�q�+��_�N�6�˶���n�1+��n�~��(CCk_�?s<��D��@O/]EUՍ?L;���^T��*Ma֎�co�=EG��m������S[@�ٓ���K�����N#�+g|���O'��jƌ<�Ȁf���`G�&�Ǘ�x��.Ru���}���鵥���DN�j��D�ͫ�D�|��5�)�1���'&�%��8Nb��T�e6��gd�c�Cec'�J��.E�L�WV��j��rJU�>�߼�������މ���V��T���Ot�^�U+ג��A��p31�����=����)8��t��t����>���|���_)�wSG[��Ţg]A/��Y*t�(Up������Bއ����Rɤ���G��ȓ�ߖ�~�`���=w������~�`0my�ӦvRƝFC3�r]�T+�N:R�q��p;���g�a���.��t��С{̡�|��W6�7����>�gr;w��U@�6[=�H$Ш�P�D_Z^e���h����H<��M���T���c&c�-rT_��,>}#���K'���t���oK����CV�2)��E�jm�X"��&�,��;�?��~������_!�}Gr]��̻aV�	�urbjZ�n��g��wn5h�C���}|;�cv�~��g�}j�fg���:���O� /��"Ųf��X`���=g������&������W���<��{������˾y
=�2s�_<NO=��ܮn��Y9�E��{eo?��S%9{���K˗	G�u�)R��ηK��g_x���v&��L�
�$�}�e�R�*	��;Q�vC�j�nc�4GUhA����C<�JG�y�$�ꬿ1�Jƍ���Nk�B��O��=_��6Ņ�*��zY�ɰY����>�	H������}����NL�_�yz�Q�Ko���A��LA�TI�R��葕颊��H�m����u}�����L�;�$č�zm�z�dQ�Γ_���ZCKW������f�B\b��������VV�}�ܛh���л�K��>��g���C=���)}}��Nz�C�C},��R��M�*���YJg34X,��`�:��"+�[gp�	�(�E�P�W�!�C�FO��=�Di�����,�H�(���[_i�[@���]�3R���VO�
�%��03���̲1i�tɝ:�V+���W�>���nt����1�?�[j�兒�5Xe��k�f��YNէ뮿��z�I4�Z��2)F��*��7�G~��t�G����ffS-T�.L�[W&�Jp���8)�'�*�*�f3a9y���ӭ�Wҭ����oٖ.:k�y��韮�9��uLgQӖ�� �M݆*}EVZۉi�V�؄-I�:9<�+�XgE<�fn���W��Т[��ſj8B$k�u�*cH삂��m)���@"k,e������g!,��_<a*�'��)��&"nqKN��e%U1���z�CA�ewz:���􁃷�SNؙ~��+R�=9�٬@�C��U�y����֮RT��>�@��˯��5��5D{�-��c��S{�@��O�7{6E�L9�(Y)��&��,[E�j/�Cm�5[(��@Zߚ54���?��O=F=����N�V3Kx�W��mK��so�颧�(W���#=PD�ݿ{�RLxq�� /W���1��L$�C>����pB1�"��L����R�0��4
.j�b��0b�{A���oF�['�W"8�並�*�@$�t2L �����L�G�Iz�C��R���H����|�?[����˶��7<E�|��t�GХW�GS�fP=����Ot�ns�c����DԻf�,����=w1��'�0�X�L�MW��t������s��ޗ�^�mfmO;��AW^�$�i�R>}3�d�Q-����T��9�O���Y;����h�w��I䱂�ڒ?S�����hG�W��˄m�ѿ�F��mK��z˜����>Ms�sz�M�����WXL�ie����X� bf��0'AV�ҋ�fPcˌ���d$Y=*4���*a�t<%��a��.�k)�16s5�6ݏ�S����$)EGU��zN�i� ѫ��t2�~z
=����f��LTO�iy碷�n��l.�؆�eJ�w�@�����
�|�4�f�c[*��'���_��=�2��N�ryz�%t��K���^:�sD4�ġ��Ѳ���A��
���Y})��ζ.�f���f���c��N9r�cޮ��S�_K�_��D����,�"Χ�^r}����C����'�f�r��k��w>Jv���c�;OO� Zœ�����S�4"�ď�RcV����ƪ4�I&���^(d�ш�*���!�	����F�%E	�3�S����.��`
T�M��s�J6���`��ѓ���w/b{{;�U�6���x�T������28eZ7[Lrn���֣~���L������`����g��B��V�C�C����=�)���W�be�����P��K��U�εI���`���^���>��{�k�j�nz`�tσ��D��NQ�Q��]X5�K��k��ϟ��n7���*��<�X2 �e����^��K^�+���ɢ�g_�;R ��JRyQx�(��.����+�N2O�hbH��e������p�&����g�~A�L���� �����S�PQWVP���uH�j�/	�>@	Hf��w���Q�!h�Fqp�P��FTc�5t;�$!��i�WA
CPS����)TD�8+���`_ޜ���b�L��,6��J	'B�ӻ����_���i;�[G���HY�q2�C�mn�#P��$�XJO�#��k,G>����p�Ä���!��ܬ�d �{K��b�l��3V����4x(�b�O���aB��Gg�t����@��q�p��o�v/�k"�
�S���ME9�5/}_`.���B��À	�C�'9]"�,S����P�[ .*�,-m
���*�WbK()m���A�=�m�+b�s��B`{��Ҩ�㤔R͛�+�F�g?	3�����������
Ѻ��<�X�%��B(=���ʉba�l�j�l]��a����*.p�=c���Y�'&VR�-䚘�n�
,���_�V�RA�H}2�GUAccI Nc!��U��G�e��J@��7�AJ?M�O�@���T=T�A��T
EN|i!)�Qc��P7(.����Cĕ)�{2�Ȗ������n��Mq/��#�%a��s1���"���b��(�^�RU��������� ��!PB�-��,Sk�MJ��!�rb�5' ��p�T�J����Zj����G�A[���yҗ�?���QT�ut5�WY|�'�<��/�k;��0�y1@��U�S���wL��NDo9a[�п��yA�@��*a9�eE�/R��Q����X�6�t"g�)Ś���V��/�`��'R�l$ʲI�Y^ &D�!@8 Ѡ{uʲ�$ռX
Jy���l��5\�y���8�R@N��8�9(Ub��3�V����0��t�s�
��d�mR����8�XԘn�P��V��51E�Y�x�� ��͵���<�����T
]Ή��pe]��]pٔ�P�֕ �X<�K���<���(
�b���yUI�����C� 5��U���	`�+tba��	��v�R�+��,��eQ���	��h��I��@�����ErA�<�j��rA<ӑT��-&$p+�l�.��M: �D.��1� ���LmF�C���!��݉�`���	��@8�ͬޯ�s�r��t@2T��@O��a�5 �
O�*�T����e3қb�R~X1��@2oul��\>��t#I�,y�A��٬bV�PJ���׵�(��6{FG�8Y9ˣ�W�P��*�_���f҂R
�jC�h� ����8�N�ιT���IʋfI�;X�S`�Pz�E�{��L&(xUQ|%��*W� !@�\p� �w6!�)����s1,0�[&B�yl+�,����Tx��[$Y�!0���y}͛
L)����!g�n������,:@U�O�*}+�//�bsHǄ��e̛��k�G���*��<Wg:M�>�� R����gB˸!�X'q��4��%�mTS�@w|B�^�s]�H}Op|��v�ڶ��(�Tc=��=��1J��1���U#��+7^I�Dk���$`(]@C��A$�
�w4��mw��Ա��T\�Q�*$������釩��Ս�0�+T�.��U�V�-�l!̢]�؎��4Q! .^�s��O�-�5��x?��TH�*u�G���z�#s�&;�N����̳V�����]�C/>��'���ST�~K圲|ϰ�8F5u}��#p�}h��?C%t(w��D�c"��x���??I�������v�K���!uN��5P��/���?w!��n�i�������A�o���@���g~��e�����(�0XT��-�4��L&G�����IauP���l�y�!�A�'�v�9��y���
��{���B��N�QřT�'�レW������_,�c����\CJ&�L�Pl��#^�iوf�;�v�1�Y�R��k��9�)���Eǭ��AO,롔W!�S��<s�|�u���\L��wo:e���5m�A�ʞ�,��3Xl�T�n��b���s��l���e��0���Ru�������fNTa�H�/b��h�DA.27~�5t�od�X�����'}�bS�3"~�'��1�5�E��\���6D�n,09'@[&պ
� �D4��giv;��� �Ѽ�	�w�芹�O!��Q[.m�������󑥓yP#�9�\�)Lp]i���*���7|D)E�;�i�	������+�E��iR��Y�E
���H~2���x���# i*�ZET{����M{��Ւ������b���b��כ��� n���q!��q�c�YA.�/�k���^#�Q#ҡt�cBj��F���*K��|�����pC�Ft���kؔ�H꧅��}��iC�e�uO��@�fٌ�E�2��{6��rq���4���3a��|���AJB�p �ԅ�&f�_3���&I���9�p�C�ur"#V�Z�� rB���$B�H�M�	���TX������%׍'u�F=P�bCu0lG5�&�R�R�M�+����q��|�8Pu� f��bԓ����F!:D��y�9N�)����
U44�k���5���yD��bh��-�_��÷�z��Q���~ �lE�ե�)C&�H7��m 6���cH G��(�v��L���-~~P$��R�����n�@��sǺ�f$VNzv�=���4t���2Y�W ��#
!kZ�����bV��L�)1W�r�4BK����gJ��##����瘽{��=� _��-���T�3y$���`H?�x�j]�d�\Z���J<��T�*�L�_I���t.��1p�2��=ߴ.�y����etKJ���{�:�M�Yʁ��߈Ԏ	<ޤf&�� l�*���}�ڵ�7����F��]�d@6By��,�8#�k8�$0��,�\I�'�(p�pU�$����K�Z�|���Hm8E)J�d�Rg�@�#I@B<:���T�"!vd���ä��@�Ռ���
C����J ��b*M�:��T�@E��GWrz-d��򘉠�x�̭`���)I 5?���Q�IٮqA��[8�Ⰱw�y'-^t�,8F6�j�~��E����˧�$�9m]$o��p�.^�.���
���:f ��iB�C�It���ZU�P`�H�_��T𹧞x�.|�/��N�J��}dQxA+v�WgQ�1�\ fE� .��"�^��sK�H�ܼ��H&rTsa$U�	�b
��z��]Ya1���Ɛ1\�UED#���(�?��ZJ�C��tEUX>lt�d��M��\P³&Y�9o�����5��%�!<�._Nk�RcS���q�r͆	
�){���]��c7Q�g��Q����^~��[Ջ��\%��~�4.��F,7|��R!2��¢�� �4ܲe�؊,�e��9� �NA�����i�+�C�T�PA�j|(�lGC�����ء����]R0=f��w��(��দ����a��Ǥ�[�,��T�$�Wzı���֧�s(�h�ƕ{`�c�ch}e�S���/7���C÷�:�&i!jd#`%�I}��l"�憱�!l|����7��-uC��b�I)�O)g���M��i�?��u95�>r�x��-�v7gش���t�q�aȦ&!p)0N� 7 ��=G7߷f8�~�ah�/8�'�8���~U��P}\��bC��J`Ѫ�}t��h]
i��n�f6,�&|�F�HQ2�lwY�jU60�\uBI���.RM[�H��}�D̤R���e��ͷO^�̵f�1��IZ����{:�3Ho�с>(���@�MD�noXA��'=�M�8<GC+¢�e�&�,4�Q��U,�()����d�|H��@�tD�F&Y�h���EJƽ./)nR)P��zS:Gi���T���b���+�F�
$��G%"{�j5N�p�X�G�ԼF^/f�����hː,r�g$'�AZ�l���=4T_5�u'�l���9�b%�ћ,�cP��O��zC)��q��M�Xx-�H��b��*�I\+�8,5��~*��V�VR�]B�Y�YI4�~����'8ҏ�DY�.����DJ���N=���L��Xz$l]m*563�UJ���aqE��d��6�q�Z��78�*����5�&�����Ł�:�(D��'�o�������:����A(�X��$��֩���br;�5G��i�u�HS�DFb�V�+)�I!�ULE\|r�tbQ�j�XR�Η�R��A���]R����|n�\�kl�jQ� wx�MK��_���F�"��Hİ�qZ�L]K'V�U~���|�:���0��Oƨ�����olA��S�E�tm��X�%f2D�IM�XNw�X���0�D�$AB�����7)
&iAb͑٤�5�X�r�H�q�J�׎�EL#=.ɻj��O<��-BE�5�'�
bڊ�%��F����b��0�M��#H8���/z2�eS�8N乮5ּß3�T��M;���Z8ĉ&@�@b�(����Nn�7^b=ڿ�|�GҬ���$��\�x	Qp������Es&���Yqn�|�5"�r�?#J��@�,�z[��@�Z
*a(΀^1D|F{mEq�_ƺy!� Z�|����4�Q��x��{��ـ��3}M�\�ډ���xƖԝ�8@�eDB�]�E��<)&�>�&�$Wץt:K�(%#���$nr��f?�'M����:�ǆ�a�s���~�+�r��ZO&�����M����D4��������f�~mD�%lisyx>�k8I�ў�X1��F��9#)�/(�f#"�ՒI��A��-5��X��5���ؔ��:I��Γ�=*b8!۳��L����bSߔX�/��0󖕇|�~뇆����8(3W~*�qC�S������3����[h��o�nh�=)��?D_}�K�S��Bۡ2���+V�A�5���[��W.ن����UOc �3���W �4��j������ت�$��_mW���'($g�hY��y�9��o"t����R,�u5m���l��wI��ύ�(��I�l)t�����I�H��:�ee�����q��rP$y5���>��8C!�%�,�7ְ�8P��Ke�cO���/^F�G�Uy���"�,�f�T���}������]��Im!I�������G�%UC�Ԙ �� �y1~��o�k��{2kub&�����Z�i��ZV��q.}���yC��	tP�L��� ذ�.ʼ���~�a����ӨR.�:&�~U�8W��+#e��������c`�D�2�Q�X���^we���G��:���t>h6^"�����3im� �ӷ/��D~����R;Rj�1a�wHFv��M��CC�(P��q��d��j&�Y*JP-A��A2U�����Te"�{��l�[ �:R�q�LS��-rR����s(䲴��QP#_��
^�z/�S
4��ç^�fT�&C�
b�/�@��K锋lR�yS�  �Ђ
���󔚳-}���h�\�t�cD�+�ӓ0�}O�@��8ڼq�.�o(�d�am����>�)ʙ��³	�#P�}�Ȧ]�Y�:����ԙ�P S@�i��zdk����#���qX%�+�@R����X��)}D�TֽPp��ՙ}cC0$�� �a�^�veG*�!kCu���Q�>M���-1� bº�<٬
�#��Uw�$�\E 4\�m�.p����!�P�sF2S�l��<�"��Yǔ؋�Ĉ���r֘;����$5Da�tB%j��d��=�|���I-H��*�-�n�z[D�� �Y���C�ֆE&�Z�����5�Ni��@�!pB�ZC74�z'	ϛ�*��V�T\��>�S
3�UA���
��)���Y� �am:���E6�Do�q�8l ,�i�]��a��, �ZI-	K�X��Ѵ]�y��{�U?�5�c�*/�a��Î��c	9�ir�4���(#�<�J�R���YY&B�9+�U�k�G��7�j(�r�(џ�������6�"T��+��"E��G�H����%�2HE$�7�xk���6`"o�0�[#ͺ9���2y)��0t��ʴ�Z�x����](�	������e)�e�Hl�Ʈ '��,VA
��Ϙɦ��pr �N��&�j| IP|� �C����AҸ�HR�IԵ�@��㴊^�VH��H� 3pS�/�X��r��{rr$����h�R~/a��H����\L[~5T:�'�A�JAL�ؒ�&X]Et�W���`��A;ɿ1�x� �Κi`�jŊ���{�[�U��
;�*Wu��PMGRC+ �(�p�>�
"���lT�\L�- ���%�D��n�s���\'���s��ϩSU�T5��}��+v�s�^{�9�s��? 6P���{������j4e
�� Gd��zm��tݼn�t���[@�.i)q6�0R��ܥ���	�Mم#m"�@�:+^C�xl����2!�����ma̜����J�,`,GS"��5� �\l����u��! W�\B�0�e�}"�p$���1HR�E�a�vN������H��S�o�R�A�K���d��bcЛ!��������إ�d����5,e=٫m��z\�ְ^_%��5�l-\���We�#|����O��2añz�\�
�S��p���VD��J�b;���v�u1�F5�,���J>�wi�BS�f�X��!���u�^(�U��He!�q�\�\����b�¡�߹J�m�AD����H�n4����v�Fq]��~o���6F��P�����������gMT~��螰{=�v>H{i�����{䋍��)<��/�6�d.�OCTkl�0�����g��U��}��U�Zް׌l`e����'�"��ᨅ�v�x�-\�l����#+�	����Ae���ρ�!�(Ҧ�����p���H桫;�R�nӊv��d�<�����L���+���%�XT����%?��=J�=+�<�K���I�F'�k/+�v�U��9��6?��}�Zg�*��[Q`�La�XeA;`O/V���U�;*yttȩ�q�/]!��U�"���tG��/Z ��@&BW�3��|9���Q�B_�F�-��X�Ќid�������2,O�.�!w�K�A�X]bd�Kaf#�ʀR��!�B*цQ6��q��ܴ0 t��U�A�:A�� �fcQX4�����)pH6Q���Y���y�]��i��.Ϣ��f* �nL-�v�%�]��ZMVJ����T�����l�,.LmC�,�'wQI��FS��_�8c��^Vny�Y�RL�GDAe�i5�5�W����p�0ϲ�<)̂���`��et��� 4J�><�1,	�6��)Ѐ��+>0s,���B�Y�m:AQuq��w��yV�oҎ�»i��*�`�vE0��'�ob�@����+-����"��L����H:F�_�"��mjC��\�{[�	��s=j�LG�!�BZx�z��8IՅ����.���Պ�]T��Ŭ9�ՙ��υ�}&����j��)�s��	(��UXw ��yMթ���؁μ�,i��PP���16���Za��U���X��������+���M]����(�o�pK�z_8�Z(åp�8<2��ƁұN4'{�_��)��ܒ��z��͒.�B��#S-I}��al��|�ν�

�͊��/8_�H[��.��>�,qU,��k7�3�Z��k�l�؄2�`H[�B��,k��y��T5AE@_'���I��m����	5zi��Н�Y1��3#
���<��f�F�}�;��L�����8�ź
8��C�ݑ��pz�b'���Zp���3o���[���1*����<F����-\f�}/�@εF%�Mb#� uc��}X��ݷ
�.D`5!�������G�\~�:��8�q���P�h�k5�.t�[>4��Ѣ��otR�s�	P��깎� {1���s_�,1NRY�s�ե�8���u� 3��֪����.SF���zt=�%*"v��PP�{�Ư(��5qWݼs$a�,集
,�P!��K�ّlKo����4��Y�gӧ�Wg���K����T>�3~|R~�ޫ��0�Q��XN ��˂�Gi�-97ͱ[h�U���`ߏ�j�	DY]f0>�&�XPL���\�AI�� ��|�C�|�v�Y .T�{�����[��Z�w���pж������5p��l��✹��Zs�9,r��!g|�
��7v�T�q�[H<�׀%�Giuu��PL(�TG�vY1�tn�,׶ �5w6�-1��q��~���7�n�=A���]�ɰ�%�UQL��?��ی[��������D���wcY��E7e�n�Ge��TaƲ�쮪t����:C6��J5hf�N5��@�����ӻ��j#4�5LF�wzd�w��r�Li�̭���`"�{鉱��(\ř~6T?�` ���**�V?��ĥ:�X%k q:kU�;}ͼ�Z������HS����}ZGr��!Υh�u�l�$YҬ%� �l��F�DE"���
��L.��X���@�x`�af���<�>�h����`�ff?�����A6t�^U�$
,:�e���a&x9L���bh�
��/�Ԡ��c�2���:�Y�`A�9��/��$a��硆l#n�2*�r��瞑ZX Q��QW�Y>�<�`�A�nQ�UH=Gܥ#��Q3bx�:��I���*�D��պL�����D���P�N�-��6�j�g����b\.��ws��2]�x�C�p�D�����C�G��%��pp�v^�8�yO�7��
0�la�]���!��Z��0C�x�WG�P���D�I��>��a%0��Tpa6���j:�қ���<�s/C�3��x���J�|�g�>s�΁!�C��~���}"��� u�-�)f0��`��X�1V3EH^W���Şu���ݕa��IbB��w�^�EB8��P�6ѐ��;�W�D�z��$�A72�@4Ks�z�|my�����Jn���%�����!�4!���WZ8(��iny�^�D�ZD���Yw���u����JS�� !�U"cĬ+mm�.��R	�
J
gZd��-3r
e4�4
�g�<!q���,���0�%.��dlTDd4���P����������P3�)Q�������j��������/w�F��6��?��r���b�G�%��l����`K$�I��eW�����\��7������������!�|;�>�v_���|�&.���!AA̼�l�O���%z$ϥ;L�Zv��t�V	���KQg�,�(��T
�\̾�y���~#�'�Z.[��W}6m�6�sM˻ ]
;+�@��
�}��f�9�f�G�j��1&�A���
4>�:�>�tSm�^q�B7+u��^p�mw�o��>Te�eH_5u�,^���zo�B(�bb���;����mh$�)4-�܋g�}�F�T�$*.��ۡN�W��-���,��.��Y�*v�y�\��
9��ݻ8ğ���0-����i#̓d6d�YS��Q�Q��w�43T��<-�{V�x���"DY�����OGd�q�0`�42���������Q4����ް��~������ŉU�m� ��pWDJ�ߎ٪��\U� 5:&�����T�a&i�Ҙ
/��̶���z�E�����~b4��/�E�Wg�R)_�ٛ+���5�C�7�ό�شc
�c&C�����Ǚ�6�s�U�E���2�-���aT��k(GU����'��T��F�`�o|��ȿ�Ux$3\�9&J劓����>�pn�]�	ga�1D ���9��N,��	>�8��HW��*�}�,�|�`��W�m�O�Xl��3 �bע��}�f�r���+�0�@��͊,L����{r�K2�K ��c���i1";�i����-/C�N�ZB���-9�d]Qrj�2�9N�&�H��̊���=�ϵ�4W��X+�G���0%�ݨO�{�n�v��6��#�in��$��5(
�?r���쇻H���E���1T>���Ԙ,�����6�g]!��}t������|O���Υ,�!��xJ-@5�"�*ɮ�z�+���'�S0ږ�΁½$��՛.f�3���"{C��I�B�}�>�X��ϋ��`h�ܣ��E�
�/h0�р��QXÒ,��K_�2[�>h�7�Uq�D[���l4�:�Z���ܠ�!F(�B����=����7��n��;�F����zzSvZ����fw���M���0L�T���Ȫ�#K���j�3��f��v��ڝ��wYp�G

6��c	� ��7d����^WR��2�hN͡GHC�����E0,��ʼ�US��(������5F�סU��R�)�
�X���*e�(_N�b�0f4.�>���Tm�HIIe���Нi^��M��&[���ɟך��~�\��w�Ei-��i��k���Sb�,n�<���F�sT���w��-�$�f1��s��4 �tM�Rr��b$uW����*��|��iw-���.�Ϋ�
��&��:53'�`�p2u�%#�!������ה��P���ke`�Kj�2��n����a�C��,�%�J
p�!u�W��P�$tY[U �Hw>^�cÓ������0�B�M�o�>	.�1��ݾO��!`� �1L�P�0\ڨ��r��ah�AUl"�ϒj�v�u1ִ��`=G/Z��f�����0�0��K�Q#�Q�ѓ�C��@��}:�=b��	�Y��\f+�Wt:��0�PC4좑�P4�p�Tu����,��@p͚�ϑ���a��r�n�|j�Vj^�>�X]0��T�;	]��ik����;�:�p9�xB�qu��C�'�Da�պ�0FCw�裨�������	��x%6B��ev Z�뿎Żn�x	��>tn��y��X諺U�0��ynGq����ð�I1��;o�[���Z��j�Lե�s,�9}|�C�ð�F��*�{�s�Q�j���7X������׿���[s<[<�w�󝘒3T�?�Y6�Q��� W���݊~�t��#?����)���(\8��' �b�Z���s�v�DMͤ>��3�)�q�h�5�F]��p�5�B[dՄ�zwӒ�#c�ӊqt_KTv�O��v��ۀ� 6��\O����-c<�5aF�GVm
�[�c4b�E_��W��K�ߊ>P�G��=���W�0�5��nY���Pc�I�d�k�{�]s�w5��[���'?����"��������ǩ��0+��6Q�fk���5�a�qQ��%�&8��c!�o��@	N�1I'!/W��(lyc�Q�<K���^'=68H�qA�B~���0���ep�
d�Պ%ȝ!�X>��i	�Iu	��2����G����MEgD�g�A%�L���#�b('�,?�C�x\oԔ[�%o�LfM/��g�NL$�W� o����F�F-W��A����z�P�����:�CW8��'�l��ԁ��p[��ŧ��1��,7�f>W���J��J0a��i�c0_��p�9\3h`1w2��/��X��Ɛ��!�e������G�����͉�E���\�z<��;��� Y�2L����<`3��+��+]ݴ��n�s1~Vj&���BSs�D:���� ��!��"��D{Ք���+y�ۑ�H��X�4PF��A^X'��OF�$�(���9��rNj�ɲF��^���a�,L��>sJ�\%>�6���H�Pj+~�J��-\J8��s�*�d*����!{lt���$T��d,�K�����v&�n��R�Z."�Mt?X����\^&���5bEV��H��G�T/#�ˣ�O��c<��h�m�-��lsЩ,�
|
��N}��qҞ�\V��F-�v������F�%,C)�j+���tz_�s����E��=��R�j�0S�si��l�[4��eyc?���Zv�%y����l�0i�\�Y%����p�ى��^��uW&���3����m4�Se4d��j��r��\�ء����׮���������XHá��W��9��r�3b�u�7~@ꈀ��U�s�p����i��3�z-���\�F%����Hܢ�(�W�ԹID���$0ʊ�0�Ct�*6?c6�V?jq�����䮖�ԁ��y�P{�QrG儮f5O�jy�8?����劣�cC|ٟ�/��V��u��:�YK�4���p�d������B��b�����zf���>��3�׺������h�lҠ^��f�S���*Vh��C]dj���!,,�Ccj��h�kDXL�$�z��=�Z�J[	w�K��P���]��13�p�uX8�X,���+wlP��`�Z���X�xbT�:b���a�bLD �a��'�@ֶ�z��6Xոb|wĀ'�wsfN�K�b����Q�k?�#�[��[��.�$��F�k���Z��`�#�� �O��fU�b�V����O��d��M8���H��X٢���f�J�#N��B�ZeZ���μ�"T�ieVL���Q�0��=�����D��AY%cS��A��P�S�qR��5�ﰿ�ܪ�iH�=�B��3��W��/*�͋�ُ{���oV��[�0�q'6nݩU�D�ٲu;��E�sF�Q��Ë��Cp��3l�n����a�����X�N��R��q�]D�]¶3��h�u5<��޽���_�+x���e�y�h9^f[b��p�w���}����s�05C(��QmlG_��bs�Y��Z35�����>Pv"c�����������`����'5�5k���{�`��p�����?���6�U�%.�d��G�.QwX��*��X,����{�w����;о�غ�Q�u�` ڦ֘B��]|�Y$b�(~W	}ߌS�$�50��*K�h��٬e��Cr�����2�ۮ�]����ڌj��ޔ܁ͧ��FA��p�9���5�Hs��o��G����5��3�}݀Ab-�A�2����$���G�	Z+���$#-3��:VP�1��e����p��ؼ�j�ɹ��[?�]7|��kO�G��AqMOd�dh57b4*�I2J���>����<Įͳ�=�sӗ����T,C;�Y��J��pB��R�2Nr��w��'9*��u;�VU��,�b����[����_��?v1���/��s����7݂g=���W��٭h���Q�"m3�?{��>�q�>�t��s������K.C�9����7��g0���	�ic�Қ�5E��2>��A�&j��_��C{P���/an�"��~��ֿ(d�7?��8��]hGm��]���|�tӍx��~oz�_cq� j�Z�6��uo§>�y�&��A��K�?7\w5��18���\`���5��?�J}Sr|՚-9b3@1Av�`�� �W1"7l���� ��!->|׷p�Eg���y��/�Қִ:�t��E�X.��|����g?oy�[�`�E(^����شq3Z�SZ�ڜe��H=��/�?f�؉�����'cnF��Զ# ����*|��r]'2V�DO�k���o�͠ڌ�_X@�x'���g]�{��y0���w���e�k
��n���]���/�Kq������=�T��]BF�(ǵ�݋G���q�/�<���{ދl����3P��&�����2�t�B�qJc��`�D-�`���H�:6NGX�� �q��.�K���g>K������s�t�mk�c�y��/~��睳K���DTd�%w�w�Kv����ڨ0'��?�����w�̳��\�T�2^8s�8Y{�sU��`����LqcZ���b� ُ��{p��b3�G苇��g�� ���û���Ӵ%!��}"�u�%���M
�Y"m'�V�bW�$B� ��oԞbc�� �s����P�R"m{��;w�x�ەl�k����S���%�r�
�9R]"!�r4���B6w�zأ���R�h�����g?_��y����(GG[<����#��h��Zo�,��7ߌ��/ğ��r�v`������.�o�q0���t�����(���O�g9����z����V{	ƂR8LgZ�J��$b~�0zK��P�g��x��]�L�,݃�-m���5���bt�\������'�u�����u�1.����܅�/����w-�E��"]v)�Ze��{�ޡ6G/_@%l�ݚFczڪ�
�q0��p�j���ˑ��T�kR[(敫�����()z�ƬW�<q��m$�k�����eg�Ш��s�]���06��!�i�u��WkX��Y.���L��&��A4�����P������J�(B�6i[$V�	1E8�t�be��)�q��`�E���#�*c�cܒ�5�$�CZhWW�;�f��ލ����E�,uPW$�PqA���/�u�zl<m¦�(DX���%��7��s7����/x�s18�u"7�e�aϡ�\o�μ�B�$�+y�0D��-��}# >ec��?J\9��g�UD�'Y�Ѱ��[eV�(����]���n?�n�zK["?����^�R4ڄ���h��7�WA�A������mÇ�}�d]<���m��#��;�ȽL#I����\õ�f��1�qq�b�e�Ȫ'đq�S��e#
-'�&J�a˔aHvj��g:[����}�k_����0]5\�/|�x��_����y�FYO���r�x�uZַ{�yj�Fu�N�眿��G�i���_Q��T_��7�8W�����g���v�]=��>�1�3
�Z8���:������N~��eiQ^����p|�<��/~/{�+133��7!�E����q;�6o¥��_��c登��Ba'N;k#��m��v��>�ױ��a|�S�ö��������e(d�J+�I��G�����`gxnu#�	5�Ɏ�e���v��ߋ��r4E��[/����ϨF)~��/Ŗٍ����1,�J���n�NO�׾�5ر�\����]���ۍ١�nD�~fozǻ�ܼw��JK�Ȼ�� ��Ѫ�(`�A/�k���S��GqD�y9&k��"�j�H�4���+�'#L�7`�����;���/���z�4ds��֔�]�y�]������w�@��x�k_���J\s�wp���ik�p�G��FP��W�Vi.��_F�ލC��8�ZX�%p��0�v{�5�������\�uō���1فn�������ô���Qco�/�S����'��ϿQ]w�q'.<{7�K�8�� z����`��ͨ�ut�4��׿	O��_��7ށ3�:��y�D��0}�#EK��Ae��ulk�9x�
�D�j�����<�1t�X�I�d\�h��H�6@��j��im
�� ������c�;����o��ضm�x5�Om�:��--���o{3�x�p�m7�='�h��7s@�t�{��:bx��<	�偅:w]k@� 'S�ud�+?��p��eK`t�߭�1Ҹ��a_Q/&C7_AI���`��D��k�����x�{��v��~���Yt�0�f��3ӱ����Y�{!n�I\ӊh��s�c��qסEl:�t����	P�q��%�fS6���qJc��H:�Ө����,����f0�]�<Ksg��o|O;7�3�M�v�=�ᰂf��5���-"B$.�]`j�N��&�/��K�}K=��y�r�M�v���cv�,���xg����5�c��5����\]j����w{#eW&U����&"1,j lv�y�
9fq���;��$^���?y�><�<l&���{R&�O~�����3p��O��܅�hl�s-q���s=�l٩�}ڋ�	z\���Z��4F9ֲ˖�/�-���,�k�Ĩl6�O�Z^�����*GKv���3 ���WP,����@ܞ��{2�a"����1�s0
U+hLoD� ��c|Э�9�S��uO�3������7p������3���r�lFD�򤯋��"dX��޲i��,�gsl>�ǔc���3v*��2 ��X�{ϋ�*
�6�y�<߄F}�V�Ȉ��+\�^�XԒ�+%��/��������ʗ}�(?o�]����0��ϗ=k�3����_�&����6�1d�;2�sH���/���*Xw�~o���=�����(ĳ47���DUm�D���"�۷Ga��6�R6��&H�@N�K���+b����#l��F0�˄�V�T��KCT�R萄�2�U��A�I�	p�zc��5A-٧�Ȗ�$�F�7��n_d�:��~��ZQa�t�K4�������>��(�jJ�C�"����/�ǣ�0bT: �щ�\���ص+��D���*��ـ��H���I�����7��P�C����C�za)[�g]`�r2�d60E2IZj(��J� M�תW:���"�-��"5Ɔ����x��/�Q:�S�a�G5R8�@��=T�M�1%�y6BK��c�F�#�r�Qd]�,C>��>Eg��{�������6�/�}�����/���G��Ncl�4/�**�S����ˏ��WǄ7b�µBy�	@�b��exGUyXe$�L���=Z��]���I�Mrg,.Á�M�،�j����>��.
C�ue��|��#�+]��/�4x��j\��u4�R<;;�o�TQ�Q�D�<*Z󡛉��T�+���Mm�X		Gz�Xo�E�J��.��A4k#�q�5�֌l�)�S��ƍ;Ā��� ��FT�<�ZA���9����)[i$���/D����&5rZ�w���]FH��MA*�̣��Z���r�X��?F-��lT��zA�ץ��/�m��a,�P�_�M�D&m�hRt��V�����J�ԇ�X_�Z�X���b�|bG��x��P�Ȇr��9��W�`�T�f�`�Ar�C�؆UӟS��)*������u
`_�YZɽ��ĕO���y�]����k��M�[�Z�i��}����l�09�Z=2$�9wؖuQY}�Y�c閁���$\��f��5��O�d�G���Z�v�7�'�v
�?&�X��A*$�_�y�AODbńp������O��Kx��_߱(�p�Q���(�INdc�yi�W��rqn�E-o��D�[�LP1Ru�Yjb.�t������h�4yds��q��ɳ��e���Q��_w��tu���������e�P��5]�7��H��}��nwZ6�A;��Lz)���פ1��8��l�-7�X����UQ�Ia |�%#��%��[W�����w�H�g�`<�q�Rڬ�R:M���ڥ0U��3���v�$�i��d	?w�&�ɯ���'��h;�R���1��͡��.��9�q(����兯����(0q�x�=r(�99Y��T��UqS�*C4�yZ�-ٳE����!R[��[ɺ����}���B��[�Tɠ0H;x�/�,^�a��)Ɲb�.����Rɳ��A)�(�(C�Q�VQ8�l^����pUk.�X�?���\��1�s n���&�ŗK���h�t�f�,D�<��Ύ�J�a�:���@��N!J0�D-)�6�f3E�S�c�&�&���Xψ���������í�G��ޗRO��yZ����EV
ő¡~N8QT8\,��OP���8(I�u.�ٝ��3���P��CA�-1[�㮽�`��I�N4�Q(dÑ�%y�G��h]�@,���᠇��ѣG�e��*�M�L�b^�h�t`�C��nCv�?p�_J8]�I��t3���[������(nc0�x�K��)W�=��Z�'�����:�R��>�w\�s�>�3-�� ���t���Ck�9��[ŧ�������.<ː�s{��+�5�������� �p���D ��j,
�+RGD��5r�O$Z�P�d,��TwǎJ�kj?w<���f�zL�<�w־�Ȁ���نc�{����9d��0�o�:���hk;��:��b#M�30X����VÊ�V�Xa���jk��П@���1+36�����%����-�Xh����;�/�e��j<��y*����V������?O��<q��cœ��P�{����=yc��f|��+��>�7��qC�,�s��H�i<��+����~���ص�¯�ʯ�[�:���:���'xȣ��o���n>�#�UG�%qp�R��e
c+K����Dt���Rz1ˇ�'z�/�Y�Jǡ����!F�mPJl�J�`k�����}����'��]g?Y��D���*�E1�?�����{j�i12E�U�8q��5���,��*�w/�Z�`V���3��*�ܳZ2eZ��D
��]���V6�S̠��`wP���	m����n���,�XJ��p�Vh��(����Đ.;���O:9�bY�O��E�#N�"#5�*t�����^���)��F��"�F�C�5�YNG.�T� �P������J�(,�c�M�h�,�6�l~c�3ч�">��(I��,O2��������'��ۂ�X��o������0l�m����>�)�+[��8<�(Z���D�b?Zn~Z
�k�5��Ȯ+���G�o&��z"͙��h�b����C�s�u�Fb\�
����a�3��^�
���U�ᘞ��+˘��h���G"�5��f;�h��"��s6��\r�$@�h
��	ϣ����A#Y�^QE^o����Bc+�7
����|lj?7P������rI��J��1*;`dń���+\6־8\�y�[G��X��,�l�Ao��O!���`>�����6o�푙�Iv҈gG��Q�1��i�dRb(��AilҖK��D�9��P�b����gU��A��F2Pn����#6��6G�B�8� Oא�;��zD@�%=s����I�D,�sLM70/�e�X�$�"+Q����Y=�0�a-?�+�0��ī��q^Tk
�dN`krĈ�=����r������13<'C�f$��10��^K�w^ V
���=nΘ)F���.f[[1�9�ƝmY��y�|řh��ܠ�	���{8e��^X��dt՚�x�J��h�.Fk*��j
ݩ"@���x�6�T#��Ē�n���.
c"U��r�.A@�������@c2�#@#�/i<�F�yU��pc��-��Cr�1
k������\�%�v���&�=��#�h]�jx^s1�I/UK"������N��W��c.��e@�9 5X'��2P//��ɀXbЮ֓=I->��AqQE�'��իG�⣂̧�2h����&����r��즙Y1X���(j	�"(��l�dCl�{ZG"�K�	H~+�H�ʦB��
Y�D��������r<��eh��6:8(�l��G���|OE4G*Z�뢥�X�B�#l ��h�	R��H�~i�dnR��ж��V�3�%�s
�h5��SLe��ĖA�u���S������A��?1w�e;����QrBC�U��P�ͽ>�M��t^��	XD��\jm�0�C���O�ǣq�mP)�l���"e�������/�,l�[@�w��[��/NS�4 	�>
۸u���Ƭ�:i�Ա����%��IҤU[�z8g�n짶Hz�Rk8,�̉�PC-�Q$�<�����F#Nb?��U�X�{���b�ʭ���"�Qè��+a!L3�>�шvz���4Y�$0�&�2�Yi�JA8�`L�Q^��`Иn4���c��˼b�Ǣ�xlя��v:4�������-[eJ��p��()�?�aV�G9��8v;��	�L�ٕIĞ^�����t|ظ6n�����&�3#~��{x �;{������b;��g<N̪ȃm9���t&R��&M��/ޥj�,��f�^�|g��.A��NG��^�W��"��QPs|�EC�Ӛ~��q0Wk�QUW�8�G��}Ypf+C��(�]�F�-gwU<�@Y���⎒��L�	<���(2�Qs��=�%hb��#t�J�͗�raA4r�UU�WmY*���2Cz$�`��N�}��jr� �p.��Z�X�����8�b�{�����"-���$�h��!��vY���g�� \��?��!�N�[��J��� �L=�Bŀ:p��Y��?�!N:��qAA���E^����YK;����h�m6�_{Z1�^��x �ZZ��6W�2n�bw$�(�X��RO��b�k�"U�Ĵ�@���2��j�mlajX�,(��|��.\��de���%�V�P�3���9-ǤQ���%�F]V�#s��+��$��0S�D��Ȇ����,Z�`h�%-i�V�e��nte��D��-��]&�LŒ�ԵK�=��@]�x�A\���fԛ��W��gd�]���_��p�E�;e��C䨠��` �;�VE\�,��~����@��ކ�:��@�SC������	Y���p��h�� %�!`�
�)E�i�x��³(�,F�h4@�M��G��b�*�R�T���a�̆y��)%	�k�.����}+SQT��)�I�+��"r�����aE(� �b�����Y���xW5�™,�-�}�E�GM������yn��p,�b`���2uG���W��r�����8~�B#��4���ҵ�g+�" ���S�x��A�!�Hu٣IA�h�*6EC��"Ҙ�H[	y�e��scW�cQ�����+�ȃb�?��NTXp��b�G7U�4�IHEJ㙂�x�ުB�����!zWd��"^����(�m퓖ss�V��v�5h��p�H�s<�X�P�8�VܒO.�R扆��}��v�s�X�	wR���,�#^���S-��E�D�]�㸳G�Q�jq99��yD/D�!�4*.���q	߉�J���>H�5��w�r��5��hFa�I,��,6����Q8�\���q�VBd��zRdU�x�$o+p��Oȭ6�xc��:L�h�Ck"�$�S���Ƹ�H;1�SӚ�]�,�f��)dؽW3�|e܁@e�\�(5Tb1[U��bYeq��xz�Z�X�`��!�������$��8�1x$0��դ�Bn�(pVK�\�x��ʻ.�'A��6�=��1���A���Z��x���Z u�:��w�`��f0i�p��5 �K0\�^�����9P}�P��-�;$�6��*v��OML$Z=�~W�c��g�f/aK!G![�@'���{-�	�P�6U��rn��e�B_�q��	j���y���P�3����(B���#1�#CS�C��e�X#�h�t���o\��>J9Z1Ĝ|@*�6�ۊ���-֥�����Eq}�u᫟�\;o#�~g���/��̣-F%#�*8bwt��҇?n�X]fkD�Ϝע�:X�9=����]�>T�9#�N��'�e6�����E�u)�U&��8Tۤ��^-p�-�a��Of��A���"�zMÓ���u��Q�4�џ��M[d�&��C��w��ϽL<��z�i�6��Gj^���1ƪ������%�F�g_��~!ww�Es�K�z'����-���i�]Pm�П����p�Tf�k0;��v��X���,1��-��>KZ���U�Yո`ʅ�X��銊�dK^���5[H[&&��>���_Ʌ���(�R:��}��m�g�]��x�����/GO�d��d�����~
ؾ��6�'��K_{�֩,f^�8���dԣ�j���[O�U/�/^�2�6�@D29�?x&�?�g?�J۩�2��^�y�Lm�Q����_�_��'��h�7 �4q˾%��Wc����jaO�
T�G��5l\�����$��8�A!gK3��M3�X��7����G\����Qk��n�����n�\�+)Vy��5�ח<�I�͙a϶
j��~��E3U#��̆vY�KC�h����2N
�KK���}䪲#1�2����U�`{b=w��k+�B��[� ���Ɠ�������2�F��%i���u�#IG�G���B{%7�S�SF���B%yr�ꮲl@ٖs4*U+$�5e�f����T}��j��e�㗭Ze\a�Q�߿ҋ��%�EVVÛ��f`!���ES��H��9Y�,;���^����=���.������o�#���^��X��_)����7Y��2u�NhT�L�z�/D�����Ci�<3�GPZ�����ל��u���MvT�n�����ǆ�ѝ�Ul�l�dM;�f:�sW�r���5 g���Z6.�U�f�#K��]��xմz�aC����Ov ��x�2f��X�i�/�հ鍜�}a�e�{�uZU^�Ҽ!ih�8��J�G����c��	�����۞�o��o�uzX�R���Fk��+n(0�pƑih{�=HU�+��`<��f�'�2��D��7�B��T�pe�h��,�dWOq�C[��zR�86��j3���� ϗ.zY����.>B4�qBϑGG��*6F��-X�6��\���3B�[Ȉ��s��pe+���ɱ_}G�T|qn)%��I�����-������Ɖ
�FQ�wN����윂�D���V�[�����١s�=_�ڞۄ�s�;�q'(:#V���?V�1֮[-Wb����2ʨZ���{��S�6%��O���y��-7��+��WV��<�Iן�5�IL���;78�����z��qn�iP��լ��<w6�� 'c-�k�v_OC3��3K#>aS���
˝T5���G��u^��aBV _�� ���|p�dJ�C��]c�T0�^�ޙ}s2�K�Ń��3�%�h[�}U�c#!M��B��%���᛺���6��u+�(�	'~V�U��:�*7���=6��;�jh�G��;\�N9�8�}���7��0���bh�Q���|��sN�K��h�u�����l%YTKX�HT���(mP�:��+��݊@�D,a�Yq��F�y�(5�9������w�E�(Z��X��aeO��S�XAUo��uP�;�2��Lk跢���-v�l��e��&4���U%�?Y����Di���r�Qq�,+��,D��!���(�4�oB�r��_�_N�Z~?�/�)U7�I8� ͦ������̿-�<�k�"�]�ܮrH�YK�c�M�����(�)���e�Ga�Y�G�]��I�`��W� ��}�}��4�c��љ�<�w%5�Cd��4�����u���5�m�w��ǳ�����}v�z;�[ Ѭ���q�A������w�,L7�ǐk-�Ά��X��_#��l�(�� ��2���Ώ������P+�+)F}DVMA�Z?����ֻ��*4��i�NT�-�����0���,/���|��~��ZB�G�ח��$'uKqƃL�I�-�rN��1��(��(1�n�[y�z*YD,��r��s~W��Qva�"��h�M�ǲ�w{,�>���Q&����O^��m`��ziM༇�S�*'WY��_23Fc�Mkڊo��U`F��ベ���a2V1Ũ�E;�wؔ��Ga��^�v�Fd�&IZÜO�<`�Yl�A�>&[���� �7����Jo�w��+>�[�N �w�&�<L��������`�s-��U��"i~��!����A.G��,!]Y��΋�}��w11Q�V,�.�(\s".�MD�-=���m��d��jv�{(�й��]t��}'&j��-1��Pv���sx��������!O�
:d#U���b^��ui2�]������%,����2L{U��b���N�aZI�f��o:�_N�������c��ba)JQ�aMI���LU��L6��}�6pE�>����T�0ꃳ*e�����KP��;�X�T�βD�<*a�4�=�������>&����W.�^�%[��ܡ�X�#�*b�,��M���Qf��>��Z�jb���F�{U��Rg��+��=:r�d̪��i�v���}�C���
��+Ǒq� [���̝�'
����U���51���`��2.)�[%���Z�2Y�`1+��P��x k7iCd���o��zݎvw3�Ċv&�<܏G��I�;-�W<�������pYH���1Zǆ+6�0��j�JcF����:D'�jMk+r�īh�^��(o��>ܰ%��z�ݥv������Z�����Im�ͱ�
.mj^����la��\���̚��H���Jh�~���
ƭ�c���G)�f3�1��%pY ��u%�WLElMd2���Z�]����N.�/�5�c�����B�b�l��zl�[��!q�f��'�Y����c��E5d�����HG�?ʞa����i��q?j�]E[x^���X_�f�z�5��|�++����ވ�Y���':�6F�6�[E��EI�(tP[��U�D�S�:�y��n1ºz��e�~��p��K+�L���fD?�J���,�8�N�;;�Z��5|
VY��&�J<�td�
dD���ŝ8��]폰�{���9>+�u��AY�V�W�� Ř���}z~����.0'%�sS5Z��Gꪎ�q��C-2He���E+Vo0ޥ�$�U1�3Pau��XSd+&���4�R��ͬ�5tF�.�b�Vv�6	��T�KSm�]��z\�'��h���h
�E���r�[\��v�-6�&������Mc>֠�Q��EaU�
o���g؊}&�}�7��M(��GG�E���{ޕ�-��mP����y��cj'EiN������a��I3$���@1��tǛ��D��(��'2�$����d�5��U��E�^֘fV��F(N�h0�`Ҩ?R�B��,�Б�Ԙ9ʴ���i��H�LB�S�90ΨA)l6g>�vߎUl�����(�x@D����x�q��H��^}�@��|h;�g��(�[-�T�`XYs��D�xP��U�6�ar���!�O<��� w�"�r4vY���uВ3�a��ݪ��X�����;�&�|�f�1�F�q�s�?�fg��.Y,O��X�^^�X-W��o!�~��J�ɝj�������"�(��v��������]���6��*e���H��]�j��)G
���h���:�*��l��#�0NZ�)n����qF}�"��^����C�*�o5��ׄ@xOfbh@,�O�4ǘm-p%y6Af��k����4L~c��d��Ǉ�K�s�����e]�0��m�L�c�*��c��ǸgF�r&��~��F%6W���^g��k���C��/G��/j�k�5���f�M��ڮ6�Ѱ�Q��B����jL�+rx��
i�Mi���Q�.�gv��|������k0����������Ñ�� s���Y�8@-D��i�X��*J<���:BWk�,k��S��f��G�w0]I13a�]�����Y��k����i[q޹�cv�F\�5���7@�kϾλ���۱Y�%�-Z�1-�G���Pm������hh�r��r��������bBN��x��L����Iy%��Yۨ�	�j��qе�Du�S0�D1ĭ�� RN�I2��3���(��.w�Ot�H%��Ii	�6M��W�;������x�_~����ٴ˱z�^��$���V|������֕"YS���	;/}8n;��-;��Qo�����8��4A�q�iC�D�f%,r�I|j��ʚ�0\�D�7J��v��s�@�F�4��¥;���M8`Ho4*�����KbC]�1�[-5�r1�'
UƑH[�p!�X�V��\s����ѻ��q՛��z�c�
䣞���Y?�0=;��z�x����o����}���O�7~�٧�;8�8m*�-�0�b�����oEy�c�T��Dl����}Ѯ#ͯ����.()���_~��#���O�R����@�*b-%?��Ǎoz�|K`7��JW���Ko�����0�˞�r,UN�(n:��,76�a�y �A(F�ᥡxm�%$�Z����8��}�U��]��k?��wnr���թ��:��=d`�������?�?�����Y��F�L,�50Ԟ��:��&a!������]/8\��ڒb��a|卯uu �6;�|n�1�����bg��KQ�r��-2�H�bB1��kk��,��+������`�\����L�A#Ws�+���D����ȣ~�"saU'��v��tw��O��M�۵ �#���,�1�%�R�0�Z�T0מF֛�L��x��G���6b\=� �c_�_f����8d�����W��w��k��U���/�����Tis�ץ+�TE���@0��s�ծNe왠$���&�Ɓ�:W�}�ӱ{Ǵ�0^D,,.��`��  �:�����u�=ޅ����	��,.��,?|N4����:K'�@!������p��	`dq1���dQt��+�VbɤV�"di��S�aK�ŗ?��x؏?��P!&Vl�),�D�q���B �@ql%��ۿ�CK	���7��]��,|/]W
�}0ֆjE)��������T�Dh5�sS���X�$Y��j�1e�]mn���-.��"���K���˰�T�⚆À� �z�D�S�������+�6���d��,ʩB �F���gl�o������ܪE���Q��~�z-���(&>���!	[M�6y����|�3��~�|�s��O�|/GufZ\�B��x��d"��`y����3���R(�>;�"��W,]$.8��LOOc~~KKK�29<6�Ɏ����D+�Sf;�V��/N s���U��"@�{�^9ƕ��*!�}���1ը���V���w��� 65]<�I5lV�bJ@���G�����Ǩ�V:Ǐ~�ݯ�E>�=�hO��ngQ+��j� u��V����	-�c�!����E*\Wq&4�Yg��Zd0�(���f�]���녣�U����r�\�;vh�Dwq���H�$n,�6���w�]�y�'#ɓc^��lLo����Gr�d�{�5x�c?������Kt��0(�������2~����J��Z͚�W�B1b����ݟ�'<����A��ʱب��*�m�~���qz�y
��%��Y�R����"�B,Sn�ZՐ�Xҹ�D]aR���͊��:�_cȍ�s��W��5>�G�+b�h�'�Q�gq������v��!� ��?"�LLg�~�C��O�5Hn�F4G�i#A>��X��s�A�f�������H�!���~�9x�[���={6�G��2��r�I,��]�ڡ�J�ȴ�g?�Y\��������fu�J!��ح2<��T;��q8��v� �4;3��
9 �L���©��&�����׆;7��׾r�^0���Ƨ��SM|e��(B��G~����\��wź�UMQ9�,��	��6Ÿ��E%GV��U(	��2ţ(�;wlBk�6��zl��n�� �S�����ᅿv\�(Z�%Gk�`��H��SSSG���V��^A��v�: �D�)=��� ���X6��Wr��䓟���k~w��\Th�E����Ck'�# }'ល��O�9S�����¡��е9NqL��ۉ�:���P9�+2*�+����_w��fkZ���x��Ql��b��9���}Pkl��%ફ�£x>�h�ǜMX~F���dn�U:-��^�?��G�B��)_S�щ��s����6X�B +z���y�,;�e	����O�����Xs�ꈰ4KW��qѹ���������%Í\� 1�Xͭu�.X�W��TN���@�	�C�4��G��hvW.�ԯ'FZET�pi �0v��c�_Lj�ȴ����~R��s�?|�׷	�]Y�����]�� ���I?j�8��5�4�fx!e%:��k�������>|<��'�����Õ�������*w��U����"Sm��Ts"��ߍϊP��L4|	��y0��6$*�&]Y�ǔ��=�d8�,C�h8���0N�/��ึ������K��+~�yY��cbpM�h-���ʮ�m��4���F��6+��:�����E[�k���J����1�!(W}]N�Ĵ�ߗ='r��a��@<��n�y6�]8&te�_�n}�(ߺg��-�5�����(��&�U-VV�z�&F{����J��v0��J�ܠ�*�ipj��q�rj�D�+
l��D����PR�zlGDLۂ~�ų�AO�\���Z���+_�v����U�A�3ϣ�+�׌�`��>�[vs%�!�[u�z��~������7��O�w�d��/���<���1�Q����W��f�b��.yG���u7`���jk���MOa�)Ζ&B�+yI�ڥ��k�7y�H"~O���q�Rڷ>C�B�;f��M����;��ٳA�c�Z�i�8Q��]GW�b���v]s�r�s�N÷��C�lQa�hvO�=i��U����%��佒��~����C�B����u���B"5oU/a�ؤ:@�Gx|�T큲L8X������_�7�.����遟�.�r��VL���V���Gj�uUz�
����V^�q�E[��I��k&�F	enS3�J�=����Z�kaLIf��W�����˗���<�"-qb������i�b260�7��e�T�r������k�ť�x(~'ݭ���G���K� ��?V��e�	Q���G#wK�1M4D��9����'��߷�B��/����ԅ�vaf�z��Ny�6��5�e��� �#rC�;���P�� 8v�C&<6nj^�a����q�RBS�#�P��Ʊv���Yl����/��.��C�-�}��a	rd�� %�*�rKN�
�:T���	��S���uo}����@�ܢF0��T�r��T�
7���Ϗ�j]t�3�D3�L��4�n5,?prV���=�N�3�\�	L��iL�X���`���5�̯}�B���i�a��(߻�?~���_���k��!q��(M��f�{Y>ծ��ط <�g��e1ІU_�k|%�Kp)J`�������4��zJ�{����	���7���"�G̘D5�S���D�&=Z�a�QK�ԕ�e��!��߲��������[���������]�e�Y�%-f��n�[��;$첋��Bޗd�v��T&���/�G�����d�ғN��=뻡l�R�"��|��/�%�_��(ƅ���:��`Y��XV��h���k5,f�i�$.�]q�Ȕ~���.6o9�����َ>�����=��.6������o�lR��_��P��U*H}dB�v��`�ⓞ�Bl}�Oc�3ppd�ܲ�D���(���D�f6nV���?Q�梫��̳X�!3�r<uʌ�
�̕GM,�����S99�yX�s ���.���������蒋A����L �/ڍ��QhB���EW��NV�yB�=�]NF�2�����T��E�lۿ����E����^�
��߾NT�����5厐P�C�^�2�z�"�*����"�k�	��?~����#��Jt��R[�PQU�м���G��J�<�����\��G/:y�*K	�(���,�3�0�w��OL��o�t�����b|�w��=J�F��4����"p@��2� d�l�$V	eg���S�5Е�Ui:ɚX�����¹|&(j��/gI��P� �Bԧ6���,pѣ�����7_������YNR�{hb�c1,k>#��g�Q��[�x՛ޅ���7�G��=�OCM�)�$�C�Pu��G��k�,��KAT-X3�P�@�GvnnN4ƒv���ڼĎi /�]�6
ׂ��\�(C�c��p?���v����+��
�R,�Z-h�hX�j-��<`����$b"PRa� �I�"Z�0S�bkD0Y�^���/�S|�u���7_���b�T!b�E��}>4�j��V�/�O^�B�����|����H��1�V����u�@���ص��%䑙"&W��sG:�l�����w{%��6�T�v�T�5V�?����S���:�#��*�\w��!;���Fy�l�CY�Ly���RO�>1���� �Zؤ���#�Fz4�!Y1��.ϡ�
Nc�1:�Q��Hda�"�ڎ��<�E������az7��m��������z��
�ۋ����%������`�9x�o���v��IQ��E"�X�A�K�lP���!�C8��*��`Q!�蛲��Fg]�����P���nʤ��\��{�Ur������Z��f�20��&� ϱ�aB;첱<)�	�յ�-TV�*'k�7.u�|F�?��~���)=;ϊ)<���ɉ�]��F0�"�T��dd�!�HH΅��`���~?�x�q6�x�ȿ�7�x6�����`�i�7ƕZQ,�o]{>��k�;��
8l��p�C�{S{5Y���w_c8�g%܂�Q�Z���"涊��xdvI���'ی�,q���B&�R�,,P�ƐH�]�j!�Ո(�#��ȵ8�e`l6��']��+��8�.�RXUKк�X�ьR���Ri�j��-�"gdC�}�mŰ����k탇(�G�4S�E�eYZ�f����[ο[K��;o����x�k� 3*������Q��坿o����z��6Av�p㐣�	�F�11���L�3�9��xt�8��!c4g��8A\ Q@Y�fiZ��n���������<��}�{o�UTwu���)�����}��>�������Y�S6�$��'7?�=[�Q��n<��@�V���[�K�#:�����X�.:��U��W��V��Z3]y�����r�)1L�}��F�y�ݻ��k���UW����/)x��d�u%�-�j2�8�/�����m|��FB�C��O���9'r+�Я��gj�;�뱃���	����b�1�������/����1�-��Y��Q���*�l<��߉���S����ִ�҅�ƙo�0����f�hh�X�s� �tUL=�#D�n��C�
9@SعR�8eۖ�"�g+�
n����_Q��9����&6]'A�-i`�QIٜ�1�K VYr���L�1m�&Y����O�"�%Gp��,�
���|�T��b�`"<���B1�y��@|!�V��vӱ-����V򒁉 koK�MOs1e2�`GC����K��d�S-R���S�qj����s_KۏW���r��Z��o�a/6�� �<wi~'��71����<�M"��
�JϤ-=�>#�v׫"m�X���|7#Y N���,�(�\-}n���	�DcV�R�`�Lf-�r>5��٘E�O�3SYe�FE[�C~r`���,�?�h�\�˼2�fc��v�1e��z��(J�J�kk�P,Y~�,���
�;��{�4)��/�5��cU�2����b��yM�Z�G�{���C�X�Q7%�.������l��-C�kj�=�^�L-h�-�b�pS��4NҾ5���e^��⏃���1m�8�������tn�
�1�.?,(>�5�S�ȹ_�M`��g;yߴ������b����l
�1Q�߬%cA�e�kMy�Ai�vD&�cx�J��-Y�mtd�X"I�E���x9C���&Β�OC�g��
Lr�q��5�{�հ� bh~	5b�,����H����	Ѧ���b%�ܻm9_O���!d��@��Bƒ�J�f69Y��U�4�
�K$Mc�6-�+��s�֢�U��6���t}�7ѥ�S^�d�X�}�z�6`�َ�	L5yv������\�/;�b����-up��r3������	�Y���B*JS������#!MS?��%�Li:����3iS��&Qm�jV���B�3�vC��3JF�A�p�k�.���h�c�v�L�u��%�,�����T��!&@�31O�l;��a�)�.�>ĝ�:jrjU7��e�l���� 7���+��a���o�
8�*��9G�A�RR�����rt'J{���MN�5��d�#6�ݜ��\a�d�D,�oX��;&I���3g���|>Y ����b�R�W�ТN���|[A�V
d��V�Հ[�+���u�Z2�Cc��:-(�؆�^j�����P3ju7;��6�u��!�ԄWC3a7A���0y�s��	U�0�N2�EExZ�s�����v�VdbҮuqX�{E�|�oh ��CՕp�	&5Q�X��e�f~��U'��z���`
����C�,��g:� �5���{�&��Ս�5��&,bm�h��h%�*)lH߰r��]���\�G��y�ͭ.�\��:�x*�sZO��vsm�@�+j���� �3ϓ�|8�Ψ�E=Nlu��mi��,�ew�|Q����r�)�A�W���%	��+'���k�Y1���]��
=�]�MPP�2�'���H�$���Eiw�Ԃ>hT3	�e7Α]X~f"�f��R
;���H�K^`��.��EK�ƒo��d�99*f��
�Ŭd����&���S-~f��XJ��)�f���Z(����y�٘yNgi��&��{�\ܥ�%	'��_|����ر��^)h;�o�P ITS"�Q��Nd�+MA�X$���b�,xWI��]C&� ����6�����{p��g��֨��/U�5�s���3�����q�a �-v�)}c��5_S;#*�}^4aQi��鉐6Zu�Dk����h���B��<�>��M��T���+rltŪ1����QI@�YO�H�S�/yH�eX�wԖgU$�<��;������d־�\��W�c�J�N�&bKw#���^8�5XV��yY��� �cS��P.�B4B�1d�\�2�RK��I��GP7Mz;�#���G���xg��4���Y*:&�T�B��&})���,'�MY�xj�b����x�ٽ���T��^�Xhf��d磂h���aW��]��y�0��F�#��"�%����a��5Q�IꚲG򋤖��H�%	wD�1������W��b�T[y_"��Si��B���٢���!C��G�g���*ʎ���F�HSi�S���MZ>(����ڬ&_�\6�c֓�4�'GFsF�rX^'�$bW[����N�7�7}�أ�:T.�Y�5	.)��/��7ɸ/bkfy��!,V"ylcnF����kI��`;09n�r�����,(�ʂ��y4��-WV��/��r�䰜"ir`����,�.��9&�����Z_�h2L�6z�&�`��;��P����U1�`��VPk����#aH!''psr�+^ ���9���rbB7gw��U��;6�QW��ب��j��ۗy!CEu�T�33"�r֋�*��k��&����햇ju\ k���1�����/�!y��'�]��T�sZ]y���VQ��\��}�w=fL�[az9Vrh�Mc�%��ИhCu����(:��%���"��u?0AE�x&�M��=���:�
9N�{p��c8�����0|�i���-���<�\l}�)1	c�h�݁sљز�Q�|�|P	�e2j��a��2���� ���5�#��k
�a{W0E�1"��W���k�И�����ĝ�������Gy[f"�ΎB�w�F����ry�蔕(��("X�>���{��`���t��L�,)�;1ʲ�W!��Ƿ�<6!�{��?N<q��.��8�����W����/���-pE �����q�Y���'�C�<���"L�\ds8�2R?Y��XL]����"���)z=�eQ����L�8��g��W����gw��t
.�����(�[������_(��)yE=���k���k��O\��\v��j���D��t��Gb�Ƚ�2��;d�����k�;	����������F���������^�w��7��~��r�;X7���{���{p�+���W��ct����+�a�N��f�&Wk3�~�p��+RS�없Dc4�r���~u�����K��{o�[�r%���3����%B��޻Lͅ��!���YGs��5o&��o
�'��ʳOö;͙��a	#u��h�Q&�TZѶ��M�1ˡkhG�J�d��1���P|����ӂ��������o_{>���?Fm�p�ӣ�n�S!�>4����?˱*��=�c�����m?��-�&&�+�1�u~م�}Er��D[��;�߀��0���"�I�"��B��.������L�;��s��-�:�����!f��{�O�Dy���ˏ�	�굸�~w�8(J�!|����g&����v\��w���l�	ڙ¥g��~�;�\p��w��ߠ��l��s��1��k~�
����}��(.��;V1G���.$QgqGփ`��M�D��y�u�Ȅ5j5��qf�8|j��ȏ��^DZO<��%��wn����>Q��h$f��\��	/74�6[CT}�+���(&6���^3��*:/Ml+q�����σ(����+O��:'���~��9�:���ߎO|�2|��7�L5߸ �07ׄ@̱6u|��:�k�|�F\��Y�M}b�E�g���$��Π$�xσ��o��ٯ�ת�������w���;n=�Qǋ(�R4���U��tF'��\���rΠ�Bn�Q��:/�����]w����β���׏�=덣�W�O㸕�䬔�#��[�S<���8���_�"�H���-y�zm�6[*!����ΐ�jc�R0)�ֵ�v�Gan���D_�,�˱t��S��xIP�`���q�
�:���߉�U���Wn�����������D�4�z�E�4��T�ڢ��N�Pm�ͅI0I�&���#|5<�Z�Q����������.y5zH �h��a`�����ȕjJ�ҳYKIN�Ǟކ�_�U���7q�2fĢ��E^/i8N|�\���,����<�� ���y6�����j;vlǘ�m�=M4��q�ƺNǴ!�ã&�W^7gń��l����<*��J�*�OU�擺Y�p���73!]��O`V���Ę�B�%���7ނ�Gc���R�c����0Z^�����߻_���`ƟϠ]$O$�Q�+�=L�މ�+����4�W�*���FPA^ݖuuOn�!��\��a�9����w��:��ΚXh���v����ג�[y�Xe9L���E`b:��RQcIGb,�%Nn=��X���[(���"�ڻ�ֹ8�k�u�n��|5pꩯŽ��BvbGk'�]�m[6c�3L��p��ER��KLy��Zr���u�8�4tF?���X�UJ����b�ú��bӶ]芠޽���J���VKZ%����v��ǛE��
8&&�"���|^�g�h�����q�[~�ݹ˦��"u�%=6@��v~35������;��4�7=���j5yt��wc�Np�l-��gZTc���o^��7�{����X�Z0�Zq�H�\��xP_�Xr�Ĵ��m�,��a�7%�r<&f�f��L�?�p���l3�Yg�ؽ��!^�oz��}'`�ګ�G,�+.��>�"�>|9N���e�0GrX�k�i����Z�ZH��t�n	���؃�}�
��0�v�Jƕ>�NΥ�	f�9Y����u_��?��I&�g9�¹��A]>�����o�����;Q�2b�#u�G�֘�1+G�H\�T��b~7�|>��_·nK46N
��]�㲋�����n��j/��W��y�w��O\���x+yR4�tξw��\���%\�\�Șah
�֓��6BKH�J�,z�����|6?��y��V��A�����<��^��?݅��;kN�㺯��]�?
�z�L�|� �;�߅�b�TG&ЊM!�U��N
�ɍd�c|r~p�#��&�]y�&��]�ɗ��^�-�o����L 	J(M��O}�Q�Ys<vEں{�z�$������	<��^�i��V�1���em��h��h����Mw��-<���P[G�-�?���pʩ'�7 ��~��=�1���?�c�uڙ8���`/1oxRۓ�z~+J�1,�^X�8�Y)_�c�0�����J�7[������U�}���Ҡ
�6nA�H�}�I��ûerD]�{<Y�T&��z�V�{�"Z"��<}�����N�yL2-�X�t#Gf����t�FmǊC��ZA��06=�F�m���y��&�{�!�6b�����>�r�iN4LՕ'
0���P��N/��61���c��0��Ąn������ڔ7j��ʽtEM<�m/���S�L!V�	�� (O`J��]?} w���L;�ȊI89G�[���s�a�B�n��b���J=�.*�5��07�f�&�Lݣ�95I������SutR��YdS��Y���4�b�QlZy���8x�X]�ZH�E����f�V��� M�_!3�=�Ֆ�ntM9�b`�R����{O���k�e�6�aƕ��[BI*5yF�¸��W�8��mkg$Zn�$���wCK��_�Gb�n�BQ*�I6�6�r~(����n�����8>����2Bȸ���TC�j�m���fՙ,�/�P�%��[��$Yu_A$���j��9e5z��:���lƒ��<p0�O�g���fFj}v�����hn�>r�os:L�j ,�,#�VEw~���S7�8��s1XRijK�L��.��[(��+�6���8�9I��+Ô�P����@��*�дgBNfڇ�R*[�]	�ѫ+IM	�YN��k�H̸dȘD��A�f�w`��v;�?D&}/���6|�,1]1m+%��wuA�W��>��,:� �.�9r%���P��"*xn�/0ĲH�%�i����3YעB���1�"_Y/X�i-ñ���Nb�gW+�px4:ME:i��r�C�%�]�ˑR�g����4-k�|6���AH�� MFnv����L'1�_o5ܒ�0^��q�E�1̙��>����%�D X�����m,??���n�G1/��4�5��}�}���[��(�=���0��~ـ����I�Ք:h�<jXGܙ��_�N��=�S=6`cv�y>���{�s�[�����g�M���Y�L�C���Z�GuxT3��-:bAl�n4�I�T��w�ƈzi�� 2ZG�3FA�^]�����_Y#k_���Y��K��Bh�E%�d�%˲���~��k����U�@�ڲh�bT��G2�)CLb;�?��ɩŶ�,�~i<3V���|��	5�[�N��~��:�X <2��,\ʉ�x2��vD>�P�F<��M��^̳F��l�'X�7�XԀ�G��K��YMg��؆S3�dwT�t���|�������}��2{� ��^��J�wy�PALu&�v�Y��ǒ��,�a�t��J�����f�h��ҋ�9�\D3��i󖬒l@�M�`
۪UK����/�ݬ�Yi��l�T�~��lz��m:T�k5�,�\�[�[�i�X�	��y�ġD��L_��L&��TL��M��fǓ&A��ep=��\7�f��$j7�a�Sd�Q�PP�D$$E�m���C����󥏃���1�ť���c֏r"S�?���5�f[i�>;0˫c��E���O��n�8����3� K��h�2��Dq����[�J3h��.8Øb߮:�l����P��hE[�0Ɏ��T���5�A0�\�J~_Mc3����J*3�=����Ũ�v���Psj�\�T�Y'jj��tvvZ��e�Y�+�0$p��.c,�����݁ߘ���R�BFJ�M�S��I-m�vc��u��j�|l�8��i�]*U�7baP�n�,VÑ]W�(��:äh�h'�����I\[39�HLN��&GՋ\<ϵ)�L��h���	]�^�B�ߑ���g����#U$Z����=�1C��Sj�����g�7�I=F/����� s5us�����"�֎��쎒PkRY�C"�?��ۊ�]m�j&��x��<�Y�K�+:U���k�t��f�f��,C��5���c�%L�%���Tr�^ʤ�G'He����v��R{�� c#Qqj��z��w��ۨ�b�G�I7����`�E��8�'aI(�t�~�i����1��uy�jf�.���jO[f�����D�܍Z�wш�9����~Cch�]��fn�5�Pt�&�DU{����/�FzS�jo_�s�xz��tP��Ư�g�!���j��p��?�-O>e�J���e�%�ݘ�1��4�3�d���Z��\DzL2�~���$��a�Y\��s�n|�~�j�l��Ŗ���0��B�%�ϬtP�{te�eT^�bM(ܱS�����SN�\'���$J�1l+δۄ��4=]t���B��	�X�UC,&��f{�+VL`�ʕ(TC%Jcy`�e"������ڂ9���V�1��;�Be���W��>
f���n��L�g�Zt�E�C�d��I�Z�Ƥ��zH��q��VKwp�
�U{f"�l�TK��0u{�ڤ�1j��hʢT��-|25nd-�)��U��wH��1?0�5��G�O�n��<׀�N�!ɉ��P��R!w�[�$�J���!��APNv����Z�S��	v*��FC�ZM�����[��<l�!A�K#�9,<��A�M�7Z���o��p�f�W�>��
Z�϶��rrg ��)=�CH��}�J�{B��s��'iڗM�jm>�(�M��e掺I���	��YE���ؚ٬՞�<K|;}W׿�wA�"��Ts�m�=ǦO:�ݲ���B�S��jwǦ⩊�S� �-��p,ڎ`�PS���L*;�\Em}v,�r����N��_�l�Z� �g������ɤ�ϜI�`�g�zb,&�Ȗ���v���G2�ˬ�h@S��3<���1�*Y2S�Q�iE΀X��Ƭ�����hu{~�Á2<o!�J�@��]���=�6�<ƞɈlNbx*L�(GU)���Sx�hV��v_���a�}��n���ps�0K%����K�kL>�)2��*�%bIP�źP>V���׷�%��d�Y}��\���U.>���YI���j5EӸ�T�U�`9fU~��'8i��4ѡ5e��quc��D���$Y�Q��f����4�~^F=f�˘m� ��1�	���`Ǟ��9L�U�]M��,SW�)m`�bH�*�}z��2�s�d8����KQ|��U��٨��R�\*��@�VIg�"���)���xP&Z�`�I�Q�X޳���S�@��ݘ�������A��C�=�m:��i�����g]�f$ڔt�8gI�.�(a�gԣht���he(��j
z��,S����������ʨ'��MicS�d"Q���A1fيI�P��pkʱY��H�-dHk"�Qά���f�i�bF{e�:�b�ٽ����1��Z���O~.��mHfg�b��"[7c�.R4t�PvB�S���gFN,���4��FMP&�K
��{��4r�u��{�9�t�qfy}qT�gO�56|����~g>�g�����=���
��bQn�>�@�'�t�5�fo6��o�Y�)�\s�k�m�d ��G��f )`B���S���ȏ
���=�B��i��a"�@�0--w)IV�jg��0��3-4Km�je=B���d^[	Oש�B�u�NS�V��
Y]�$0�����ޖ����2�$0:r#�Ly��b�fy���p�H�e=�M��3t�Y� �D6Dq��
�m�HyRR�Fj�����ܘV�i�΁����P�ˏ��t�m	�����)���!i�l9H��OTS�-�Z����I���+5�:cΣ�.Q�����NK&�.�2��_��+�{�pjd��[��\�<fe#EE>��06���רFI��@vl��x~>�D }8�y>'���b�_������J_�fTE ���$,������Q]�mnik�x5�g�@ǩjL�����S�F�l�+j�԰�e~�����*�[Q���\D�*������{�pN�4�:ن<��X��.�U��@,'1��b�9%�˫А��jH�|�Y�c���g��� G��`��t3�4_�$�4�i�D3M�}%�=��E�@D�1fs�����	ztݢ��rSC���RfB�D d��_�
x�����j�tt�o��;��m,]o>6�GY����x,�NytT�挋5|m���pJU�Ϻ�cȻ��E�p�Eb%lD�Qv�f;%��2�8�o)��9���N�xEF6Mb:�XFY�܀����9;���Q��M8$J���&|��;�"��l�*�\���Z~�d��d�A���1�;����_�����j]�p.��e,'����Q��I�I���D)[)�4/�-:2�,��r�Y"V���7,s"�*�zu���� 8���u%{N�k�
�d��'M�O��f&����۠)Hb�VB�9�T�ihW�*h�A�(���ޥ֘�?���$�+0�6!/!���`w欦�65�ɓ�yyͼɵ�^(�/C*|Ij2�� d���u���NL��TK�r��Ӂl$�.�3���0f�%�R�JD�%���s0&���G`�,��؀%�z&3o#G�5�-�:(��+g��/+/k/�'�0ǡ(�f^�C����k�(w=8��7�'��Kר��-��p�Zu+k��t"s�U��O�AG@n>ߑ�5���"��vC��	��0A&(1�SqR�������f��O6�Y�T�+�u���ԛ@�SG�K����䞺ih�H�^W⩮�0W혓�(X�A���`�.8�RDCE6M�`�]�-^�G�rd:6�L�w�ɵ檓�I2_ej�2�s�r�5��h�S+�y*0C��ɤ���b��b��Uu�%a����[�=E�u�[�9����u c8j���cCs4���|�/��#�8$d�]4SB����=�;m�}B�{�N�i�`�+���Hh8��	4��8�<�иè�e�ш-���X7��	-'�̙�Yģ�ڋͳK��Ԉ�蘒��`Q�}���ibx�X	mG1	���E^o���3�Q�T:�}��"['��,�����Q�nhh��:�M�I@�fV�(��\��ȘoZ��(�{��q]ߓ#�����6�v����5�FNO(H����b���z"���Wa$ECО��B�]��X)��2�<�ג�9����O3�f7҉ɸS=]k"g�+M���?��S��(3a$Z����d�b����	f{�q'	�'uc�IO��H9@�U���J��.`d	�����O�V&b1@�s�`tc�\7�ϹCb�9i�T�Փ�CS�x�ߡh��Wn^�"Q��y?�Ė/jy�Q��p�-TGdG5v��D���f�i�b�;���9Vx�DF!���5NJDǸߍ��|�:��sI.g�.�0B��F��]Y�Ey�1�gŁ��j<�q��0����h��>�h̲mu�K�����{�%��A�a��e��1���T�݊�ĵj��YBN{'	،v� 	��ߗ�):�޿c��C���׼t^��r<G= ����~�|�=��m�[��"�yG�۠�.�Fԏga �!���W=��:k��� ��Ҵi�E�p.�̟x�BŐ��ۋ�ʊ������H� I㚝h�b#�^'�B��=O��@OuQҸ�=H��5�����������S�v����Ǣt
�>Wұ�fKE��g�G=���C��Tk0�<���v|�ǳ�Ug|��z�0�[q���\vT>�|Of�4~��|+V3��h1�Ӗ�Ԛ����
�o�ƻ7�MC�9\ks3N�&?��������a�El�LD����az�?�隴��/��;�FF�l6���O����?�p]o�k;w<�X�Vav��7O�����-��M���շ�cc��x�ٍ#pm���6�s�|�������_L��%�\	�\��_�η�������������߽`>Ƶ���^��7,w�,������۱�T������9�\p�,�а��r���߿�'����ј]h+���^�����6��f�v}����N��/�(�l�Y�c9��P�0�(��8��_��:Ђ�a�S]�k�A9�ꄫ
��rX��2/?����A��D�B�GqS����Ǳ��)�1Q��e�x��I	,B�l�Q����c�ޘ(V�rf7��/F6��wʬ���֬Amz�����n{E��n�y��W�57s<�q�K�D�^�Hշ��q�qL	F�T^YL;�3�U2����ɏ_��|w(_*�_��bg�b�8�4ʗ
y��d�/�(�cJ0:����8��b���0q\vC�>�sD�'�v$ʣ�>����e{�cJ0d��O��xK'�\�p�z��ue�JQ��'ը��7��q�	�<��4M�M0r�eJ���/����a��A��˭��֣z�k�����Gl$��KO�^�؟�`���8�#]47�aG{.�0KGq�ɘ7D�� ?�C�����R1����O?�`��w�r.�����V����hjO�G���ڗ��Xf�8��_�c �l� ;vY����L	�Qǔ`�_i����r^�c�1��U20����5�����܂1o-^��c�s}�Dq/}$Ird,|��_��1O0�Y��s]�h/����e�d`̋O,��V�����Q�,�bj�Ʋ�ǔ`d~Vl��5�?D�Aļ&��I��|�M������Q���.'���(��m3�	�V����jy�Ϝ#��.�qL	F�[fa��o��,H��lCCCڈ��l.[ȟ�����5���pS�Q(��Z�P4E�NҞ庶��z��Uv�zY��-��2��cC�,��]�V��Qǔ`\|�ş���V��eq��1{�r]���/���۷�#BY��7��n,���K�X���T�3r�8���6�o����q�eU���8Jc�ڵO�ǔ`d�h��c��W���3j�    IEND�B`�PK
     $s�[���� � /   images/bf314729-9196-4b76-b154-4ab11fec66f9.png�PNG

   IHDR  x  �   y1�   	pHYs  �  ��+  ��IDATx���eGu ZU'��b��je@�D�1D���/}�`��؆��������4k�`���<x��a#�ƈX$�H���J�R��n:��f�
�{n|�V����sn�:��کv�r�l�l�<#a��o�l�<Ca��o�l�<Ca�	�;���Gn���O�͛7S�~���n�l~�����q̛�oN����
���:N����Nv�&Yg6��c���LDyF��B����-��,��	���'ֻ��	�Yg�U��x�W\���j���x��8��r�u:1��23���@w���	a#�8&[�l#KKK�Z��:���G�6m!�g����!�J]_dׯ����ݞ�����s�ya��Hw��e�1'�9֞{�u� ��ЗUL�Q�e#���kc���#P�5!�
�C6 N%!��/볨�I@����lD���ӄa��9,c.i��$5'�^���$�	��@u;F�� �/�?-����$F��p}w�'��Z�0��+_��C�^w���>�!� k&����s���o����G�Ւ��r�7Ά�nK�dzOB�c��O��O*B�N}J	u=B!��$�"µT.�k&��꽡@�T1?����q	�HBe��|��aD*��V�+Yf �1�}��|G��2��k���c�摓�'Fί!8�w�8X��0�q^#���~czGd�`]�ۯ��g`c�!Eob�sO�����w���|���������m?����͉������ٛ��ٽ�R��Q_��=�N��A�q��v�8�$I�}�*���8Ү�	���b�A�3D��p.��n�ڊjc܉H�S��i�S���H�+R�'�x���(�x�����g��t�t���OY��0��#�-�Pw?���<������sg��O
����]})ۯ	�y��­��ĉ��'Q���۷|}�����^��w]}�Ս�6o��UW�j�ā�WJ��pl�ȋN�<yF����:��u|P���S�v�H�Z��ȰH��~|K�W�'��wK�Qc�RI�����Q�J���ݖ����XK�����kӤ���7i�8����ܰ�ޞ:s!k��jޱ�-���f��W�s\�رcgA����n��?��O|�S���-oy˒��Wcxh<}ӛ�4}߽?���wC�.l4S��+L?��"qG�&n=,���<�y�ylx����~��LK�\�ez/� O���o �#x-�����I��P@DQ��GѺ���@�?���=^�)�=���s 8�����~���>���Xm�c�~�J�<���W���;�\ j��9L2�O�����ˍ��I�Ϥ�?�9���}j�4���c�`ĝ��Se�]>???}������W_��E���m����ɟ��^�W���e�aʭVG�q��igx&�ɇ���ۀ�A���=�!���,��ʾ�_T�U�H�߀��@���X���o?cii�;��MG��]Y�q�8�:��^�`���p�5��p��:�X��t/����Z��+�zի>�'�-$����[��}�{_y���@mس��`�� w�9�n]�V��ҵ�a�d0�aD��dn�R�mC����~JC~��U�d���9v�T*��8��j���}��}���I�:��ԩS/��l�Pm@���t�u�l�D>[p�_�S} ʍ	����O_F_��y$�t�
�ϒT��_��=�9jS�P��7��~�l�}o[���Pj����2C�K��3��w���'W��܏x2	��LJ^���K2b+�*���T7�<��a�.X�hOYh��摸�A@ڭn-��=�����k�B�֨������ �Ǐ;�������m��j��� �7��@�B��	%���{�#���[��@M��]�F>�|ҝ��A�)�ɸ�<ۯU��n=��*3-�I�J�J5H���������v���D�i��H�eЅWjn����"��߀Shn���GQ�,����|�y��dR��~iyy�¥�ŝ�f�у]���S�+6X�Z�۔� �p�k��"乿����!O�G��*l���	W`7
�_�TR�p2(�n�R
��o�@�y�t���f)��iX��g�y�B�3_�T.�ڂ�}lc�i#i~z�)�0e+�\�3-lw�FU�Ht؅0����+'*����1Ǵ/=.�$PvIm�v�tzB�8��r�reb��G�v���f�l$�����WAYW{�=�ҼOXO�4�3 ^�2Ix:��z�e0��OY$�R�HF�X0� ��Ab	m��|>6���Vw�SFg.]�#<��x������P�<�s�ݱ���j.��l��QB/4��d�V��@�Խ��5 F5����h�[.���V{>�]0n�*���@���_fi䠍�y�^#�:!~Nz��� x_��/|�K�|xT�������tr��A!l#�N5l�%ж�333�wG�Ѹ���@��g'��퀺���~��������k_�y衇�5�\#���w)�:uJ�3����`���u�MX�r�>��2S���Y.��'�!Dq�G�F�A=R�uf�'��C"��-���&�p��D A���J��r��І��>�a�*����J.�2n_�Z��jQ�Ў�D��ԣ�*���#��_�
�eh|hc�]�!v�
�Rf��:����"�}X�=J#��oG����'�:�Ƅ��l��{i����=IP�|�O���X?�Y%\�����C��L��S��%�Y�M�J%*���tNK��N���a�,�p�0v�\�%.Bq���N��i]���!:�j��ҙ���b=�t��~���&Z�<���7�(	ı+�>��*��L��Sg�{[��6R2�V����#qO߅��:��b��1#Tt�$���,�jI�A��a(^ 4�J6/�z|(��"�yF�vx��>��Mp?V����[��������>�<�����p"�4������W^y�я}�c(~�,�(������[���گu�F�^�ϧu��I������b.�b��K����&{{-��o�O_X\#mY��0�+'̳e���~���5�����{�m��s_�73�^^*�� �Q��bá ���$4�H+���
���`1�Y�mp/�|��͛7_�җ��� �����	�=	�D��6`6`0�1�ךg=�7�����
���{�?��G=��V��6��[���8��ۅW���-{���7r)i(�隡]�j�� kKʂ���'y����_�ћo��N�Om<�_�s��痖��}�� �}�^ܦ+��+++��V|�R��b�|z���=��|t��E�'˃��7֏iX�#R���}�<�����vY֗|9��+:1-{�2������b�4[=���>(O�s-��`yX����Ԧ�o�i���x�㦷��_���XƤ�������lP�Є��Ф���J��	LM>m�{4=��?k�'�e�4���ەϗo��vr�j�o����L�k��������jE�~���Q��������� �|+��3�.?��[�}�=�ɮ������8�Z1[j-��б����^�������?`���>����?�������;y>4v3t�l�u�M�@G*(�S�Mޘ�+�\�FS4�x�\��m���h�Q�p-�c;�m��ڕ�	�קж��L�Z�3B5���yU��z�j"ԃxӆZ��9�f�wv�KB]^͂.�s4GA���1�3<����JA�4'<P��
���������h���P�p S�?�nA7v���(a�*����ȩ��L:~����x �ܽZe���$pH�R�L=֋��:���u����r2ܪz�ɧҍ0]��~���J�4�r����S�{�~Of�i<~+ R��Aa|�o���zcyT���9"�j���a�M�O�cH(㸐L߳lli��>�O�n�h��18����wC|����J���,��-[ڢ�i��|�6Q�R87����jj�b�4�7$�L�C|��h�7Cp�N\��Ӧ��o��9i��sU��ǧ-���`���1��:�xC;)�{H��8p�q��_Rvs �(������_t�9G>��O6�ſ���8�����c7���}���m��؏�ZRe��tCZ����C	�9�������ceH8U�s��چ�^�W|�W~�W���B���L���������]PvmI�����@�	vg�M�u���CI:꣺"ͪ=>'�7�v�\�	��H�qr"Ӑ��j=#̫80|0$��â�S��D���(��-ևx2��;��P<�nl~,ȧ���4����f��b�J�:2
�׭rK��MI6�fqq,? ���,T�8(�t6��.��E��-N�������R��"`�'M7�EuS�oU��l�>�^T��~#%�!�1���ƬDb���si��Z��c�'�߹��}�I��<���s�w�9�� �W��m�{;�E��<���s�l�T8ı��y���U�~p��D'	L�"�|����m��5��}[�K����,:q�ʵp��-��˴��`�֏�1i��v�)M�p�����|�]?��7��6BN�T��O��c���C�=���@u)����5��>{B�#��"���yf�þ��l�A�9����K��ɾ}�J�^{��`��Pw�;. P�a�D�C�q@�q��m��Һcҭ�XS�u��wQC��=���ȼ�`��fS)��ϋu��l���U�ly���u�yO%�Jby8Q��C?������@��q��
���q�����f�*+�<�a5�Xk���s�f�[�w`���͝�f���9v���Q`��֍!?�A�Z�q�VP�20P���sA�m��w�܅ʁ.> B���~�]F�������6�g$%�[��Vb����E�:���/��%(�W���{É'�o`{a�� ����#1?�l�� �=��ը�45��������'q�Xaj��B��x,R�Wq�Y1?Z���xz������
KP�x�8���d�������u���<~�}f��+�y���nc� X���d���ݵ�s: �NˤV�>$�vN��h8�H�@����l�>SYYY�ܯ����]3ܟ��L��;��_����mG�_5!`좋.9��x�_Zo�?.�=	�U������}�c�9r�� ߳�Ν����݀؀x:�6�) �/K���T��\��Y9�y��m�Š%n�ߞ%�C����瞑�{(��5+2������4r��/��{n��������Б�mOMU�qT�'��2�px��6����!�^�;Y/�Z��Ux�����o���\s���%H<|g�#K'7�؅�Q��$�����w�uɦ7��3J�ҋA��Z��������؀؀�X��5���R��~� ��{/x��-��?z���8�l�Тǩ�?�
v_�w��$���/�����|�|�#�n��ƽ����9�Y>�ώ���L��!�������s����o�#ʇ>���[n�s������N�y�ZCJ��0�����l�J+�v�z`߾}������M�r������tW!�h���L�_�k��sY^XX�B0�z:��,o~�=���f?�(�׺���q�hF�oݺ����Z���+�_��_o�۳��+�â�ݘu���a�p��OE��&����ŧ�*,�:��sܜ���1���j�Қy�w�	{r�^4�l�f�J�h�jM�^��R�i����I]�
�����ٵOąո>]�х0uzkƈ��{i4ȞA�o�)�#^��&���+'~����<���ؐ�|��a��p1q�7v���u=��<��7�W�$�����㹔m>���&떾듣�h�	;��c�+��
,\(�!H�^E%�ٴ>��MA���̟��z��8Չڳ�eq�A%q���`�I�@&�?�VW<�J�����4I�!�p�Kp� wq�U��e����b��.��D,Bsm�{
�#l���zW����υ
(�`���c�g����ףO�������]�,q��&w���g��q���wא����{IL(��	��Ku~5�+Q�4q��cY�1t��}w#��ru^�o��L�/u��X����z�z6��NĄ䉎T�"7I�HQi;�3�y�E��d $%P:K^��C�x|�qWܡ���e��#�g>�H��i)]�+��᩠�1Ȯ������d�.����n�| ��#$f�.Dw��U]��ꯓ́��h(�_��&����(m�G����jE��
�g��$	i$v�%wi}Za�#=�sJ����$J'��%b.D:�+�Kѝ�� ���}��S��ab�P�a=&.�7�R��	�Iߚ��cJe,��2��S*�<}ǟ�O+��K<��8�c;(ɢ�=-q���]�C%�;*l��*��l�' )�aI���G�l;"����^髂��hr�����i���A{�����h^:�Y��`�h���T��"6i8cV�C�
�MAJ회]�>��	i}qc��H�
/�9t{�.�8�r�]�Vj3N���t��~�.|fO]B� rP�ԦX4"ZA�ɺvї����qfq��w&�+P(���t082�x/LL��mW�=�wϞ=z�0C��j4��Cs�<�V�VoB�]xy���J;X�s�O8�>I�t�rd����u�aÐ>�j;[�5_�cN�K�yb����홑�����vE�C�]H�]�O����]mnqrIx��ƙ�헱y��k2	ᮐ����R*�ۡt½�O��U�qٻ*�ql��C^�֓Us�|U��m��J��'<F�앴��)��ca�oj�[t�$LK&�g�O,H҇!����S��&�>c,O�e.-����%�U��ԏ� ���I�=c�>��c��5ƺ���&�(0�ɯ�ی�֋j���gԫ1ь5�FxI��Ә«D.v��"��u{�d�^Yo�N��ʢ���x�F,��a�l� rU�a�J�ѐ�y��L��<��O歂��� �/ޚ�����5���a	����@��%�H�}�Z��ޓ{�"�<��ܭ�P�'?F��Bb�J5%�������tz�h���J��?ƘS���v��z��X4�i�H��d�*�2U�H�5'�&���S��恧��0h0��&$5�g��PxǕ^��'l�rq7�5��R�jAv�	�2��Oj���ϭ�D�r9�V�E�-q�r�,N@]�u�|�]�L-Q0z�q������6-�u�L�v�g�ړ2,��+�#w$]ow�`kV�יY4q����
��Z��D���M�~�߅8�����S]���t�s[�B�����x�룿(:�'D:�G�����F��!�Oq��~f*&��p��0\�扖��yn���ES�=`�`��cw�-Y��b�Ԥ�(d�	M J���ۘS�N��j���5�D3e���p�#gRH�l���Z!r�G7����_�z������R�*�)R���]�a���C.=_�U(fF���C0HE�g�u��Jh`�Gҵ����U�T3��v�q˳�Ί�Z��f=���r�s:�=�Z�^,L���+�+�W9E��rp������L� *���M:x����)������@�Q0:��(9NY��B�X�9?m�n8t�D8�$""��^m��8��1�D�3�3�0}M�B��Ƃk<��� �;f��u9�Sh�Z��B����)�.�f�Z�Ŀ5�u�7��8�u{�J� ��몀ǁ�v��{�'��%<��m�M''lw�F�f�x�D1����L�6	ꇁc���l]�:1Tu�A�G9�(S&�RG�IMG��AH�����(ЀT���՚�r��-��a�f$7��O��w�k�:j�P����E�%i.�&�-��|��w�D!��53Z��u����xH2RD�qC�C�\��D�:⑼�L벹�+�����L4^yZ��Ig��R�[�#X}�9�� �'�$��i�a+�LRuUM�mc�I��\���x�u�Vyا��CY�-T�my��\X�z����3J�]�F�$k .��4�%!j���~�)G�r�R5v�9�6E����s+1?s!�;����0����5k5D�	������&��+�g�p��.�95R�1��,��dz����{�V���mI��?�!�3G��|���M:0��9u<�IN�ܘ����i�z MhLJ9�� �%^Đ�!����vN�s�F�{�(I(8��cH���Pq�{U?�����x��- g��"��~�`q�ұ����ڵx�೼`��ˇy����8j!/R+�]�qȌ�&H��+%�'�����v��"V�#�k�|Z���X�KJn,� NĴ� �SO�K�WԝI�W�uL�_x��#�J%����7���*݅z$sus$����zLy
��<hZ�t �\N�ڜ�8t@��+��ҵ������>j��vsg�}�҅C��,����%	�����Li�=X��X5F`#&��ߴ����샒�-�I0��b�eY��8�j���o(B?�WW�7e1�ށ�����߃��r�*��kx�!��\����NS��f�k��\8�,�Y��=��"� y�G�4TR} d�=m){w����u��e�Q��^�.v���C� 
�7���b$��[+��:�D��t
�^�]��L)p��	�����X���c*b#�h�p�=���2�Z���^��������+ ��u�X�:c��a"������GI����1���R���H��e���f�����0R�g����w�"����'���IR�Z���w�q�s�Lﾩ4��`��1g�.�~�X�w#�fK�
�����h�M1�T� ~ُ��n5N^��.�G^+b1��C�ne�q=����ឲR,EG9�������Ȋ�Ĥ㵁���%VH��;M�/#��pZ���J%I�4f���;E�8�r]���c`|l�HDB��L'�W[��<,�s�o������z((W���b@L] �����7�� �&�2���ν�R�z�M���o��_n7OtX�M3?p��2�5���#��J�:�ë�.���v�;e����ca#jn�ߠ��	��Ͷ.�#�0��-�<%��g�?�#�0�h� �P^]��1u��,�'x��,A�x�%�8M�B��
_��1r��O�ѱ�+�-�������sI{�c���k��Ȃ(P|����3���FP���׿�����׼�E�[����de�4�����#��>x��o?7G�������։�W&퓻�*��5�"�c�3�Qլ:dy{ɻ}w���;+�vy�O��)������,Q���HD�6�`�`�$�T�S҆/ޡ�}���e��HhGA��s��t9j�	(��%�͕� �J��^��&� ��,�0��WE�B㣶c1�X�~7Q���{`� Nǁ��Y�ntdYT�=ɖ�u����?�/� jB��.��y�_U�P��k�F�hXjc^#�^qcS���B�1���[���-{��g�/~�O��;��3��=�v�W<�����D�^y���t�4 v�;@0�Y�V��4|^![7�!PSO�%̉A �јL�yV�� ܲ�,��uK��� 
g�$�1鴥L�Āք�B�D.�!h���lJ@Xe>H� ��V��b�T;��#���,�� ��d�yr��,޼��~d�S�V�:'����%	�~ϗ�D�� �#Sg]��m�]v���������Ǧ.���;��7AB+���"����V@	�ȃ� :�8 -�S2`x
/��:ٚC���E{��hN�o��(Q�s�g�T��'���j�č�� Ϡ~�L)+���Z:a���He-�%@^��w�����e5��+A{����T W���	צВ�4B^;��������_MO�����߉��$Ѳ�I*�j;��,Uc�D��s�Ww������gw�G[�����Sr0+?�e�JL��$l�B�O݀$Ǚ�pA3��	%XB�9�I��A�� %<��6۲R-I��4���}�r�s���w,=|�}'��;I��9Bv@�i��ق�D���Ͻ����ߜ3[tO�z�.�t��縄{%ޚ�h�d$���$ B1(�0������D�Y�YF�	���@���{_-��3�n	1+$�.��)8�#5U	c�T�is�eǔ���A����������GO�s����M.�'�+�1��G�8����Q�kf$21������b��`$�cN�nY�Oz�v�t�9�|t��Ϻ{z��Wәs~�TX~I��hP&��H�PaU��Ip���D�m��:L�%��bӳt�촞iw����e�l�Z��^��DJۥ��h��{�b�\�z�Y���+�+��G�S��(����v�1��9Mg�ޯm�z��ӳ�s;/~G���y�:��I��!`�S��&ԔM{]5�����A����ΈH�e�Q� 4[2ci�����t�d��8��7˘]�d�C���H�{�~��V�qIL���������Ն+�~����!�����ک�F��ش��on�������m=�e���oqj[��q+S�|�wѠ�$�p�Z�mˑ)�E�!^%�(��א����>���+w��%�T>$�����e��Jӫ�D/���*�}�xU�U��\鬐Ʈ;�J���!�t��ڔ�M{O���w����N���<���[y���2
K$OH��+����~p���?����=S�_�	ۿ;�r�Boeٍ�Ir�WA�I@Ĉ��h��	�	�JA���q'��!�]_ܱv��V�O���rO]���d��Q��J�_��bY�+���,�����IR��K�J�O���l��g�y�<ԉ�B��;,�k 2��.�s�χf�	�>���|�h�8��b{�_>���IR7��fw|��+^���������xꥋa�{f�&P� �^_J�E�H_V��[����KV��&r�U~�q��޷?����ؿL�6�c%������^�~���G�en���+��-���|p�J�{lv���o;���s��"�w/�ٖ�!Lf�Lb���:p[�z~h��mYvS&�b1ץ~iž���J�p&�|�s%C\�S_��
�11�͘t�3���o'3'��M�t�'��S�����-����[o⹒զ+Mo����/��󊤼�y���ǖ]r���*�	(h��@Z�=Qb��BO*�	%�p�w�+�Pc��q�GR���V���
W��X���6�{Ƞm�����XY�a�5c�Z�M$x�<G�fs�kϙ�t���(�?���y�w���#�l�;g�ʑ���H筩r��_�Tq�7�����g�Hi�MJ�o4T.����s�Q~U���@�^�*�9�C��@7�� Ф��E���+PSL����W����\D1�o�)Mt��4h9:f|���|�-o�>kv���)��M�=�����]�.-^��|���(X�)�bg��ɺ�h(� �+��lv	�
E���3v�:�˿����>}�Im۳N�"�[)��0j2� ����J��d��� ̱��}�O��<_ز��$���T�� ����jy�����7�3�|�/���o|����Ti-m��~]��3u�{���tf�T�מߡ��P���ȱ�$�<�\-,)?iV�i ��*|3a=x�yN),��e�/7��qh6� \*-JSU��l�H��Zy��~ij�/����~�����+՛Qk9��������j큟���?<ј��Vw�M�۞��2%�Lj��KH����V��D���Є�M,��@��5��"�;�þ��_��sM@���Uw+��g�y�	�吔� �W�l����?�y�s���黿���<��,H���Z�~M��_�u�ܻk���U˯��삸��D�X̉�0�H�+��q��7}A�J��I]��Hv�߀-�^-���ȕ�����ک�a*��[��V"i-��,
%���o� ����>������;�w���݇�.�,�ܤ�$��5;���49�Ǚ�n�w�;�@�?�����(J��(!�}&&����Nח+��T�J��S=k%���`�D	md���告!�H�����9�0��{^\v
DƸ���g���O��}��R� ��,�ĸX*Uݠvƥ�?�r��[�*w��DY�df���GB�r���'�թ���yg�Uv:�Q_u.��c���Jt&v�'�-�u1Ƭ����jZ��*�#���/�H|.�$p�7��&���I�dC!�HAb�d��2	��D�2Ss��6��e�|����E����b}n8;��@'���ڎ5���V�
�K�S љ�2wV�>j��gڣeR�g�/���k���S3�I�W�5L{�g�<�}c"�X1��멓���49|j�2̾��������wK���w�&�R1b�%��+�V�#+3�W�Qq9�<宀>�x$�uʵ�̄�iH�ٲ�
�gD��_���KrX(�Ahc!K��8����Z�"CD���;�t�;kM�\��n�]�ԩ�س��Je	��%jɹ)�Q�H��M4j�KA[-Bns,S�DG���	ʓ�Mw�8�?��;�8u���+)�I��eo�f�x&hT�0;xB�7�옉�&��(#�2Q�n�UwР]\���q�3�)C��Mj�*Ni
��4�j�Y4͸
�DᑚmQ�$9�t�nx���ĝ�2��΀�I0��U`p�ԯ��(hu��s`\Qv[����	�u����h�v�C;�X�$�+/?���؝�1�սJ�ՆO��Q��Rf�"�[�6;�q�����A�M?� u$��cھ+i&e���t:1�3�Ru�M�_��3�?߶���F��׬F�uD9O\ѡ�ྋ������8~r&�m#��x5})�a��!l���tH�z���A��A���E�M4M��=��q��p{�ظՎ�w��qw�9l�y�q�)��uaJU�b����5�����'�[xz%����5z��j��K�Y�e��v�.ou��t9~��I`	.�삇��EP3�l�$��� Q���l��o^P�b'��)� 
�a���ӡ�B�F��K2��U.�@�B��T�)��3_yt�`�3t��>�'���F6�p�,���v�̠r�W���3�+�������[��N�*�`T��]W�+�b��fԛ]��%i��0��x�M��N�x���z=-*O
���Am������2�B�	3Lq����N���{�O,*�m�iV���%Ɔ���P�w]s�ZDd�vѮ�Z�LjEI�Y�Xy�WmwW���6�k/]|&��#Ǆ�@�e;R�k�AruM~e�HɈe�]pl�@�JAP����?��&44�1���������S�y��*����Y �݃IE
��s(Q���D��U���B�Xt���&�@4(Z[��9M�=�@g��Q_��A�#����7���ȾB����>��=g���s�RB������˞ ��B���5������r���7h�Y�[m��u�u���_���F�Q��I/qV�%R�n�*�K:g�$����[���iI�_��b�a�p$@%�'"L�]����5��4;�N���#O(��S�'���:�]�-W+&Z���U\�O��F���ߧ�w��0�v��T��{�j�+h���m��ʲ5��g-�M���AWB�](�*���EɽǦᚅY��f������8�����k%,(n��3�;8U
99M`O�[�#��ٺ��;7��dqz��4fJJ��3NY���֫�E��8R����j--���̞7��L�H.��Q��i׳��+8�u�?q�&*��K��ȹ���''���&����!�9�@���6��H�=w/9��;�	��8j�����)L�p�*�G.�)O���oG���%𲀿ޯ�1�Q�˯r!�<iG����,��.����Ui�l��	���͸��q�I�;c{�0)�E�A����HqQ�f���6����҈Dly�>���m�&��8���)k�ɦ�]���;ϲ�$jm��"��0в]���&%뚼B�s����0��ì~䜁|���������?K�F@H�"ؤ��F��ļPEbV�x�$��Ψ�������z��$Q6s��_F놮���8e�)���T�90%U�C��ri7j	L�ͼ�
��Z�%ƃ��P����<a�֖�U��Z���e�W�*�u���ZѽI���YJs\B���v՞�5�~3�l�EPD�Z�]�	x��]sB�"_,wr#�r�D}0�d�'z�z�X�%�aJ��'"er��`{o��Цh�&EL� >�����`iZ�Dנ�S�"��u���t���nO���o:�dI���.����.W���D�RMz�3oB�^5٤��H4j!˼g�i�+�^B����#�@t�Q�?��!��~yq5lX;�eՄT��úe��/�C�3��;ه�6��/�:�*�@ #���Z�I=�8�	cє��\b��p�����!���$�
k�,~>-�+����ha�ELM)[.]����V=��������;�'ݻs�b��D\&ڛ�C�=���[A��~Z[��^X���P�DM1ѝ�ϫ�7i(�2S^'�6h�w�C�S�T<��|���S�!>�H�A�Z.�%xQX�x��1�(X\nʤҴޮ3奀��5(�}���"F@��oB2��K��
M����.M%u��w������" 	�(&3���M�2�GW������ے�a
����^�cSƾa���e�j&Tlb��|qP{�����͆ �ِڭ�n�kv��<����7"%_#!q:��6AU%�������e����*�sj�!�=���p�Z�ZYrh��̊��# !��h�Ĉ�Do#K\,����]����BQr���
�MS�HT^���'�����qx.wF����x��M�����jw��u4�ZNl�7~�c�
98/����Ñ�5*u�Y3�n&�&�6��v�{:/~�V������"�-�eQs� �4��D3�t��2��l`�D�qr�:hW�@5#��]/e���sD����*�Ձ��L�5W̹ H�q,c(�jC��R�M��"�M�Gŕ�����g��5�͸m�A��]����JL��]����;ٻH����4�ki�O�6���f�t���*,31�dH�q3�/l������z�D�Ԗ3at�b�N<�њ�Txf��a{��z�HW�	�^�V@�Ç�T%���NH�J��$���<�\ו3[2Ĺt��)l@p6]�&��%�� ��c�A6���E-��M@o��46x��MN/�M����w�]�nC�����W'ϐ�Ҋ��t�_t�#m)��.m�E�RU�WmH�X��D@2���9�Mx"�m%�F;�NFcA�����܇�Y3�"�ы�nB��8�`���
C-u��z��o=�@X'%J�YEeO�Km`
f��4�.;�T�h�Aٶ磍j4|>~r���:Ep�o6@�v��>|+��LT%�&Ƹ7'сzr$	��^U�em҄���mRoSL���A�NQw0�!��&4��8a(^����0MFj��#
 o�H�%�?XP�$ی�-���0V��c=GrY��Za��]��r����e �ӕ�$i5�I���L�ߖ��mCXU��]|������K��:��[�[O	��C��	9�§ϔ��s���G�i��-����	�+F
d�$@��[R�R(n�F����i�al��n�U0��<4a��'g��_Y�P���u��*�"u��$(� =�ݛ�)��$)�����q��F��@�@\EU
�ч	�:	I�OPʳgJ����kW�9ax���<E�\�
��D�m��~�*�K��yΜ���~��z�p)�u��S�~����s�40ӆvӹ�0!u��YRR�4sd��(	I�A����G�P��&+��oÄ��w)��;f�h,J/�h��������9��d��hB*�"�7sb��|���N�P*%�����6�a���'zq8IE��y����O�ax=\��]W?�a`��l�'R�Q_Y*w5u]/6X�����4"�2F��I��jG<����1LB/�{��=���A��k�v� ����}��R6��>t��X&1�an��n�[��VA�I@r���C՚&��ӎ�m��&h�S~��K��)ǰ�N�-�k�8&�c�m���5ȴ��؏�0�XF8��RiE��yn �(�7�9���)k�)nY��T�AS"��\M�a>�!W�)��J�".�y��5�W�k1�0�멎�E=Q� �MO�0�)N�ٸ�m��{ͧ��6�I4�h�k��N����
W9�/��l(��s�W�w	�#�1p��Iɦ=g���?ڎ��Ch�h���%c��#��j���]N� �?��8�H�F��_9�\\�$�jQI,�m9��6�2I�iw���":2Sʂy�;��n'!�+H��Q�	��%}?~�����5��Q�``�"�������=�\��������N�A< T���!���%�?8���z�߇����4��Z�N�3q��6u���D�@�,e.yЇ=g�N���J�:�	�����/~��!�;ʙUR<�	T/��K��nh������hK���j,""H�.n�RY���R�9Œ��t�6}Wyݻ)k��3-�/���s���m�1�-��*���$=��zt��5�l4�ä��h�Q�
N��O�c��@ �����͵SOs�w�q�Lv��J��F��_'��T'SYgI>��x�%�*�al��zntꕒ�H>>�vap�]0�!��c��<�W����uDx���Wc��K�mE�0�^�\hx��C���#��"��N� ��j�S�����G���c+�+!���g�]�PHļS�y����C���-Y�}��z4p:�ڎ�%TϞr��,4[���:���&?{����X�B�T#(<0f��y����ط�P�bѨ5�׽�]��ۿ���J��V5*�	���e��Augx��F�� *e4q�?��葄/��27���ҩ�e�\(KD$�r�:�7�nD�S+�+���s�Z����d`�8f֝�X� �k���JS�h�|��S�!p:	���,�U�t���J�x(��w�r�M����k���k��οwۆ�?�Ձ7�F�d]i��DO���wm-@�z��ס#1���g�D�HZ��8X�;4X�7�p�.�p�輠OF+��I�����ϖ?�ƷV�
đ��������b�$ ߅��H��Kj��>��/
FL0IR����|�y�h�0�p���r��2��8i�~��n�zeRY�Ҷ3g��|��޾ݓ���2�媫����3H��d�i���7r'�����<>/��[�+�;hD�?s%&4��Й�� ��0$3��)�	{�z����s	�K.H�s�P�`ؕ^���Ýen�m�.��
�,nvҺ�0�H�lvF���7��d��H�/�����眳e�UoD����oX�`<���T�����_n/�F)^"c��K�ERs@�(�N^n��O��jA�h��`YVS6x@�wj�A�a������J׹g�71|O�xw��꛾��[����׻?���XwE��"
g<�-��(��^�>�gO)kg���v�w} 5��m��-�Rq��\ߔ��2�}��4$D���(E˫
6�8�MR�ɂZM��us)��ֺ,�&���ib�)�F�@\0/� �i����?j���>���'����JRsv,v���:�0D!�����j O蕉��&��$1xu�C�kq���#d�a�Ϝ\�Q��s�a���a�Q�a�B���J�>ϴ��;�l�O�_X9����k�]�{��6��8�O5Nl�yѩ
'��%oe�]�w�%��߽����#=�X���;I�&	�(3m �DԢ"��(��M�&�<���\�C��MR	|��|��m �&ʙ!�O�Q�Q8�y�vB�4�ʤz&͑|��%�+���1b}�H�Z�ݠJ�߀��{eI�z��a�x������f���;/Mn��;����g*����&9U&�Z�4���[ë�G?���ny�'�x�s���sf]�s�sH�0`�s�d��u(B�e2Gxi�r{R��ʥ��?�=��L�>�A�8X2���LP�%O����J�쉔��x4ญ����������*�{�!z�B^uU��_�=�s�����g�f����j �t$2��=���؇l�����%&D�( 2s:��·{'\�z1�}F����2+Nl�W\y��2fqO�ݛ+z��
��G[K���cf�w�3��]�R���Ss�0�D+$�z �9J��w��Z��W�L�k�b�~����|�l��4	h��2��U�}��v}�����v�s�x�O~"�]9�5C d�z�pT�_6��WgSkq,�aȂ��M�-ip��l�^�oey�?m=��{.��ȷ��N<z|o�D/c���Re��|��J��-_9����z���&^z)9�G74�g���,��ߡ�?KR�v����ȣC�������X\8��sR*9d�2M�V"��������M\M1E�{'�	=�J��'����:)�cJ�K�����t��ʁ�a܉O}����_h�{�t��[�\⺵=A�u/��X��x�^y,����G����+w �<N�=����yy�m�-mn���mA���c%�Ijm��w�v`j�M�A{�w{��kx��\OpAy�Wm��Qx�5P��!V��FHg�!&�8�!x+�ܟn��Gν���旿\Qp��������mz�u��w`�ܠ
��[N0���k<!7�96o"`�UP���
:��
����Efќ�Uښ'\MF��*�d	��QR6Ś�6e�S�����s��d��\��ǏEg~o���AևP�p�qQ�^�̅!%�V�za�l�"=w��.R�K��p!�*�(���2�%�vx-��L�P4�y��c��<�8o�MD�]�g���9r�5�w���%���;��b��+��<��zT�ɡ��������Kw�k�����@��|�q�2�g�.]��!��� ���@�+�-j�+L�f'&�!���8���$	���I̓ �K�{��i+z��v�`f����.0�q]��P��Ven�v_�7��7���E��_BX�u'd[�J���FTg{KS�o��-���_����P����.�?~c���ωN�%z�POy2�W������N�<.�p�r'�xbm�t&'��v?�j/Q�Wk��o�"�4��<?	�z�wrf����}���|��n�;����׿���o�e�/}���詟PA���hNM�˄4����N(�Dz/�b�)�`Ɖ������1��PO�L�tE.\0�C�R�P0�M���M'���K}���&ʍ8�V�T���ݹ/aџ����O�U��5���M_P-��U�ow�;K�E��:�Cd)��I�m|P��]��Q��1��fƑ�ʹ"�s� ���x���t{R��Y���)7��Ӈۿ_�г�,=�/U_�����P�[^��T�oxfA�gS��-���#_x��}o8�Ⱦ�����t:�e�LK����+� �	1�;κۚ�����R��(n��cc��y�= U��Ro~��J�m?R�,�\VͳH���jS��[�b�R�����JRYh���$
*d�֟
i5�-��E$�oy��c�]/�7�E��:�P=���H���N1�n��P���m��M�����aܬL5 �;�6S��*z$��^��Q�����⩲�h�	w'�h����L�`�cG��_p�x�C���ۯv��_������L�=���U�W�0775�z�6�`dDK��>��$�:�Ϳ�����|��b)�} ���i6-u�Ym��~��P���{�#�^�I�L�
D|�uo�:��o���\z-Ϳ�����Wݟ���ջ��N$(Jeh�k6���\���ތ��L�Q^4��R)�X"ҭ?G�q���w��Ҿ�AI�Bﺴ�il�:N�>�)̽i�0{��b�;���g�9߹҉�)KaⱲ["A��L,�;�Nq��R�U�7m}~�>��9��NBW���t]�JcV�1!��Iz}m�$�b�4�C�/xPEq�;�&0����+?����a��"Ѱ+W?�,XZmf��c��3 _�{���m�"@��/�ЩZ]mCCH�����8���C������Am?���D!u��q�S��2 8t�0=o�~�p�z\��G�<��|_pr�۳[����<�Y!�)q�4_����_�3��}b���zP��e.L�fg�������{�k��P�|r�nǚ|E:=d�����&n�I_����q�I��6��	�G�c}.�b� ��O�k��_�EVbԸ|���Qfb��m�b,<�T���5�i���_���W�+Y���!�0Pd��(���oM�1��<�O�����z�'Zt�!0�yK���n��21�EFAO��
�e�	X���U��K/ѻ]�ZVm�ur`ia�ys�V,睗��[����!���h�[�_'���1u�3� ��FB��\f딶�܃��t�a�E����2H��a{E1�`��Ct
��o��T�E���$�qHb�\����U����0�6̷2�Sa����?/��RG�(��၀����7�2�^��6L�v�8�Vw�����^�I�D��P��U�WCa`8�:[O���&���G�b�҈��[�y\~��-��cK�]�i"�y������������bM��r=����]dD{�z��4�m�0o�և�#����k[��P��}�y�u��0��Q��m�fX�5 <.N�o���/I�y�h�}�C��m�bϡ�K�+�6u 5P*d2lj�m��kĈk�+�F�`X\��c�0�#m�}��Z���:�UҶ�T��'v<�n0�,U�����Y� -�!i�b��5Rg^�p�f����KN�4Q�wl�=���C蓼B����������p2�;j��s.y�:���l4
���a���V2c�݋��"��?�y}d.�6��fDv����B��@�f�Jd�ف�������J@��@�m��%�Cׯ���{��l.�q0U�e���E!S���#g�0����Y68%s�LM4}^��Nq��5B��i�5s2��]�T��3�Q������(w���ge�go�^�-�(�֢���y�Cﺃ��?ւ��'*o
O�({]3�3뻰��1l?����cܱl�k��*r�A�O�G˴ E0e/�Zn6IEz,(W^�X�Jb���E�;-H~�Vj���N`�6�F3!xbz��B��bhA��v�W�M�\�g�Cq��Z�"�I�-�R�E���܄��f�� a�0&5 N	H?�OU�)�8C�� �j�ѸAΪ;�����o�R�
�ڀڣ�Nd�q��ԑ��4�q���0Ȓg�_�Y��$s̥(;���F!d�R*ƢQޅ��}ya�.��$��i`���^7�|rb%!�JM�㋋mR��i�R��Z) �VB��Ou@��ΗX%��/�(�(A��9��b<�
�>s���q�T02o���j���rYn��.��8GD:	�PF�R�܌��WM��j�9�ǜĴ��H��� |y!I���S��狭�TED/�;�
�~�Ԧ��h��o߉c�������1����\Q	�����N��.��o�C��u�OH�t��\�.�c���n��-���0��9�����z����M�������or%�Gy����5���FN-I�ǙRh��%�����4t�me,Z�-�OZS^�Ȫ�: U�r���~0��k�_�ae./B��P�å dB�Է�X���[JE��ō�42�Ȝ^dO
b2c�*�k"�f�6�����ʛ�"'�@�=��2>��	���L������I�Z��)�)�N�������#�C4��x��-0(Ւ�֩6���/��{�����[s�b*�$"�ѩ��kNn�c_!U��h��2�b� ���Z�\��V��a�ee��hW13��h�x[�p��Z��m?Z�{:�͜���*�w�HP4�p�p���t�6�qՍ�A6x#�	�6�փ�ض�D&I�t��3�k7��'�����t$d� 񍳹@�"�eJ�Ҥ�xν�>����/�o����w1������ӳ���s�>v����	�_�<w�ѣ8(����8���K�1����:X�r+���T�%�K*�����H�➓ǷCQ2p�+�3Z�M�ŉl�Ԙ(���c%[y�\<u��(Ԇ(�k�ȩh�r�	K�%:��,�#��U9CM֖;��q5_��0b���"�uQ��=�!�P�X:�Lת�[-�0����ͥ
Y�m2Ub�Ƥq s���;{!T�m��}�/*�rȷ� �*�4�������{������]W��ɒ��aҞ�Eh��d?^c��m��2+�懬�w��<Z�*�J\��Ԇ Bmb�v�VA�p]y��ؾe���]F��,���t�ԛ}pE��H@�x\@8l��c�e���:�������9o�+!���3Cb�EPF��3c��oYP�p	½3w�� �d�5+�zf��W�p��
�H���-[.��_�P^�����O6��ݴc۫�+��d�e�SFXr�A-�J�z{�Յ0N��@�#'�+Q��;(%e�	<���jǉ]c�Im�6�@���&�D�ˉ��E3*$K��~Z_˲L>�K��u[i�V�P��c`���!�a쩣��ǆ�_ڞjq��-���^(��"�tPӻA�y�!7^�����<��I�~�ę1�_9�4�>B�q�ML���0[�bT�%�1�vH��o|Q�W�TH� C��4E�
^8�\���~�V�rY�'�e�j}�l�ԧ-iF�vvE_����K�L���K�;m�z.�1�w"ٹY6���o�Ԧ����r曷$/Xh���+e2�,`�m�LiLD�B����V��E�	rXv�w�N)�kc)�����uDB�"��g4���6o��Ȼ�����3~��~����Pڎ:�\j�Ci�շ�ඟ^v��|p�k~�������WBI�1|��ۇf�i����и�8���0�"�a�_�F'tH�	:ԟ�巩��^�w��1�A��b�TI�hB�Z1YVc���+�TIG�O�	O���(͍SK�G�m��e�_��,F���B�X�2�/�SrA5����5Pͧ=	������f�>?y�ܾԊ�������|e�b���Z�2=����y�!����K�mN^��u�+�'d�
�� l)��Qg�ݟ@��@�X�e����l��\A��QA�@u�j<k�V�_���P�x������ց����;w�Oݕ<J���&g>xh�F���eR��x��&�D�[�j��K��p�^�l뎭;���2��4U�V[�*��ҝIMN�[w�FZ29��y��7}�(�������3�l�(/���61и�͕�������>���C��fY/c�8��x�{�ے�LpG�����|9gB�I&�L����-`���)�U�]ZK���ի�H۵��ҶL�B-���%P"ʠ�/!�Lrz/3��7�ӝ�ѱwD���s��/�ʎ���{��ĉ��������}�����7��/l˘h^��u�����ط���<k;����XB��']�LT�1�M#y�J^I
��ɱH6�`��:ϓڶ�����f̖l"�df�o��'�Fg&d�1�(��N�`\RӌB_�FIH�v��Y���a���&�5�8�ƱS�O��F�Er������?���}��H��_���p�K	W��g>���JjΧJ��|�yf;��n簪뱒4��z��VWfy
s%5�XxX�[�p���-�G�P�BCM��LV#��P(�# TF�$���ev����_��z"��2�������?�S���ޭ�.��ou_>(��\~�n�IE�rE�04),=%����x`����|�(�$bE�\t�9��N���J��0�ų�J#�i�I���\;CxU����U/��調>8}0��_[����a�<�v�57�����p��������%q!�ٚg�M��,8h��+.)��.�\1?�U�T[���ھ����vd�)������k�|h$��!�l�<z��`b*�ORG�[_��Z�Rj�;��l�=�a�h�	t���ڐ+<����m22�����	9�F#qh3z�g�_9�	����.��j�����>gPB��b��=N��)9o�;wX����,+u��62�FC��@68?��8Ip�|��`Lo������D�6�7��J���4����u?��� ���c�#��SR��^ȣ��~��T��n^��<�s�M/*P��"�C���dx��9�s�\A���ݶ@�f��"��j�1���@�G����d��K��}�]uÓdQ����hT�;���C�c�,�݅�U�l�eW���K�'�aw�u�C��y�w�����w=�^�k��:�������T�+"��A�;�MF�!	ڃ*��./�z+�0CH����8��r�^�Z�	�_���G�X ���yFzז�R3`��X�6�\I�d����>��VB���3g�P�i'+~+��Q���q�F��9]8^��õF,� ��	��N��s�y�ÿ����_|Uv��?o�R�׿v���>2�1�(�����nos�0~-�Bi'Z���I��.���	�d���v7D?���I�)�A���xo�}�|���z~	�>��8L^��'F��"{�0�ڭk�_�£�q��n���>y�5��K���ko]�&og�ڧ��9����T�6x�|2�^n��I�g�@�j�1���y������q _����G�u%ϟ~ts3�[[t�`5��=`�k�M/|�_����9:s�g��<�)��k��w5����80�&0��+Ӭ�h�mK�Η���e>hSDD�Nʽ�� ��^Vb�)�zRԮ�^�U@m�"x.7�Z�)ʐ� $I���Y�h��,��uB�Q.1~�âqnr��NV���	)����c�8�Nz���V��f����|�����M��ϸ����XI�tYd�B��a���o����}\@)�����қh7�!�J�fY��R;�n���[��m�i;^Sϡ~�(➫	zdO�%ڌ� {�
[1Y�v@%'�$WZ;��d���v原v�O�����{+��wM����B��b�ߖ{�c����,`+Y^����K�|?<q�ƛ����N<n<��'�3wߓ�Od���%�� /��Ccs���ѯ���e�$|��ݘ ��� x,�j�R���dBO�e�Ib�:�G�}3��������yN���=o��u�G��g��⭓B����d&��z꭯��'�������G:-�@��cP�~>�Pz���a�SH�2��i�\�ޚe)I��lL_�2�(�#U������tu^�:UtU�e�*��ѹ�9��3�$�yK�N�3fb�-c���V豢-���E���RqS��g�14Bs�$���@��ΰP��Mh`I�����q��odQ�k���W�M���)d��=�N<QcY��@c���3Ғ�zE��X(�g�n��v�g�-H����԰��P�Z�}%3�U�-� ������s��W?^�k�/�W^8R]��W������х�:6>O\��/c�mKQ3L3^D��D�>7�,-��w~�q4�ی$�Ԡ���IRQv��}$�%�8�
η.�YQ�k(�\]:�:8�L�ɕ�ncG�a��Kk�e�%Ļ�,��Qn2�v�q�;)�����!���*�����쉟��{��+�O��U����ăcB�\��;sm<�*� K�&��l@G0"q"�JVJ�m��L���M�J�W`�V��[D�	v{���m@�"T3`�F���Û��Z��������g��R1�o~�L�=��M�C5���d^��e���N?�{^I��W����}s���,ϟ�1 ����YI ���8�h�eLq���iƒ-F�O��L�X���(���Y���
gS�/�,��e��7V��$�i"d�`l��;@6�Xo�Ul�	bU�9NV�%VĬ�{1x�QV��S+Ɋ�|��#s#�ˍ���Q��#�3��f�m�A����,	Y��<�zУ�=;�m�M^+Q �L-:�>6�v0[�݆,��͈\���zڭ�>��!}�/�����?6�7����\_Y%�;vl�����a�b�wWzV��*�F9���k�������;���;[m˪xD��Z��Vo����j4*F/<����Z�V<)_��p����\<��&��E|�B�[�
�+%_�Fb�"��j�?�9��'O��O�U�����x~��х5�Q���5aa����a����V\Z"-pq���rm��r�JO@2�!��� �E��+?~�y߼���p���+^��O|���/���3ꩾ>]�����I�����7���[���;s���a��3�wQ�K�3�+e~אR���r�����0�
����Z�"��Em�	�0�3�f�5�<�����t�ҍ�'7wV���0I8�%�$���X��{Z�d�X�<�2;-�$�G�!6n�R�B�yR#��u�Mb���L�TMx�ז�#R��UV�"Di��O�V]�Ƶq�����{��ܯ��[�����;ȿ��y�Z�j�����#׮��>���=S6Q����;4����r�<)�2��:�C�`xz�~���~���0�q]�A��i��KDk�1E���{��k��B1yFׄSD���$Is�}{�Rnԡ�������"j��1��.���#'��ӯ����<z�����Z 8B��KxY3ɤ�G�.�(���I1Fg�)W��&�N(	8���n����s/�Z�)��H/�#?�щw�+�m�a�SQ�����㫫�/��<g�67��;!z�ސ����ȑQ�_�����6�<K/{es�[�1_�����K�1���D�>D�_tk�Q2��q�h���4TZN���Ji�h���}b���"��~=`�a�0O��J�[�r���%H�ED.j�YI��l�d��������e�iɒ�lc�UV���X�89��D=�gl0�([3�)�����C_I=�>��~����������w�����?��?��*�M2��FBNe�[���7־|�Bh-D�WY���B��ڡN�������^򙲜����l�䢎u>0L����o#C�}^��l=V{2����Z�Όj>��J�� a���Ba�3�e���{�WPI��Qo�{��nRd���C�,�nu�+��,��l�+>�W2�&4�R-��Qp�=6�L���z��Ʈ&"ZRz�V������=�?��?��~c��W^�xv�c,=�C�rG�����>��D���N�Ů=�����y���ߘ�����}����ܓ�?�m�5�)-=� �W>�F�`�Tf�R���/ٗq!�n�L��0h�	=F�pf� �Bz�����伱�E�Օ�=*^���.�崾���d�4&?�4���v�W��s'����fB�,u���h�)<>Q�ax�7f0IET0Π�px×"+�r�On�gx�f�w�����Ge���@�
x�½�����0P���r>3��
�d�z+��3�?�����YїW�wY�Cḑ2��V6u zy(LtB��D�j�:�%��!z����ƌ�}�<��e�v��sB�l)EjPfm?�d\�����mtWB_�s��cNm\/��e����{5�d��%s�Ī�kw��E&�a֊Vx��{�m����������v��V!e�Pd#��-Cؒ��l���x�<�:v4G�)I��p���wj��#;|�h'緩�1:Gv�
6���]�ª獈xʈ�X�o��$[�#7G9�}f���軁��Sc��snV\mSt��MƶS}�U�RB��w�*�1��f��E�I��t��C�<$~��\�5�vT�=Y��I;7�T��)]�D=/J���v����mn���?�������[�����O��+�֡��Oot���2Lr� \9P��
��TtI¤ŵ��2��s	� ���e�}(Ip�*Rz/���
(>ʚ[��Ԧ�{�a���իh�9s��1l ����Ŵ�tN��	q��;�W�Aq4�K0�S!+�@��k�Z%��Q����F�e���B+^LΟ���MF$M�+!��D×���Ҝb��^�2|��P�P��ՍG���m�}������~�P��U7���[ۭ�`Z�C����?V�w!WK���9b���:GV^����	�'�}���a�A?�Y+ha��n�|9�������J�J,a���-s�ˉ@_\���B��Aq142��.%@���Q����ki}�;��fZ�f�'��Lv}����';�mm�(�K���Kn(�_e�^~3���P.�hZ�R����$]"�k�0�8U�B+WO�a�(�[�lW�|x�����zR��w����������>�w��l㍻yz{��/(��}�Qo��B��܄WR˪rC�c)��5w�}�ʺǵ�MiR��-:+�s����D�e�zxSy�s�f75�n��=J���'�߆��4�Ad�w�(,���#�5#�0���aU�v�/�x�o�)�/�B6�<g�:���Y,��m>����4?{�Q���e�oJ�#��n�\_��2h����~i���.~�g_�y��� <kt�\������#����� KH�M�Z�8S�v�3��cA�pC���^q��c��M<��~u�P��to7������J5V�JK�".W4\����I��XP��~����6��Ƅ�c��˒y�����<g0�����&:i���2�>�i��zQ��3�gp��E^�u��(�0�C6�d
�|Ҙ���&����N�g�[hz���4�د�2�q�5��K]����3��Ŀ��#�E�/>t��}�߿����A|�ןP��ڛ��ܡ�[�O��,�7څvҸgyAҵ�6��2�4�}���g�Cra�_��:A�	~n%���=��$QZ^�o��c����Tᷬ��F�F)�_�*&6t��Bf蟆2Т�@<�S��C���j�s�\	�ZA� W��d�7���Mu߫�xN� �zē���;s�j&�w�٬�v��xK(�(?��6�7�0�0�g�����j��o��zx����<9�o��*���/T�Jv���D}6��ۇVQr��x��{o���cp����I�D �ߢ�+@�-���\E�1րZt��R�g!����$��N�K�MQ�ezN�4��0�D��1Ӕ����Or?���X����<Y��&��+M|�v��u3��d���vn���c%R-3
e0�c��S��F-C&)*�x�Z�=D{�(�Ɵaܦ[���Z�6��y9%�:%�u�z��vURm�<f���0�bhwW�,W�{��c�k̴���P����7����%��	�x�ԷE��Ⱦ�-!�`]�<?b0L�p#W�<Eh7|�zu��(㸀�0�rA���)�[�_m���*�+��-�����b`6v9��PYY0_��2�u�J3~@���@��~L��mQD|5q��4"_c��#u^��!O�E>S�3$TGcm�j.g)����P�4�G�|7
�������3�BJ_���2���av�R�>/�EyW��X�<;�5�g5�8��=w{u���;����z�����r�N��d�0 o�������^����ޖ?���]�Zߙ���ƾ)%��]	#�zMG�YՄU� ~H]Sɚ�H^'�m�����Ub}��_����u��8*E�0�pQ����:��+�NV����axv�\U);��Kwya�������!�����',��N��~���~�<��A_���َ�ׂ��d��%�/����&����'���/O�����8�Ш@s�i|�vh�)�&LĀؤ���pU�e�c�_��qθN3av�dÌ��惖>Q)G�,%�:!��8�
�b����F��;>���^�ҏ�{�_�e�x��|şV#�n#�$ s�h�������F�T��O�k;��3�����ŝn�zʋ%����?�/�'&@M���((N�y�ꥃm�D
E��x�c�@,#<�`�qޗ��B�He¹�U�}5�A�z/OvU��]E�=����j�]�Y�^&˶�kG�\n������G�r�y�� >��'��#��gpC���Z�F�S�,&}�oNC;$�CI6���^�H}��wE)<�O<1��b���
+����ϸ�{7�zW_�uW�ſ��wo�%,˴CA��Ċ!T���"�Cd��Zg-�����f���/�����A�������J��BM�R�����e\(�7+�MM��6�4�����c<	���\��� :���[`#�l�9�-��&��6��q��	�B�`�-~σ6�i@��*I�ɋ}�=uY=� E[,�;��/\,$�:]C"��T�c��sZQ~q�����N��9c��}��k�_���톆���)��L��^β2Rtg�R���54<�����4z�V�=��J#DZD�[�������6���SA'�1�VTǻ�p���n\%e�� ��ڔ�I��Ӿ��H��É�-��Z& ��1��{>(�F���6�\�7	�:���n�2�cY���#G6��Y��Û�WnyƱ���l6x�[�w�_ȣ_���u^q��BI~���S����E��O��3�Y�6O=L��/3�19��b����_�ۜS�}���/�lj�����M�ɯ���x��_���$91�Y��9-��0�~�(M�yek�2��e/�C�-�|��Ȼ�>��}���{vΞ�R+d�Od0��.�#��vE���q�Y���&Ȯ�ju�h4��a�TX"����V�0��" ����Lv��̓Ɠ��m���/ ��Z$�����3U�t�،,����w�аMbv��Nٺ_3DxItqT����JE	~<P����W�HD!v�<��#F;&�-]��ݘ]p�˳��cu��u��?��g�è�eR��)(�������[[!84�����~��XF����B8�&1fJ��"��S1e6#l˚�7ױ�i0��N=r��n�E���m����[O�c�\�>��$	�3�M�KL�SJ��Ar�3C����O����8}ko���[���[p]�@���d� +r�e3	w�O?�����Jt�B����,qɕ��r��c�}L�h���ą��R��s�;�K�{�?Ԓ�V��2�I�b���]_TvxR�8����F,��љ'�i�)��V��V�(d��v����!\�Fdjo�	*аxr�����W&~�f�{�s��r���h�x����#�ϊ�Sn���F�V��$�L��;e&ˤ���te%y�u�ԻF����/���O�q5?:��L����C�8v��j*,?������ �<![�uR���,uWh�m�(�c�r�^�>�	�_8%c<��j�wV}_Q���k�� ��·�}���O��Nݧ�j!��C
�g"��?�+�6�~ݑ��߃U%.����N��?���3/�+�#�����b�P��yR�����D�P������v�W�Q����๲�����n�K7����od���u�˕G�ky���r�Չ�y�����k/E�_�7md2Y�pE3�@i^b��L��|��1_�Ӹz��3��V���'{{�׿���#��?��tR��ro��j�aqB���g"�L��8[e քE|"B	ʠ�)��k��~���]���}�k�AH�X�j#�y�B�W�i���l��Q��HZ�]�����'��m��}JJWR|v�\�։�D���6�l�tᠽ��k(��@&��/tM�:D�(���������~�o$��BC��U�@[�T�/a�t�N��sm�m_1	T���/����/�H�8)���]tn�_�_�߱��{bEY(��I�Y�XΔĢtOF��"�$IA!,>h���#��/"Ų�Q2�H$a�eKm]�;v綱l������ny:`4ѐ`�0R$qՕ"�9W�j�Rs�/7��3�*��PJ�u{��a�҃���v��	�?����<?�w���zw����Y6� ��V�K�O�u&�������7�ޖJ���a�a[ p��.�vֈ�����Y�0��[��)3,)5I�d.\���̩�aԠľ�,9������j��O~�������(�1��ܨ���bE�[@uU�A6m��̂ ��c�.2`�rp?ֹ����g��_��v�����d9��+j�%i��V��+��hq���������Sm��n����������%�hZ�1�2���}X��X�R�A���y��x�=֐ix�Kؒl�3R���>l*����%/J�~-Y2@���-L�!�����ؿ9�2/Ӑ��$!���E6xI�S������ְ��H��UF����\t�Hig
�q�/L�F��@�����R����#JZ�E)![��Ha�}H�b�X|��"�Sr�����8Ψ핊�l��!�����Ń�{/���q{�!5L���c&1S��Үj�0�eL;���DL�q��b�i/9�g�H���vv�TI1Y�{y����`�|����4̋��FK�ȶ���a��q>B2R��7��
C���<A;<�ɵ9�O���݅� [�s�$��m�ř@`|����zS_#r���'ıd��'h�i+�w�,J��JX�
1�1�]�X�;0����PL���{�����N?�ߙ%��� -���1I�&��&/;������M�`��f7��L��#�/������7[]Z�$U�=��R�\��aV��E�,0�YHK�mҢ%�Jj',q� N�˩R12SC��e_�[n�b�+yB�]�>� ��L������5L�����PQ26�C8���am*���B�Q$�g�����;W�Y��Ӹ��a�3M���$P/��!�z)t,@b^@�ow��;�E������(O���'�ʥz����ơR,)�B�W�B�����:���I`4Z/������w*o���d�!lRDc�P#�Ԝ�+!������"E�|C�\�h]Q�\���/���h`B'� �cq�p�l�A�]_�UfL1�S�#u�K4+	U�I�Xo��ū�hV ����
�z�+/�����+��u9�C�g���Yjhdt ���I�5��5'���$��4̋J�g�!v5�������Do�:��V��X�d{1���Ei
5�J5���U�ʱ~������UK��M��o��x�������T�VJ�j�Ah��'{8��ϖ@�q�p>��(�QAXRUg7;�1���e��#_��d���^Mǵ�j���\�� �D[a�e�0R �院���T�ƊF�LWRB������"
�����eh�y��IBA�_���8P�6�i���F
��+�����i[-�ߐg�3�X�3=�"H�ҜG�0�v��K�ϮE~=qrd��Z\9�鉔)�K�	%��:�0��ªl�&L^�4��^�
x���q
�|D��s���S���lr��6N)�S�2,ЇZ"2>t���T�
�u(u	q*12�uM
S�(`�3�QѤ��h|~K��r�N��c�Nj߈:y�E&Я��V_Dh��|�;3�P�R�M��B��J ^*�Rz��Z�P�^�Ydf���	�N�f�3Vm��>��Z	a�ț�6/	�5�	s[f�`u�G� �
��)衵��H�=5�\1Ք�[��2C"Kjs[��h�t��%�`��<�9N}����0�X�y�3�Y�WW���2.%C�J����W��0�м*|]T5c^A�{�G۷�L�{!�h�[9
	R�����あ� ��Jb ����J�Ou�����j����~n�ݧ9	5<���+�c_[u|^��^�m&���l��އ�b:�ς%�IY:;޺��M��ڠ�Ț�T3l�`���`�1����>�0����'|�g��ewr�t.sҿ�8�jnj�e���Ď�D�����1�TIL!��W�Ʈ=�E	o(s�|��L�AN��0R��@�t��ʐ�#f=��%�6�������7��g���j��qBK�^�0I�ݦ�d(��W��*0��F#*+�	���E� ]�ڂE�4DJM�Hq�Ki
�}$���~�'����Rb�~
�,^$gZ�A�Jy".|2�p�y�oa��b�2
�v.� 0�q8�eSc��bb<]�N���<�������%E���X_1 9��E�ľɆ�K#t�#h��D�Y�_�f<�w��(a��X��ω��a**1&+�ʩV�D�n��Bi�X6�h���"<xp�Xn�'���c��Jn��>�ig�R���>��2��Ŧ���׫ƈ������ᗦ��%�e�g�?��R=���G�D4\���3x((� �©�Mm�A\;>��4�ތG�l�Xy�Nu��B���IGJr�[��$�u�Yy�M�ߦ��4�#���"�  �ԯ����t>C��g@N=�&���1��Sq,�f�Kh+�嘑j�~���d��څm$��]Y��7�ZI��sq����m�B�.B��I�RҹzZz���ӆ3�d�� s�ŉhA��i��$4�7R����+��̠MA�"<��	c��4zE�]J}	�3��*���f��>��g��7@֦Bm�t��C!#��s>b��D,�����3	��π����a�Tw�Y\vO�CO��K�Ͳ"���\��7���$��sMX�'37mb��x�l�G౤ͨ��x�5�ˋ�K��ϗs@b8H�J�e�����5NN��KD��0Ŧ@g�G𬒾�jN��&W�J�}D�XcU�����l��+b7���t����M�F3�أ��
N#S�19�	:�z�$O��b�#��U��r8�	�Gs��Z�/�2���I6�a=H��ҳl�~��M�s������L'�&���$�l8��G��nD�#:R49�v%���UA6#Q̩Ĥ%q*h:��[X�w��\�8��1���ZC���l�|n"�������{�:���3Z���#�4 �Eh��Q+����)�������qN���m;��|��p���$�j��/��a����_~�V"�x�-�F�IY��EmF.��%�qqɾ*\��<]���	��Q���P��Q}2I�ڒ���H4ѕ4��y��qIX���Ǭ&�x7��%�ym�1�0�R��'��75|��l1DcU[�o�]�;�ka�cZ������+s����./�UN4�r�=¤�,"�������/�%�	��gr|�ѳ1]�U��#�:C�;oy:��'��c@]�@uo� ��+��h�Ԕ<�J����(��`�V9'�T#��4��Eq�0>o���~�ƫ�l=�f�C:��L�����Z��И��� �Ӓ@�C�+4�/��+}�!�0)�0�3M��+��u57�C�Z�L�ː/�����ڲ ��<|"� 2��
2�k��x��R&�E&x;���Q�
2�'��D'E�=c}�f�k^\L8)�6�`���>��6����ڸ��=����}Q�h�;�d"w�H��u7�M�B���,���J�ऍ�F��:���:4�00�Xf#ࡺ#�!\��]��|�ʳF�)5��� w�]>�i��L�D�?m��(@�[����pU&�	�k6�U�v;�+����厡t.(�#L���o�����@'�J��w�ҚB/�[-)�N���9c�7�O�}��<��)1��:B��P�=LtB(22�ؽ�(1c�z%-#����in?���T-�zJ�'�-����$��=���A��|%I�Ѫ,|�8)��i��z���|yY~R.���hؒ�@i���WVtU�y�Y�b�IO��� �R�u�<ڡ�Ԅ�hFEeE����RJ�&{F�ci�D8pR�b�3�p����26�[�w��Zt�x�g:8GM�\I����8�7�qnYq@�0F�ӅX��|�%��H�qm+��-l�MNaZ�0R1[{z�s�m�\0>��Ǚ�H���t67`��,���
�kL��1U�3+A�����K���>�_�>�*��8�f���,���Y�5���uk�
ǤqmNt%y@J5�-;A��e+���c�i���l�7l�6gz=퀗4���Di��\rćt�Œ{ᐳHp�R�aD�zg�ݢHnl,��9����'�o�)�매`#�Q��(����V�F��u=��|Ţh��\4I$�����ě�D��	���K05���bz�t� �܊PP���
�|M,�g�z�Ձ=����h��|Q_3�t���0m�uI���Faj�b���>�2S��((ԧIK'I��:��I��"J񴨈��8F�sM\���#MG���jIzzU��;��[����ߝ���$���H��������υ���� Za0�	�L�����fa:��Q,1P�� R�4����Pn�Ff�5��ڻ7V��nM�h�ZS"���fv�"4��98����Z)6U�Ə�X����d��i^�-�~13��H�w߼� �(b��+�Rc
�(j��e�ʜ)��4� �aN�i�&�(B��`[�)+/t�_i*��0Q4������'�H&+��AP6��>�\G��!�L��B�`I>T��~؁���8Q�cGG��!�%r$�86���Y��O�H�8���H2�hJ8�Cfr���8l�9��-0D���Jh���t$�t��rm-Y��c/Վ^����eE*�5�2�J��DѠ-���tJ�4Б�:�ˌa�s��xv_-:E�G��v<����3����"i"c�E?h
��J�0�g1y
����� ̸�̾I�9��-#�Z9�(��D�Xw���,�
���=]dc�s�(��\��Z&?c�R���T�7�[�H����d�"Е�}տ<U�8�$�ig�M�E�9	!����U��l�13�IB[�N0[�`���z���\V���i��Yr�θ&({��#U���O^*���ZIV�B��;�?0q�a�b�i�VhĻ���bRK�aufb�#���gEE}r�ʈ�?�Ť)���ߥ��M���%����]���ir��>2��W(B��@�d�
�R�F��̻��*������d���"<!�b�]����r���	�S��͂Cv4�Gf�&7S��N+�����Fj@y� -��(.X$��o�v�Rj�`�~�)k��Z��H-��Bf�:����~�ii��˪B	Sk_1�6!�aRK�6it���I�p~����8Lo�?��q�D.�j�^��3�6�T�MG�"�Zb3�$X�4S"���W�����&~���o$)M�R���湙G�<�M%'&�h��8;^�O�@��z)M��k�j��Z*�+��er�3�J�({�4j�5��.y��$C�b�$0����3Nk,5�s���%�D�C%nX ZQ�&����h���ԲU��1C"&��ĝEH�6�'��)-�;U��$5��o4h���<��c����KC� ����@5���E|����hjp˴�+ӏz{%j�X3�eD#)�Y�(39l��%)�,����0�W�d$�h��G�T�RV�I� �\�>���~�me.t~'�`M��1o�8�������Z��ra0�e�^�f^'��Nf*�9�\���i�M,n�h���j���x7�~R� )y�����n���}�����љ�~+�=šB�)�+A'��= V�l��H�5Q��kn�!8Z�?�:qu�����pǿ�u��n��w��'G���f�V[I���K��[BҁH�V~�
��eM�<��s��z{۽��`�x���\13�:�j�TR��vЄ3�uH�d������D�*����G6~l9|��?c�ޢ`T���&�[P�ײ@p:��}^(M���Χï�G�w�:T= �i�Z��,˄�ٞ,v��`]�?R��'��@�M�C6���UX+��i����>�@w�]��;>6oc�V��Hu�ݴ����fK�4E�Ŕ\Yd����BN*����iZ��%+� P��J���2� <�%v�B�g���W��m�\fsU\&�Z�dI���2�s|�jc�Y�}lM$�d���n����&%߶�v�1?�15��4kN�%��/�yXE�q�KH
�Ǡ���*�M��7�w�����W�z$�}�W�G��rs$n(�I��ң2reR
2����d.�$T�cF���+9I��`���y�(C$QZ��3I��U�ms5�[�U��~��*�d�4KߙA���h��ǡW�=U]���Wl���7>����������Y�*�1�n&��Ao��n�|���2��&Lh��3��t�GF�$����h\�sBK�����m���40���36j�)��Wi�01n�{�~���K�Ef�Es�ڹ����sO��{�$�^*,;�Ak`2����׿�=p&�p��Ɂ���Q��H�#h03�)4��1��������m�2�d�Sm��X��2Vk�w�:��!b2��&��> 3�pR�!��G�q��}N �D\�.��ì�W�Yr�l��}��?���[��o��}}\�:p��{E-�}��PU;{�sL|_������Y+��c)�rsVn�v�Rȿ�_�c��v���W)ܹ��0�U_F&���7ݖ��_@�].�h��,��$J�i,O��ޥ�[v��V�����|㹇ZW����v��o�ݥ�ҞǸ&�`S���j'��S�!�N�ը�цjl���
�	�3S~�3"���ƶ,%��R�����qa W����Nd����LOv���I98��k-�,����KO�=(�?���>w<;��+}�qB1a`��l�h=Y^-z�m4�xO������~�:�g)镊����Xhۮ��MV#���V����)j�5f�8��w0ω�Ra=��X8� 7V����Y>6N8���)4�b�߼w?�y(���D��?��مG������o�}���p�k��'���"�z���H;����W�,����RPZ�ԻRQY秒�'m�8�C���a*JH�Vm��9N��q���Gz?mA?���o:��j��'���/�s��ڱi������3��s[�߹F�� @�?, �������?y*L�f5�/;���!�h�j�����A�Z�(��Rj��&B�&��2O��Ϗ�GJ�@z�8��5�̊�<j��|n�3�;QD�6`Њ�<:~�?1H�m$�z�����#����E��|��H�S�I�hp�s���{�9��׽:�t�H��=�M���zY��uG���+Q0g9+�'�I�+XA�v�O��hmF��p�0��N�ct4Nt%��ncH�	��G�%���[����c��RK�J?���~�Q���X����-Th�(֯�%M���[��`<�i�B�}�T�O��
.G��'��|�wGO�8͆��g��+�d��)?����q5Z-/��p��c�(z�k����߆W��w%��׭�u�dA�dd�T���+�� N�G��KD4�PQF2��{>�X�h��ƴ��!�H߅�=�[x3�o�1�X�
C0t"�2J�~�#!�q&^�^���M�{��h#=�lQ�	x�^uc,F�����'vv���ҙ������'��ǊB��0�^9tI`(D���s�ݿ���}�g�����t�e�]U� 
Ct`
"���1#��>\30�a0%g!�ep/E�0c:�QUL�mnсrV�w�h�#�y�z6�(�]�P�Ʒ�Z���Ef��m'�Լ%<��}�㽕X&/M��w�D�64����FF�P���������kQ!ߟ���V~N���y�&���>�W���B�~���I�&.��(�0jh��ě���ua�63�����;��L�0K׻�8+�{K���k�B�f � �6�"S%�9O�I^fg,ѮH�ic#�&A`3r�8�){�������DbKɜ_��?�W}8n_�h8�m���XM�!���@FJ=PD�+V���)��6D�qő�=;������y��ӮZ�R������G���U��D���$������7|�;B1�P)��)ZkyBl��c�}�s�d �~���z�1c�Eb����Q+j�త�m(���޷���>2H_%���������o�=y��Y��б�RT�ܴf�Q4�}�E�'ٛ�G�שּ䓝#7��Z��A�8n�q?@[_ZJ��$�>ce�F��y�x�Q�)ib��ƭ��m�@�(1x��cF��Z����j�c�s�xի�A���\Q�D��Hq���oP�Rz,�O��(r1D_�����!E�X̺b�(�q�a1侢��z���}x�<�T�S>qYP�j:mm���w�����.>Td��yS8����Ǐ�-�r��.*
�b^��}������a𨈯���������<�-����Y2��'�KGfb� �'���Lpf��,�<�~%��d>m�������QQ )V�җfᔆ����ir�HH��$��h�51ݪ>
���i�������l��c���{�K��}���p�:�Ja(�7E�N����[���]�m���|}'b�Ǳ���ë�O�y�j��{�Nu^.s�`@K��������)��:lW�9��2����y���}D��܏3�Q)�����7�oԙMH�D^"��h���l�����=v������3���a)u%cjT'q�w�T�D�� %���$�_�/�0I�m�rƱ��W��.�~��'�u����CGo�D�m~!_{���`�x��ȋXK��>Pn���Q�%�yi$�^�Ʈ��0��@`�uV�B��B����ȏd�T�=��%�2���V0(����(��I?~���W�e��M*S�
Y(G^�(_�K���B��꾁L<h�s��z�k�.���E�Z�_�p�1��/���HI2�,�\�ج,�v��H{��p�Ƞ����'��z�yj^�����6w�z���K�����&�w|�?��f���@k�Ag�\�1�z0���<	G��@Q����a"�P�cy� �9!˔R�J̊%����gOFà~����y�+�j�B��\i+�W&:�p���W���s�4.|%����!^��U�%0^<E�ò���y����=Vc��=�<�|����
?�>Js�����K흋��/�^�]:�����I�`�,��{	Z�1��n��+��n����x5�����/2�uM{u���8K�|�6�[�"B��R���"� JVЫ�.&��\�[�Q��H�I3�ԑ���eY�Eu*2�(�J��-����}�T���D&=,��y��,��uN`�>	^��O������O�}��/By���n���Gʽ��Rwk�X��{��<�{,-��]ȳ;����b���������E<V|8�"'���C�ҁ�vJm�+��7�����7�3Y،m�0��3�����̽X`�Q���H����3����C�\9b�^��y	�7����o�Retc&��X� �{b�v����(����S�!���^���F�("�W7�NV�hm�4�B�;�������z�����m�8�trWQ�b��}�hJ&���x�_�H�4����^�u��D��. ՗�8v0�8=�^U9��ى_{�!�}-�>U8�c�r��-�/���Q@9�� 6�*k����t��D��MJ��JQ;�4�Ң�F�(󼴗\��N�z��?;�}�;�_�q/��n3?wco��@�JthrY��ʱ�)/�`��g̢��������8�_�y>���s�ʜ*5Ճ�T�=��}X�ւ�$�T�kBE�<��LNdV���2cy�p:�==��y�h��`����~�]6Ufh�������n�������[���VF�}����tم��`�k��;�i�7- w��6���+�7=hl���lb����.1���Y�lk� �{�mVP>�&�]�����!UBPʎ����������zK�ߺC�-Q�J�R87��X�֔���3^y� �o������(��_���mA;(h����`�H'��i����<���ѫo��-��<j��hEȍ���w�X&��:�<u��n�a���(���E���W�d�T[�@T:�Rt���@�W�@�q,l���|�8,і�����9��U�:��`	K��4�ޥ#�l�|��M���2��*m�$�j�(����cD���4�!��HG�H��U�����yIV�CU�z�@��V{�'�`�z*W��JѢ)HI0�`�Υv()��Pk\�˼8&Ӵ�f���!P�o�Y�l�ɶ�ܴ�l^x��J���ØF���GU?��Ҕ�&�-�2���Y�JE�j<ǦÂyV���6�6��A��?� *�M��PE�y�S�y���,?e�"�R(�'���D��(�wisP�/�ӽ#�s�ţ�͇à5 /�x�@yQ4@���3�1�*2�j\wVo {�w�Չk�l[���z��=��d~ӏQ:�[coT��nF%yy�WC�r����
k�VYSk �":�p�Xo��[[o/{�OWwkIw�����u?,�d* ܖ�A�~���;Q����`��G��^������&���-7%��4-ߜWX�3S��
{�%>���J'�8���-�B}Y���,3Z�6��:�r����w)N�悲��?���4��X�'���w��L�����¶��
�)C��JN|�N:���g� ������� 䩳�kSui�6�:��`q#_�!.��K��j҃g0���(a�����06��^��@�]*���)����	h���Lg�L�+��D��H`r����9�:w�����JDa�b;h�K�����i��P��؛�Ft�0K�\[���[�����
k���ͨ���q`�1g��E�GJ�����a��ķ��to��}=��`YV�g�C�_W�ϺʨT�<���?i��ڕn�r	�c�K����N��f�<p��H��ʔ�):Nݔ�a�~_H�ɧQ���o��b�f���/L;jo����/�9��[��i���}Ne'�,g�":H�����K#����V���f��D,�GԷ�$��h��M�&LCS�xu-SG|2��6+9al�{f�ފ�9x)K5���"B�,S/����[�R�|{��<V�G3�9w*aM	 N��)��{:�<��1�����aV�f������s�q����3���>i���|�qd�w��;��&�(�d�c����j�<��<y�,�����x��d������%q����!��m8L>��Kե�f�F_�FA�F�ub�u� fP�u*�USwg��^ҝvr X�}�s��c�69蚳��IO��ײM.��=l�N��������52�[_�e
��ϥ?l��c��h's/ ���2[�3-9Uw/���
Xz��g3Y��̻�4c''w,�~V�����0YO�M��
����mm�;�9֖�ac�y|���<��4 \��M7ŋ��F��Rz˲6��m��9��66ȓ�}B���gY�YH�%4H�2/�9T���u<�t"��k�}]�R?��Jp��f"kU�����Xb�_m�,\-��o5ͤs���5�`N�̊��3���{9��DMqíYN�sb�{��}?����*���܊������q�Č<㍡�P��b<��֢N2`OO�")����&�am��z̛��1Lѿ�zn�q�~O�[{�e�_��v9�1xc����������L�	9����P)g�C���|x��ә��ls�xrN���6��q�Qi�i����b�4�=�*�m�eS��)a�3w���q�ݺ�W��Ye{��ֻ&m���7qJ6)¸̖5���b`
�Lo��f�On��d��?�w��[G�l@3��ڔ��.�Fhb\�q�Gr� 9�����B�92�}���ݺڃ�Ʉ��s��n�UBɘ�˘*�l��.��LsCL�s���	��f ����i"Hk��aE�����훹��=���@��c�F��d	����g��� E!9��A�PN=�>���>���͙]v�-\T�@f.ĬL�ː����?J�d}�]�SX6�{[C�]�u�[Ƨ�h�����	s�J��dT���3�k�i&�F����n
�_m3�]�uܶ!��U?\Z�w̼��M���e�h_�%��x��A���c��j��:�b�s���B���g�K�^)`��~���29� '�0kQX�g�a'����Fw��	�5�S����ܵ�'U�L(�	7�����Ў�y��>��ae�1S�/X���>:Y��H��UM���M/�Y؝�֑�pڱ��0v��i+�?��O>C��i�>������󘒉}�5ea�ɞ��t]Fg#�J�/Ox��6Sq&pC[V�8(�u�����
T�4�
"���D�1� ID܉è��!a|9:��������X���,<`�+L�#���)�q۽m�x��?��B�'�TҠm�H����(-��;��d��Z�Pω��1ͳĜ�������ikU����q|�w��~a@�����x��J5f�$�Lo">����F�s�$�G�Bp`Ť�i>ۯ:���sw�e�*c�2�4�Z��2�����������h����l\W2~��0��Ǽ��B&�V������yI�$Uĝ|lx�5PB�⼆�81�Gg:�4v�Z3�.DG۳��"V\B_b)9s>~��D��ҽ���j@,l&�醰g��#tw��x��E
���\(Ϧԕ�pѢfU #S�g&Nk��_֖:�U���sTV�*T�d�d�Y�3���L(r��%��-d03��^OL(ʎ��*��Øμ؏�s�2}ȉ�c�ho��p��E�L�>�Zx��̾������)��$�4�X�9�,���88��S�,���ye��e�M�lm�!��>��*�v�"����B	[�O$�t}E(Q����-���H^NPZ�"~Js �4���HMV��:p�`��4[a�wy\�F�����Ԙ�Uejl��.�S��B��E����T[B�c� �#���,��6g���?~v��"��8����M���O��6FIU��M�h�UzNk @�ybB˞���'N���bc�l��_GP�A�?��ج�67�D����h	��p�+�1�i:��N=�����1_�c�!"O�F�8o��H��%x`O)��b����aY��]�C����.AOSS�R�h)�&���� TH�#�x.����<�JkA�N`S�-V�l0�B	�b�ҤyZj)Pjd�a�����
ep��/n�(�$�@Nx^j�n	�� Q��C�(|��O�\��1m���P��+���1���;j>zk��,��b��Q�/�,/�,����1Fcek	W�ٖ�=�Iw����2�?����
G]1~Ң
W\q߂)�ǭM���� ���۱+�3�d��L���;o��T�E�|���iG����z�CC[��/�X(�L�K�$�y�]5h%(M��d��ۺ�:I�7��8`�p���y�����׶u}�	,+�BGT@�*�?�D���0�Z�q��q�2���^Z�FϷꊴ1x����2J�Re�����"�,��^��ϵ�Y�1n6.�i����lsg���"ȆC(Maqb�߿�V��t]V9J�X�|��y�nLJ���١6~I���&(��[]��t���bd�Cٰ�{3��e�w1_�۲�Z��*�;k!��pN���n��o���s�*a?������>�m����g���}�΃��'�F�_�n3ԉ's�r����h�J�/�_u��YV^�(���RUʚbE��u:���](�⊭M[�� ��
���*��*\	1�(T�B:�2͡���_�F�!^q���SO=�pt�R��<�!n�%>���T�1��"��̏�,=���#�(w�d<�V�����QC�`e唒�O�1�7��Y����1K��@!��5���x����m=nBZ�N�@J]`�߄���ZZ���T��|oڏ"S�LV��J��1߃V؂~ox��b�𨨕'=�E��<i�"�,���e�W�Pt��%��!�F``T&Wc:�:1�C�,�f������K�4�(SJL@0[��F�[AUV��7�`��[u߱#&	|�wQ�)���4VϏŹ��оw�~��2]Uh"{<��L'O�o���Ą�^܏�M�`P��L|��;j��խ=���A�olA�}i��d�s�Z�Ǣ!��D�k�,�!/$��վM|�/΍p��s��9�����Cėts#\�d�rM��a�/zG���?½��������ߜZ�����&��|�$�ʯ���"O��� ������H��U��7��U����n��װ�fK��E�g~F��m�҉�.�B�����0n?���+wvN���S���fOV���~�%ɽ�Ó����8z͇}����_�=���?�'�ꄢ�4F���q��~ꓟ����?��"���E�0��c�p��y~>H��!s��w��+�{��8q�D�9��o?������vv_��}]��z>��+ ��!�u�4p�~���H{��=+++��~4"�@a�5nD�W���`�Ub�1�(d�m�l���|�	��7��P+���*D����`u0�]�����b�w�}K�0���zk|Wxo�*E�����0��ѕ�?[m��ԉ��\�,�#=�C�P��3I�� t#;@@ǲ-�{R�c�5�X���QGG.��g�����`��]�K#�� �� Rc_yJM߶-$��F9��eG�Oۍ�^.a0��nEk2����
>tۋ~��u���k��|��ϝ�x�����W�����-VP���y\������������͏3ol�J�������Uh�a �[�]rqυ�y��41��"Ӫ	W��s�l$9���a~�KW�PP�SR ;��R�}��d��/%�
�ڛ���_����m���<�ेN�(˳!+=DՖޠ�,{v�"q��y���o���Xt}����_���w��������c��!�!�"�9�����=�ko�~F��>�LM8�(�ڎ�C�B��d�u���/|N;��q��֬��Q�в�hU���ě���� Ed����l��e���=�Y�~~o���gc�e��1Hd,� �@��ʺ�J7�ԧÎU5��U�{w��s�9��Q�kW����� �x����,�Z�_�4.�}lзp��d�J(�Hī�:��'��c��'|��z��{��:�?1#xN�#ޡ:��!��c�'���;/�k���_����oKO�	�[��fy&��]󾘰͸����6��� S�͎a۾��s�?���-��b��\�_{�]݃?x���kPX��W�cʴ0�ڲZ�"F����6�~�l|�ҙ�#������x��#�35NX�d�V�Y���9���o]��U������8�y���&I�P��--O~e�ߦ�3�@+�O\��.ē��g�?��_��os�o{0���tZ�w�D�M��\T`u��{%��?����dF�N�*�F�t�H?�T�$G�h�?��AA '����;���W��Y\u�K7��o,����\ui!�Z�<�!��_���e\�V(��6��ԁ��&�ʜc�0��tI4�T�}����Z+/Uh�)��e���ª���t�d����١�|FK�V�2
��h�f�:_��{O=���>���n��}�7���3~笋�+��CZ�&@�섳�ʩ6����7�һn���<��O��33g]�F�uV�]���a����SLC� ���V��+
�����F�\3�J�ហ�
�Th�����;������6IM�ZX��Mfr��~��+@k�8���⨍C<�E�;�������_����{$�(����d�WJ^��j��~�F��q�ߨ��λ��粏��<���~�k;)��xa��]��d���')>�{\�!=��-�8~`l1�@��:�0H}�%U�<���{M+��/�`�ஂHJ��9���%�g��� �J�h��n��K��,�]`��1@K���ΩV6���|	��
Zȸ�d���0�x��/��u�����>/�S�����(]��WdY�S���X5�����A���,�?�V��夕\�^�X�����4|Vw2��3.�Cx�y�xR��DZzZ�&K\�-F���k'���g��quƴ�t�@�<9�FW֤�ʋ��2�Y[���|�o����;o���c��f.l����t��v�U*{�M��43Y�j���Y�o۴M�t���~刨����۞���O��4�f��+����\������Lz�>U�f�ϡ�`�X�V�0��6[�Va<# S$�e�
 ��h�{�c7�o�i6��su��+[Y�u��q�}�����&����8[?{��#/���a�^+H�r���o�������_p����ڶ��w�'��B���:����y(�rx���
S&�m��W��U��L�Bm'�3�G�������,\ᅋ/|<��?ͅs�NY���}��g�D�c7��!��f�t�Y�ۯ�x:{ŉ�s��ޯ�.���4ء�o�X��H��
J<�U����(�O@J�����t��@���c�$� ݠ�,����W����_W�����)O�SM�_@�:B���t��za��B	㗺�ZxZ���@鍩�)V^Aj�{�\���T�Y��Cz_��x���9�뢏��Ȏ_�����|���ꨫ���鲻�bާ.[�n�u�S��(�<�}?���+e�zǔIX�h.7e���8�)77�o��6h�����J6��r;53��E���u�ל9�=�đ��'��|�_X����<��d��#��T�2f�3c����*f@�:鷍�A��4Ө����]|'��}�����׮Y>�!��P�`Rha�� ��-HjFER��k4��:��#��[��;��lHҭ�&BN�C� 1%#�9�9j�?k���M��^����;����A����������xy5[��f��B�]�g��ͤqί-��ss0��hba�P���`�lD)�(J��KB�ɱ����P���J��-��L49␲��U�7S2�F������}�/����Uo��S���.��;�J��6w�i�1;
����ַ_�"ܻL�.�鞿�k�|n�0RJ��E̖2��@2R7B�3�ը�����-xu!������v;�5�Ǖ�V>k�9&,K%�V3������^�u�{��p!�V�=�\<�����a�?t�����x�zf����J��ĸ��T���o�3���Πv���S��^F��\_'"�d�d��C� �7�B�%i$��J�TIu}�쌼��SiO�~�^�z�
��>�+�,X-!h�G�=_�խS�۱{׹���<��Ͽ��_����?���^�^����l��[�N�m!�<Z�B���#M�8�����y�bGS�G��zsy��zۛ�]���}E*��S��yw9��P�r�D5V�'�(�d^!��U[y��=1ߒ���ݲ��0w\R�kj����W��F��Ϳ�λ�ySq�wV��tz�&Gb⍬r��D������]{�7��.?���,Q�0��@�Q�!7L�N2c��t���Wkԭ|o�sp���":��$t��P�ޝQ�|J������_��g?��k_��-�ɃIo��][n�Z�V]��4�{nx�/}�GG�s2g���$|N���e�;���+�"'��#�2�A���� �a�c-_xEL7��s�vEE��G�J܎���`;��A@� F���Ăi�֜�Ftu�Ͽ��3�xֹ_{|���D��0-�4�3A�d\�Ŝ��9~���^���2��wi�P�S�S�N��k�a,-�8���ïsLҲ|����*��j_����*M������|��D��M
9�����G_�U�I������E����˯��+������ʉ����
��BA����clNSͧ3c�ǂ'��e����m�U!�Q���V���[.��_̘�\�d��f�1�eh�`��t�hb�-y:��	�~�t��e��q�ݓ�����[n[�&�`���V�����g"ߙ�~�y�{�m���Z#�BB�-P͝�	��Lkn��Ӌ
Ǜu�+2��KzJ�6)QZ�W���=w�zF����1�R��M?i�i��m"54!K6�R��!�������ۚi��N�ަn���i�@�:�7�֑o�zw���h�s/~���������T.�*�Rg�z((��Sy��(�^'mG�~\n����q����n<���C�ry�Y��ބ
YKw��s��5���}�^����H�hxF�2(�G��Ł��k��_��^��#�S��H���N�kS;�{���Y��l��-z|���X�'�"���=3.��>�oWj~FRV_х�%d��ҍ�p�U��V�&��󳽥�}�x��U��:�w�~��d�m*�#��YU'kc-��)��+�}��\2�ɥ��E��v�D!#8�D�� ���u�[X��k8O�<��׍~Ȭ@�P��-ˑ���o�1�����ۏ�*6�y�+ߪQE�,)���Kc��!�Fm� �t�a-6`4���ff'�$tM!()rr�#I��`b�@b�H�j�~iL4d�uV�}�o�ÊY��jq�"��|0�~	o#��4��Xr	��=���i�jDz5��C���$�j���|�a���m~]��M󌸾O��q�%i]JXp*
�~��<�iZ�l��$S2/6'�N�a_��v�ah�ܗP�G5��]R0���a���mKi''��i��?2>�Iб�N�z&SS3'^M���܀�����jW��t���lO��7��L�'?�GBj�F��A�w��	=�I�<���.��Ǥ�Bט'Ċ]:X��4 <r���4�2�r����ortpZA�J���Tp�u�\�@	�<ǚ�N��D������W�&I�V�Z�S�
7�U��DH���t������1N*���u:�LN�z���Ʉ
ŧ�*}Q�Qw�nL,�$ÁyG�����T����4
�x�J���J�5�77O�w�'�P�2�7{_xL,����ꌆ��=ɉ�ۓ-��v;�,����8[A��)d@C�WH�IW�	A��=x���<�Z[c��1�)j���	��hV�J���ɮ�A�.Es��¦�k�:���b3-��13�����$ٸ���!�H��P�l�>TK��{a�O��e_��C����}G�{� Q dNKQ&9���n�[�M�޸v�nֆLs���t:�sn�\�=�yGQ�I`���&�L�k�pfh��@�V��4��DZ^������c�6�,J��y1�&	�b�!����k�l��0P�hg�E���5���n�G�A�
�3���Н4�|��.L~Ɇ��m�*`�������D�=�:q�͗͵��������Ú�X�6G�<�s䴴Pϖ�Rjr���^�A};�����
c�R��!l�܈�h�|"���k��B����a����Ʈ�V��sl��0?]Ԓ(�d4WI2�%!�~նtjlG�_9Z�/<lK����=�l�IP�p������<υ���%������J��!JO�L�fI���'�I�ث]s��dAH�Ͷ0.{�Z�	y����JI���o�Z-qd\�1E�9/?��>�m��M\_ &��\К��:&#70V��5�_ɸY$<��d������Je���az�b��B���l��lqyC��d��)�i�\���� ���2�����sV��2ch���3fu�aB~�#�/�m��>��iW1Ts�u�Q( <��*jM!��0�Q�!�������=�z]��w�3��3s��g�F?�?Ǹkk�@/>Z"I �Zb�>���^Y�*ll�}.@+��J�b��A�BOp@�y��AE��̵�M��4��V�7�~������߇��ah��䝾zu�#���_�3���m�Vi><��x��-�I� ͙Yp�c�pSmѱ}b�$�-{���K"��[�܂�j�sˀ�&,2��V���4���WW�{1 ��ѐF;j"be
���[cE�(�� H(���\:t��]q!�L=��i^����қ�ah��i�q����6�F-�N��`궵�;��6J���0et�B��~ �w!�Us-|�3����)�^-YB�L����=NؖN`9����F -����o���6D�TO�,Z`�ۜ'6>��������0�^�	;];*�G+89�1Ӷ꿪�}�[�z���
�ķJ�L%Uo�w���V-q�D���辐nEe��@�@L2��f�������ELƇ|�T�A�`j�m������`��~���9��&�|Џ��7��Q0��Dk�>��]���V���$$�b6�W
��1EK��T��:v�����O��lc�3i"�8f�K�$+ӷz��ks�H2�u�M�`)���bږQ4b
F�j%���7:ST�k���E+,����d��Hjq=3�q����V~����l�:�����Mj-?o8��{�ͪ�KU�W���Qj�N��W|��BT����h˯<2fg�T`|4�s~&֖�����H�Mm���#��J�
�k�2�i�AX���7ob�n�y�?�e�⑩�I���q��*
����&x@�駰x�e�����Y"+�������4�4�0���5������@�����Ew땻Lڌ�ݓ�E�06�axцPO�W�*�	O��n6��2A9�K]�_�pm�#��JWu�;��J��}l*�|�mS�X&��͒��`� B��|)����
��T2Wʡ~ܚg�f���c�"�Ü��D��V|�Jgi�Q��ڪ1�<�J����
H���C����dP�gRI��� /���	Y�h�C�8��&ÔqYH6�?�`���X�U_? M�<���]�"5
��wUa��P�aO��i��v���JHy<���8��h�EK�,
��w�Q���Os~l�U#��D�
R'~�2O8J�;$�ljshU��h��
Ċx�r�ohp���U4Hip-�ӗ��Z��@C�����gZ�����N�a��J��li���T��ENR�3c$�Pߚ��� �ѭKIahWt���F���C�glv������	F6�n�gq�	wF����I"Q`�9�}B���Og��l"h&�(MS�3�����a��'�q.mT�G۸����I��%;��qM���XJ����F�^E�&ꃘJMX�D�X�i�-��G%~.㠙#�U�۞˼�lp�i�����T��c����%�T����E�٥�����6�8��1�L+�e� c�s:�GjQ�<��޽��!�o��*/�Mg��e.E��a.y�)�J�@c�ep�*,5E�\�R;�cscE@2,*�b���Z�.k!�1��I�y���ɸ��K�"-�{*0+�@��ZUq�{�_3��0� � e�B�<ɹ-�FL��Y��8���r�J�m!�+avB!~��vcU�}���D$0a�����B�v�06<��`���wu�oX 6�W�ީ���6%C�	0�Ih�0h�w4K0D֚��rT�%%BGV��L9S>A��L btG@���Ê���6v��,4�˩�/��/5���6u�n��)�߄�1����GL:LԐ�G�fT�/H�ޥ���Ô��-���[���>b&������|�J���x��!Z�I����X����I_���ce���7���I `��5H�m���ݜ����?4��|7��Ꮳv�����=;ȫe�'t��}ҁT'4#
�����L�͍����s\1��(�8�����B�ܞ�c�HdH�*�]��l�j>{��
��-��b������7Y�kb��v1�P��/G�L���� .o&L��[�fS�a���ΩCj&����)���� s��d*a����<t��8ƼR39iYP ����Qj��2#0��Ȥs8�Ml|%�pc����4�h�B߲�ׄ��JX�:-'&�o����(�CG�B��I�f:��<���`�~�|�Ͻ�%��ߐ�^WV����4Յ]��ʁt�r��s��2}�Ѯ����i�#H��2�\+X8��D�j	�:mӨZx.p�&T��3�u�gb>��31���J"�oC�	ͱZ)C����A %C(�z��c�W�����fj]�Sd�;�\�A&�9��_�oL6�`k撥�0��ch�k���jĵOb�_u�3�XD�&ըX�C�j8�6�!6G�Z��$8��pR31B�o���v���8�@w�s��Q�
wy��AB��d��\��&��u� Q����)9�ox��F]#�3�̪�������z݂4#ЏI[I��-����yFv� : 3;�B#|(��>�Q���6�&l "���O�`uwi�Y�1���?��mꍮZ��HХ��" u2��Z��b��yK(3���J[�2�ai�>yJZ~@�$1��"Rd�rB`*)�Z����qf4ea�&�8j���fgT�W�J_�x�dv��]�z��۸�|����IB<�Q�T��s�o��k��R(c5���;E��1VT,Y�ƙp�$���XA�`(�p��3���2!�  	d���2����8B�I����H�^'q��i���`;�<7{l߀!u������7ʂ�ƥ#|g�e \��Q5���^���	|�1�"V�MT���t���c�z)h�p�s�����@��,���~G}��HO$�$���#�p��_`[����s��2?T��:5H[��ט`%I�� �gLN���# !�P�IA��u_'���JM�љة�Yja4\ג<}?���C���!&�L]����`�Ì# Z�U�m,24Wj��b?�A�(�fFQU�kb%���iuap[0� d	b�w.@�B�UɅ��c\&���
������H͇�5���T	���Toֈ��X�a�J��$L8�o��X��3��tvρ�^���
~�3d�q�S�� ��,�!����i�B~�@�0�j���X!�7}��\֔$�=*!��#s/ _%㕺f�E�6S��ͅ�0Y+��#[���FQ�f���c��P���Bs��q�ǔ�2S�ņ���AL����� 4��ccp�Y1q�ҡ
���ȵ8%s�	@��k����"C���`�(��n$gL	}u�X�q�blŁ�N����>1���������f^!����,�8j-z�1NBHȗ4T+(��0^�T�M���Mz����M����Ġ~w�t�ij�E�ᐛ%z�I�V�j�]�z�K�7�u��z:�X]w�w� ,t�JG�5k9��Vƒ���"�z����?	� �Y�Np��qӶ��d�4���^H,H0�b��1f�LP=�����c��VP3�� �f
A��A�,�ryN����WY��ۙ��t}�&�R�Rg6��S�M�<� z�0|n���dZ�~�o���&4�D���n��6+]�J',$Z9��p����:>_M�y*��=2~��JWP���fJ�`� ��  ��χ�"4/DM2g���ve����L�
�i�^l)��{��������'��������~�/�4M��>R܁n�o�U�����t8�g�>��k ��G��B�m@E�4�ȕ1\H깅��<�
�E!F֓P$�ϡt�Ա�%I
O��L�W�k���ϥ�W�J*7[]�<�g�����RVv�,��Y��&�Ha�c�H���Şۥ��)�M;]��ę��b͗)-������ܳ�Ѥ9[���.
UCV�O�X��z�f�" Z#f�3Ӹ����<s���F��.r�ll��,�b�&7f[2t;�p =�'�*7Z%D_&F�b.���k3�*��V$tĚK��q�^������߽�jw�k߿�vV�{3A���yB2��j�F���FG0���6ա��:�4Zu(�Pyk�_�?���`.q�V��3��	�����|'���f�Gk���J];5&��<����J;�f�4�/WJ񻕎�<(Cf5aa����	�IN�*��6��vJa����b��Olxd(:�.�SS�b��eh#$AYYh�P��¤Ih;<5g�+���l!P�Z��Pf|�&{��V��S?�T��z��ц�P���f�(��}��ש��Miu(ؼ�͵�q>����{3;>P�LW�d���Q��ӌQ�?����p��	�F�M�ޛ�y�{��q���,�$^R��>T����Խ�������V4j�d1��d�+�ܽ�.ѽr�?�n�c��7LT����יw�ju�����7���!x=kNiū���WM����REҿ��<Yk�I������{��������_V��9I����W�>Q����:�KR3�N�9�*}P�WO��f�YA�_�)3Ӹ 6��2S�djB%�s���-��Z����K�.y���ɜ��*}���K������Ќ��__���Ӄڷx1��,��5�>�:*���C':d�l��z1�����C￉1�Ep��7M���'݊�rR+m��
�E���_���B]��}��"������m���0��^h�;I���lu���U�>B�.� �﹔n�Y*��d�&��p}��5[04n��f�
�Z��@��"?����@��D��,�R4�s2��Тᒬ�����O��[���ފ9�r�~F^�R3ξ��%�@��{�#σ���2�{�"�į�G�|��'�7_!����@	Y�fH��V���QW�K���O��LΗ� �L�z�ث�_�H�*bUӬ���2"66QF{�ebh�Gr%�"�h!�k�H�?���/;��{.'�o���Eu�Kp.+�\�F�+�����@!D�/��mN��MS@F��v*����(��Y�:����o�I�B虰�d?�����#奞�y���b.�R�
�q���歧�s��|.
f�����̈́(CDu�!����
�I}�s�I�L�82��d/}ޏ�����hn��4J6��LC��`��TҚ5�-��b3l��`�t��Ѭ�]W����Ģ�	��j�����5���W0mHX0��i�����/�9'����}����{����E���b0��_��>aC%d#ߛ(@*Y��̡87/\Ρ4��ީ�c+N�CW��h_�UQ)@��/�_���(j��+d�~���t�k��]����ܗ^Թ���jI%}u����u�?���{[Q��4��W��,��I���J�OO��:z/���jI����E�Z<�m
?�	�e�M�~�d�I&��ݘ	a�ޖ�\��}�i��n�/�y��?8뼝��y�t�}߱�N����|oMm�Gj�n+ �$�{dE���:ͬBf�bpL1"ܑ�oK�h��M�R�NdۓƦo�ym���|�����[M�wz&��_����Di8~r�ݒ��'��l�%B���p7� � �:3pf�3�v:+��\��z��˂�B�C�$Xou����i�RҪD䚪 Lo��gh�s�fS���8���8���Os��W��J��˧}�gg����o��O~����w�sh����~�o�������U���Ok͵淫nO���}�`��+x��B%�Aѐ�����~�M�VN�!|�i���m:��1�c U�w�ծp��Z+��}���;+t�+�{�酤;K�>��+w��^��Q_|�\��j/�A��˵(��?~�����c���Ƕ_y�#��WB���-/y�w;O=�� ��W��Q��D&������B�ш��vF�$���7�(�iyv��|���K�B�����`|��Fn��@bȠlz�2럿��sz��ֱ���;���]|7l���FQH�j �i�`6"$�!�m3O�όZWp>�~R�P5��
��6ZTҔ(���D� ��z�|��i�V�#s�^=)Z�d	�\p7���Xm� �?�
U9-�,������(q��\�/�y��o?�U��M�?�ڈ�ڍ�"������O~�����EN�d����?4ό��Z���U@*2%�g�^�(V>���_�����᥄��O��򭏾� �^�O���Z�Fth9��|O��<�̫�q9�Il�}"��:,u�6:o�N֑߰�L4t*���P����$���I���� (���c&"��S,e��%���;��U���:��t&�$?�S��[t��-?i�n���<���O|���z��=��_�ƭ�|-=z�������V$�B+
Ƹ�L��Sj�j"F�gş�>��8�2��s��8xV��3��jb�6�=�i�+
iЧkb~�EZj!�M�m�T�Ea��D�R#L
ᐆ�Pw����ߜOS������s���=��΋�4|�t��,�P/Z^k�䝌��J ����}�R��m�X��(&�dڼ1�UX�s��P��P?�{���Q��P�[E�H�����!�C�\&?�x�B�x!�0�TȸoCx/r�9�Ie�d�o��&�Q��m՝��"GX�-�Bj~נ�a���B�U�o�|�ż
�W�)'����) y�uˣ��N�@[�z&̔��`���HwLêN���6���6��/�P��A��?��s�{��4�_=�'������o�w'a�K�d�e&{���>�A��E4����Yշ1N��{6E)M��s�p���>�f.85zIJ�4�
0�+-�������N�yh�Ml�X���Z5Xc\�J�<�ګ'�]"z
�>������>ĕC��k\q��]R��5u��?����|���j����G������p���=E�3`/����9ҏs�Л�z���~Z�z�`���Xjl\HM��m�S��D3P��_�gE�H��Z�9�B]g�ƐQ(d��bn&�k.�}�?K���#��v{���¿4M���������Je6�&���dJ��ez8Ja��/m��tBű:����T�i�t�����u3.4�F}G��8O�6�u\/�x�V8Di�Xt�v�LF6�?Z���c��1�GF��#����yի��u��隇3L�»Ɏ�e��
�6��D����%s}��B-�!�
-�����>;��g^Y������z(J�s��Z�f�o�+����fz��{��?~F�'��#d�T�v�Vy�Ӎ"��!��C�)�V�k��i�:����Q�ܛW�B�Tf�x�~= ��6�G���u�m��V��>���N+z���V����oZ������Z*0�@I�:$�Y	|�B.�s���,'z�H;s6xA�15�l�Ш%��q>f�X�2�4�>�4����� ����"]�f�'Ev�;v���"�����Kɋ�ې$.;���D�t�)���$��H�˗�Lu�j�肛�l�%����Ӵ�Cϩ�#O�~gMW6�Yh�+�Ry�8r%�S�DE:�Ŝ�FÙ�$NX,C"�X��> ���3a�xx�\�'u��<�	V5�Y-�U�w�<�z���Ưo��op0�$��ݰҨ�U!^���f�J`2YFt�j|��	SB.��O1���ٯ>�" ���������8�'����;���"�ǒo��q����$v�:f�W#�N5�M�g��1��P�N�m�k\c� ԴN5t"���*\-��8�2	J-Њ�V{df�X=��z�Km����t��Ύ���v�i"%�|aǢ�z���u���3�f�39���mZ��: "a�ч�Vo�1K��Z�D�ȵY���v]����:�����5�$⥏\v鎯/.����vu��np�w�z�],�xV��/��Kj����2׀���u'
�I-��>�jǂP����r*<�ᥡ�Á�l@�d61Ia �n(\��$��<�qO�uu��Y �/G��a�,�9�L��fG��@Pr2�j���)�vx���L=[�|�;O2��
�J�lDj ����31N���_��V����Y�,&�~�(������O4:wmPs^vdI����\����V��Z�!�6*3��ve�ȯz��q�PohC�j♶ �"���o���	�o:�l�7�?t�.甉k܀Њ`NC�Ӗ�ݟ�&!o�#J)c�Ǐ�֡m�^�H��|��t9T���3e݌��h���gTf�3a�9�(��m'�TǞ���2n����A�T��T��Ȩ�@J����$py��t�+��v���e��[���9���o�;����{�D����Щ>�R�ʎ�A�<�\��+�jZ�(��6v;ZF4�(`�L��t��g6�R���Vk���u�2w�uB�z�j&�F1�[!q��)�2"(�� Q�.�ye�Q�����	(4�A�z��
}j���l�	���%r��������6J��W�M+Ջ���1�"�ݙV���v�(��-��� u^�dJ�	e��W�Wǅ�'��@��A�H�hWg2 �4ަlս� �;w��E�D$��	��ǂX�h�����{��'�m�<�^���X����Y�>	�#�I	z�f�bX[��}��/6�rw��m'\tH^p�cFb����7j���c�t
r&<�iL4��ǯHk��� ��s�{o�k�����Sͬ�'}�>R�^F�=��i�p}-{��hk��$�n��Bf�Q?�W�j�Gj�>�*�6̏B5g��l��IN�j����	�J��l��l���%,R���,w�BR)ڐ���#��6,�_^S
P�Q�SK`����n%�c�Y:��g�g����X���7x���W��<��B�܏�}?@�o~@
^bEVSu`D�٬Q�o�^"x\�8�;�!�4�=�����7�(��������S�uU��MJ-�k�4�V���`���d~{o�M��Jʭ��{��!˨Z{1�~O���Tll��E�d�AɅ�������R|NiQ.ouG,�I�q�
��[
�w"%��B�k}��y���6o������y�D{K��,�C����L ��3�@,��C�铤*��d�3c�?���ȳ���UuEبZY���S�wFT&��Z@��#�����lBYh�I���3��?��Żx��YviAZ?���s~���	R�ytqv�<N��S�$D�3
��L	}�a���4U�G�8���(므�q�CY]g����� �pu4Agr�dug���0*V���#3�ܚ��1W)�J)����:�Μ��[�
.\�&�Az?6���bV�\�@�H�w������Q������0ti�ed�6� �T�mʯ)�(��vb4��id͐�Bɬ@�q/o�t�/�O4�����Y/:��'EBf��Vr �
@�ѵ��C"Lp�tFB�-5��8L}���I5t2kzJR��8�t��B=��h�Ol�i��kܔ�R��_�'������U�l�h�r�y�GjR�-���-(2'�Nb�%��y��fF����o|cc[&~���.L��,(���3GxB�3�	=cB��3v-t�e����Řh`��BLv�I&�`6vc|��(<���e}07dJ�K�]���5&n|�^r������g�[���1�� "�z�����G�:�����}S�(d��@0;����-�­��4��3�Y.&'%�<E1�Ѹژ	A���e�4��uE���7܀q��9�}ֽ�<t�&�캵����pW2Vw�w��ݛd�E2u�U}{�J.�R!V�������R��u!JN����t��Qc��|膤���	�{���P}ҩ��p@�>n��}��Ō��|H��o���y�.ڗ:l�Q�Di6y���2;��7w�s͉��ޤ���s�#q���mn�H$Ḭ�����PpO��©�,���`	��1�N��:�v�m��N���Hف��@X�Kɩv���*�P���t8�������%d����Ŧ
�{;w����d<�%Ki�G!�/����ɻxmG����/���������J�P◂3���k�$�5�U%��.'Slk/���/\�W���V7�����<�/�yC&9��Q ���Ή(�S������@6���d�fxi�L��F(��c[���s/[��]#��?L~5��O��X-�d9��,�����\f�Ӕ�,9J�S]A#A`����1�ֲP2�������L�?��`u�Vz�DlV�f�{ �N5�^/'!��G(�2�P���q+�)i���%$.byų�vn��{����.�(坫�@s�A�%5pWrL��Q8������=�<~"�Y^o�\����m���e��_�)��%d�ڻ52ɪ�5_5-@?A���*m]�?��'�m_ՉNdΫQ���
j{ԕ܅$L"I�V3aX��&
CC�zF)��JI,�VjBpkf�A$6$��=W^$�h ��x^u��;��D���ܳ�����xd���@~����H�G�KV��z�5W����/D�%Z5=S�F]O�M�p9�*�	p�T�m4���BD��Č��M��p�$�)�5�9��[>�2�wB��4<���-�yYA`��������7t����<un�ǹL��V�&�!��Z�f'����{]��f~���}U=��K/�'�N����f�t:��P�����Ix	԰7�>B��������f�o��@���[Wy��%���i�)��ls��;�-����CZǿ�`3�VvT���)�Vs?�AT��?�;�Z�q���5I��D{�4;�w"�����R �J��b,��bd���v�)�U�*^�' �j(������+0]ܵ��6xt��7����M�AX�%E��rf�ه=�ƣ�㫯���;������^�\�y��]�)����U����m�zt�t���f������/_=�9��[�y�e��L�6'�x� ��F���Q��.W*��ˌc��0�����2%�Y����������V��҅�`X��ez�8�D���7�+D����s��������dn�����\��cu���4#��d�so�,]$ꨰ��߹㐼�c�[�F[���9���v�4�z���B�M��k�p���R��&����
��h�w�(�S��F ��ĸ�	�;j�d�Z�1�	^�v���0��6�ǯ:����py�����ճkA:����;	�W'dM	��^G�`O��3;lhq���U���%��= Ni(;Aj�ҍk^��;T`)�/�Ј��A�Ma����B���[��|�4yח��E�U���[!��m⁂E�B�
H���9��� �؁���hn���i����Baubl���&:s�\��O,���,t��!�eȪt�	��dVȖ��c�+�T��,�Z"#��  =����Sw=��hA�o��|@]G��������<՟9��ݝ��B��J�{
<���!:��1�儔�An�����I*������o!e�&�i���R:�J:�JKT|��^�gPq�1ԇ�6�+=`5�:�^�G�>v�����od���:W牼z�o�����!3$K���n>*������������Cl���c���x^@2��(@�$R�lø�������y�8ݐX7�!���QYMt��ax��O[�p�������qVLp���'@�߻�0��{W����zw84��c��֣Zmy���T�ZQ�=��EFt��3� ��iS!�����ʰ������ ����s�(�	���R�!;y���#�q��ߺY�:�|�S���L�uQ`���9�֊"!ଧt@��'U�@_��U�c>MwU'�8���M�JW��E��"Y�	q�8�񽦸M���5<���t&`�B��gғ�(��)�%���T��3"���r5jԮ��?���]�%�|۷JyD|$��X��R=�B��(��1]y���GU��#71DyQ��BMZ�s�wȓ�n˜MH��<(5�I���Bf��Ǫ�CN�Uն{�T_B<�-�wd�a��������Ǟ>��}��b7f?]�?t��w]���q'�i��w���������o�8ҽy�c���� �$6��ܐyI9��ce�����5��|��4]�z��6�QS���l���h�����!��=�w_��߽�O:WJ��fJ���a��q�Xr|~8̂'h˻��7�p˭7}����j����r_*N��¦K���TxީDߟ�&)[����rZ��m�C+�RLX�U6��|�Jjꀑ��je�2]s����6�Dh�Տ��ƭ��G�ѳ/  ��IDAT�����_'�ґ��I�^�_�3_���� kH(��B(����)'��:>㎏�\�-8m�g��7�J����B���2�T�%���6�U��Ǳ�%��*Fs����13$dz������_Pi�F2��H�1Էe&�>�j����~�����+�;�p�w��z��M����G�o8t�y!��qI���_P�(�m�,c�Ũ~���	c�aL�I��/����N�)�O��P=	�t������甋<���u[A>u��a��]����)ġ���<6ǂ�/��������k���]��8�&��O����ǹ��c7J���&���l)���M���S�T��&����������5f�~`�a��h܃�b8���
ɛ�7eA�f���{����W����4t#��)�|*��nz~�1����ܭ�Ó�?���^��{�<y����<O�f��t}��B�)�P�U�}���&Z=�ٟ�x�M��h��`��r[XF�8��ʀ&m���aU�Nx�@ �t�Ɯ�Ƚ�P|�M����w�������ns�7<��~�9�;ܥe!k���=��T!�<�E�Ay��υ�pz9w��Wc�Z�٪o+�#�ncw��'+�v����S��J,M�Ft!�T�
�>�$�<&h����:�O;+d&���'��\H���_z�r����W�{կ��]�O�������
R���|�\.٠iX��m�������P�
4Ӽ�l"? i���4��fP�Ǔc���}L4!6�1���\�w`/F#�d.݋��_�s�~��Ot���B�����$V1�p�G�8
b��<�v݉�=
��봳�p��_-�Wí�Lu0��r�NvH����M�Si�A�B��ss	����4`m�&dr�t���0�}we���L��&sf|��y��Z~�,4w�hG�y��>������>禛��_�����Gn	�Y*�(� I/�lt�&���g����<��)O(%�t�E��@���	�8H�NV��,�`��A���P l�!D�PG̲⎦�?�+��q��(�=k��x&/��n�s�ݦ��ۑ��|I���C#�^ϡ򈽆Z���y_m��Sue'c�)y�R�ϑ�p���(��ӫ�>�w��KaȪ��[�hj\/D�L^VK��c�azR��v��
�8('5���Ai/��!�a�P@[�	\��l�]
�L`��B�'�N�'-��Eu�po��'����y�c0Z׸�=�ݸE �Mh>`�����fD��{�u�$q�(R�a���v6d(mL6r��S���$���oP_�\�ᕣ��u˫>�ܽ<w�鑧;���ˢ�G�uRS�S�JY`�����K�����sjbu���'S�V�|/�9����6U)�^}���	�VG��@��P�P���i�� �K!t�R]���38ĦqA�#W]f�'�6M@^�� ��e�X'"�̋��+,��s����m;������Ï�����"%�B�E���\s+�]���Nd�(8v����d}&邧n["x���[_(=��[�]�m��&:�:Y�6�ᎉN&(Ԅ�2d��=�`& �/?={OO�JHG����s0D@��d:Q��1G-�뇬�=�fy���#���T8��*�)V�/��5�6���c����GY[���������9��BZ���8+�J�JՕ�`���3��̈́��TI���GV�i����Z����uM{N��zi�Ē��P����v�Mjr-CJ�iE�L��8%�zD�4!�R+�������SE�ŸUH�g A��ܛ�X'��+��"x��3jHմ�l��fW
���/�$�b;#���dY��h3<���uu=�k�s�Vr�߬-�D�S����}��ɾ�T�胕�2�Uɑ�.<3L#\m㾃��h���8����pS�6�U`����}�$�Ŷ�/�I� ,"(K�b�X��ޒ��5���O�>�g�]���w��>����,.������v=�t��6a��1Nx=ht�>�J�t���T\Q�Z'�H���$�_���Zv��mu�a^ИBB�I���j��b���N6�자K1tM@�%X�^�����'=`�N����)�����㵫$��5�26�,��~��G����9��,���4�~�q�jh3	�d���a����"��~-�tW�{�y� �e�Ҋ\�p]��}?X%��\���I�h�-nF�'�����<K�9��U� �'#ciX�LX����Y������V�Ў�^p!�����4 �3�9��4P�j`�1��2 ��3Ƌ��j� �~8�K$-R���K]�_�/���P�4�|*�X��r<,n\}��T��4�LuW�SQۦ��Kyh%*��+�P��jT�����T�_���9a�w 6=���P8��\����8�#���tD�E&����x	����VÌ�[�I�ff�ȕ%m*�)!�4�ZM`��I�TO��9�#�I~A�@6�_��?�z���+~p���L'։j�<�\'�ߖS����i�O�7u����Ju��r��["x=^���n�C�C�&|\ �bf�������W7bC�f���Y���'���ߔ��.��f^$�Ә>xࠫ�'�P��-y��;�<����ʉC'>��:\n�_��	Yy�����6�ḥ�՞}�J<<�Ǫ��{.4j��3�ԑ[�z0˸F����:�N�4ۘE�N/x^ �^���f�D��D@�*���p�`�Rv�C#���zWm?�
Q��3��Ot��B��(ՌZptR�^���x2�@x�M22�ϔ�L��?��wI���h��@6V�vi!jGMD�9B��'=���P=�s}��rLxN\o�>d=}*Џ��/_����B�֫��Sq�Ug�#�}�Qz,nιю��)�� ��}uÖ5N�O�e�]�*mk�aMF��L4 ���*u>�����W���4'�u�eB�����q��'��}��z�����N��\�����Ş�D'�mf�;�&+��L�`lrM-g�?e�&���	q�m�n���PYr+ �,m�6C�uptYB&��Rq����A�8�pg�o�s	N�$s}���RD���8�G�+�>�"-h�E���޿P��>,r��N��+ȯ�:�E���zow��9�z2#��T���A3���0��=�yYO�L�: Owf��X�
��&��b��fC�˅��X�W "�JlGj�Pi�T}R;�%����!��k5�z�`j���זZP+��B�w���I������B��i3�3M��vR���(�R����|���}���81�}\/�mZ&��F,U��6k]�`hs�� 	� �9�"?�����i�>Ÿ{�[H��vȒ��0��� �2'�F�h4�u����کT����I��B�SR�Lj�5JMcV��PRE��5���6x���)@b-ai̍Зp�e�6��5I��\�|Y�O��P�n=&��J��4#��j��m������"�����?W�fmu��|&�1r���M|��7�-i��"����┉:f�h�[�5{8��5l@���^���ɳd�9�k���� 0�x�2uA�%�W2@mG�̓���&HP˻+ݕϨ�}��N�9{/lwɕ��D���U�ʂ6)��(gw����i��L�h�t�
�;�����I�6.��ցd.���k~��X$[�)�bd��$sL�P<�3*S�}��B�z?K��#�?�x�c�����C&�3Ё�soՒ,#s3>I�9�E��TG����(�Hf�h�봂W��H՘�p��A�"I<�e�T���0�����JI��Jbg�=�X{7 ���"y8I������ ڽ�Ɉ��9a&o�1Tu6��*Ѷ�r�m��~���_u=�n��W�Џ��c�񀸫Z�F�p����Mp=�hnfh����o���@���v��M�L�ӨZ�n>�}QPO*<.����P�F�f�$˫j��N�F�U�j�G���]�v6$���_���<�ƻ-l��γ�^�w&W�9�����:,u��!
iȄ&v�t��u]v�%�l�#���Pu�"Mlr�~�I���*��ɺႇ�'�N����#����1�QjZ\�H�Th1- �$��D����5J�)T��8��N5!;�u<w� �� ���s�$�lC�F,�(���|eד^�ARپ�|4�Ԅ�9f�Y�HH�c�����Q�Q���S�@?N]F9c:�R�AVᆐ68F(�S9� ��߷k���_������8����{{Y�z��o���s�4���1��ǵV�'�j����0�H������&'K�E�m
AS5�Qסl��w�d�L��a�󌐇�@oh+��b�����?�o��k���z�]s�w:��ӭƜӆ�3������
!�������yŵ;�a���k��{r&�&P{�!u�FJs&�HV}A`�=ߧ���`�tO/�x!ƒ�W����P�\��;���+�/.:K��$�d~0��M��T.�����$;v��J{;���`��^��Y���@q _zN�_9z���^�Q��|������O��muVc���Vg7Y����并D�2�F��y� �1�� �#`�:L/�N��@]<�ِzo����Ҭ`�fL����"��NR�c�j��T��Jj�����ШP@��j���ay�Y��D�1�$50 �Y��ns��qB~�^���S�9TN2��o]�G�]�DS��v�Z�E����ѡm�Λ�5��d���e�89[�k^ߨ�/<H�Q2	��lĲh.:�պ��>p�%Ͽ���,䍙�q�ɕE�8)�,�9:���-S�+�{�5�~s�v�t�}��?}#�K>+6It���y�R@J��h~>ɩ�9t�)C���)L�-)}��ݦ�^��[�������\2����=�g��Ƴ_�_��5��ƫX��%3
�ք��X|׼����ϛAS�/^�څE"�Zc1�a�>��}���Š	�k�"�=�Z��)���ScL�pU��N+H�H	����5��w�3���m�����b�N��9;h���"��};�أ�7�p��_��ݽ��_���
�[?�>����	���&�KwJy�Bh�|���!���?�B0�gS!J�m�zS� ��������:-�T08�8'k鈕��J&u��6L]��8��H����2K��4��Z�I�r��*%�[��5�K�Wr�� +9D���R���Opf��Q���K��e�f.+��M]�%ӕ5����>#��q,��#FfH��֡����8�.>�Dq�:�s��?W:r��G5���ـ�ΐ�c,9~��ݱc�9O��j���Ͳ~����{��Y��)U��%�:����|��<uy�N�^��V#P�T�3_��4�RZ5ь6k
���D��
��}�ٹ�&Bc(GS��>
����{Ld�_�/�ta��/~���7��{?#���C�h�Do=�KwĲ���CG(�J��b����+v��J������r�����Mݛ Y�\eb���m������w�[��F�@B�4�d������Ǝ��q��1�!��N��c���`���ǈU ,�AH$��Ւz_����z���e��yo�[��{�Wu7J��[�y��<y�� **	5��B��~�;^�=7���^�J�4��@�V����F��Gd��4f#�M�]�o�����d��\��/�/mR���e��g�Tv�x�{c_�'�h�S�w�����]��/�3��_v���Ǜ�wn�9X`���7q������=)^k<�����Z��d�
�b�Z���p��U��ZLՠC4���wݜSp3NV9�?ĄAdWn��C��h���*���	�2����C"`ϟ��e���4Jn����>��R �9��`)�YE̹:�1�2x_O(��� ���L.p�|Y8d�%y�=Dww�c,�M��l(-��[�3�@�ҕ���%n|�w�����'�������7G}!��'��J�o|��x����O<̶�Z��f볟������;of���B[�8�ߠ��Z�JR��i��٫@[0�K�^?a�iaIƝSV���Y�V	�`��L�����
��HH�Ɓ&c�p"���7�]������W� Li	V�V���K��Ψz�����G>b����^�;�ޗ?���t䛧ev�Ѳ��r$*���~���N������C{~��go��ŷ�&�%��y�N̼[c�uc��ͅ8B�$P��tEq�VH�A�����<c� Cއ��E��I�9�tշx�?�gك���/��>��'>�Ϟ��wΟ3vb����u�}�n����`�������Ŀ}���7 *G�rS��.���ئ8����z����@z��#�����}6��>��
4���3@�7��Ʋ�40)xl㚯�LÇA*��<���]��ra24���H��4!��Tqr�6���
�T���?D�-���l����L����گ�W��mMd���L�1�	y��;�i�o��h��ϛ:IQA���5�+s�c���h]$x�a��:sM_M�PI��� 
˽�7��;�x���p��,JW&z��.{�'?�>3:ͮ������h����F����l�=��S�o�>�9�S,閆:j��. ���M�Sm+��a�C^ߏ,�����������������4N8�8��A�������K����K��5Ta`�@� �$Su,kh����j�e;&��S�_�N�?v�)ֹi�o��3����O�g>�_��=���N��N��������'����/bp�e�~�<��.���>;|�3��N���d�L��!�Xa�8��g���	�f�m��E,�#��"7���H,W%�7�Ш��R�Rfy�l�έ&c95�e�c�3ށ���;X��w�11�D�j������>�E�oa3?�c������~�7���w�ܛ����#��^���(�4Y��ڎ�<%V0z}�,f�.W��
a��<��(��2�󤵹��*:��X��,X�I�:��оÜ�M2LsCj�I���{����[ ��l'diE��R�On�ک�`i��;�+~	�s�$���#�jB�n�U%�Y���yo��{ȳ�ɻ;g�qմ"�m3ݸ�}��(���Q�'�I�ſ��b;ϳ]�y���C^2Ӌ���[��/=���ҿX��kwG�k
�n�&J0m�;'�}A��;^Kk�ͨ��;8d�Z� �o��ﱷ����_��V\�̭��8���$� �@���-4W����9+es��4N�.�j�B�^�rg�7�����0���f�_}�{�^����E���1��+�C�_����L�{��^�i�͵��*N}�߭�0�栍�v��ճ�ϼ�f^W{O��H&��*���^ͥ��f�>c�Z�,r���\SJ�qV~���ۯ|�����r���������X�=2ݩ=�+�&牒qYL{����D�>=��a-�Y�)s��{T�q��9���-k2���b�BB�,nK��;�0ud���O
�Y-TS�'Jo�T�^�Yg�?6/;Էv�J�ؼ��0�À%��|���[���4N��ļRv�p��}��vXs!zX���+��}����ȟ	%x��FiTΟAз`ʒ��i�ڢ,_���M�����\W��Ԯ�SV�����sy�~��0�L[�7J�r��pۈ�$�`P�bK,x�%}��k)Dm���6`��]�%`�,$�@!7�@|��(ʩ>�z�?z�`h/l#0?v��g�U�����ʰ|��n������������,[+�e��"I��{م/?{�[�2��bwTV�ȍ���]�c�G��>�8� p�e�gƲ���"��$�k�'�Șr�_d�Wc�}�v����ǟ�Ɲ瞗�=��r<bk����FK�z�dGZ%f���&�N�U���٥93TL~����-aZ)��s��n9��$�53�$���Y��A��b�����a�������3��1P/�B)-&UL��D�;�ƙ��#�8�����9���-~�Q�"�EQIHbg��Zr�GƜ�V�[��C]Lú� �e�To�cܝu�bH{��J��,o��o���k^{_X5ܷ��Ե��3��k�~�Ϧ����~JTh�Ts�獗lg� 	^/����ݕ�� )��9�c�+ZZ�T���z��Ck=����b/�ѕ�����Zˊ|���l��{&�ٸ��J��㞠d2��v���1�.��d
���\F�a���Rn��=�s��@�=����K�7��$pA�0[�yf�秺`2�Y��lg���@�'U�@�}��E��jʎ1���A>��,�ɐm��c���ʭ
�n���:ҷ;��������C`^�!��8�8�4m\Tc�h�,U3��%��}^��QGی�����R����mݳQ�����8��L�Lt �Z1/��8x��}V�.��0V�1{���l�Ճ"t|	��U��	ZN9�#�!5FK�}���� ��\L��+Mc^�^���t�ya�3ߘ�G9�N,C|�{>�w�{B���S�!�4$�`��i�.�0#�=�Tci��Р��>��o��h���d��ss_�j����!�Nc�^�Ǆ*��^Ɇ|<x��h8%:-Z�Hz��$`��c�'��F+�:��������%�7z�-p�Zb8�K����
E��\jN���$w��b��L[qQ�5��ي"MQ4K��oc��W�Ǐ�	���j�˸T��K��;���e�~kK,�����U����5:R1�#vhq���v�� �h� ���h���%�"���'U#���_�Ą^���!�T�c�}M}�ha�Hrd��ᙻ7mPV��1��Y<x��Q �U]B�pHȚ��������o2� � j��*�&����e��. )`�Sm\���fX��qbڗ�!
`1��6�rJ��=�7Ti��<G?�Z �V��(�?f��qq�r(Ю��!�����ފ:�Ee9 fUVƃz�+�=���3�~��@�Ԕ����u��e��e��ᬱ�Ji�%+�+HP���%��I�Ӹmt����`��aB�gޡ��_$�����9��a<K�(����Gh�?xA�E�<�ن���>h^��AH'��p�|@zm$��e{�����=��-F���J���q��ߴ�d\��3Z�n��>
`�b����%��>X94M,q!(�>��8m�����7����ZV�䗵HBMֲ�۠�s�U�\<�0O)&���b�9�u���1w_h����ǧ����>�� � �O��${�"r�u^p����Ֆ�O��4�������������DLh��&�d~�b�m���Uc���B�f���7�2�$�£aĬ}E`�tJE!�P� ����!]*��G<T�x��9[WVW�sN���+�C��ٴ,��
�Jׯ ��l�Q�μ�˿:�;{�g��@�h�vwoB���w�x���F��@�o[�kK���営eL�G�x���#����"t8L?j(�����twy
��J�eY����X�h��7�(;�	����+qwo�M��~Q��eߞ|+�Y�!}s���Aa��4i�,[�* k��4��*�9n�4�-���<�IӁ ?(�B;��(�$Ovz��ؙ*��t����<g� �3Zw \�EF4��
dR�~�mG�f�43t�320��2ђ�s�=l�v����y��A�9@�R�KƛN�Y��z�?C:�.��r��߻��JQ���?a�{�&�ڒLV+7��>�:l��	q��Dx�5�D��G'�������nO�[�1ų��A#�{~߽3)TQ�����v�����{z�2�~:T�v������1�����h�K:�h@�g��ut(�k�0*�/8{X�#x�[�+P;uߘ�E��q��U��݅�#dzB�A�]��L��	�-��!�\�59r�@�+�1�7�3}8����rMXt6��.����[�0� J�Ql�3

v當��,�<�(����(�V�/ۅ��Yd�|�e�LYкd}p��F@F�D셵XBTI����KM%vl���hD�MJ�:x#<��d��ڥ�	^x����ĭo#MʥQU�P̀%���i�q~Xk�1��T�׈J ��/���9�� .c��$�����%S��)�U���Z}�.kh���{�!����~���>�c?z�vbq�l����Re؀��z=�gV�Q�1��=����p6���-��,c��&ƚ����QMP��G!�=�-�m���3�A�'H**@F�#M���!��j��ss�EԌ�4��dΤZ�]{-�5NSH~h��1pz5S�� i�x�;|�����;��� 	>J�d\��� �Bo��א�j�]��X�s�*)2zJ����p�>��c�,���%Y��]���!�u�ȌǛ ������t�T�HQQ٘�pp;���j�I�r���:��X'<1�5�2�򸛱hyC�i�8�W��]����Џh<��"�tς�
��Z����<lY����3׶�2�M&f�zZT�I��8�Z��JqD��n��]������o�Z�Ә6�	��?k��Vi���<ϸ�f�*9I��Eˁ��4�c�Q)'�d�$&0�)�T�+�$�bf�hs�z��1w���9�S�$�0A�����v�k���)�����l�{vD�dل�t�ˁ�4�p��o��ν�3�eE��x��pr�a/ͻ��<���&$�t
�܂͎g�!zW��S���M�C�w0� �{Hp��~�#�c�H�G��ڇju���mA:�X��.rex\��8�ň�:@�D�;�r�-.6/2������xKg�BjBƪ2�������>�*~i?�?�Xs&F{��n���;�E���J�zE\���؂��U�����=�R�y���wqh�Sx���	�X�s��K�%6a��p��PO�������CE�L�i�K��0V>	��1S�f~��Z�h�s5i~�o��,�L��F��Q������?�����K���hN�d2'�F��L�W�Z4t�9Dp�RU4���b�!���Ȑ�i\z��g��C��o��,�N����X��5��2����T� ����9�S�ὄ�v�hh'ád�AĚ��e(����	F�,k$,���
AO�Aܼ("���҆��8V?/#Qk�̍�,���z�$_5��Xw�R���W�U��N�o�e�}��N�ޜ��`Sv�.�;o���_� P��:��(ݳ��5bS~wW��@"����K���W���Ԉٻ�/�m��%)�T�k�uq&��y�ţIL���k]�a�S(�[&�����G�����ϟC�k%��$�\s����6xD�3�f�<,I�'5�E~��y9��q�a��LX��Yӥ�@x��7�UC��d`��C��@ډ
����d�)�G�wlf�֣	Z#��/p�Nz�3M�T��@ͣ��xB����Q�� �6��K�c�,}�
�l��_�<�Wz��ޕmE��{�f�x:��=�>�0I�rd������lf�!s�F���8��7ƒx��,��=�1�i] �R�!�Mҍ�i�W�U{�Ca��3 W�|	�y��V�0�>ksp�C?�<	lo��L�����e <��b՘�u�.��1EQ����5�WV����4�/!_o3��ƃ�-z6��R<V|��!��(�c��-|�t���\^�0��+�`��ey�b�U��lk�/}Ù��D�#�,��:�^�{��c�Bc5�:�>����{:L=���^`�:�!�2w����1Zn�!��~�R��8m)\pw����BWh��ɪ�ReY���W*���鈑��P�&/�C�j.�a��0�n/D�<��s
��9�	��Ef�U޽��j<�#]��ɺ�~�|�L�Y��?��k\�i)��a�����ҳ���C̠��D3�ǈD)	j�O�F�s���z	K�G����o�W�]n�!��c�����UZ���O�6v-j�*�
��dGa��!�K,��K�"�i���p̼��-�;�m5B=��n�Pj��6���|�	���&@�$I��x�Qs4fK��J �K��E�K��\�=�h��{ߪ9΂c@H^�.F~&I�2u(d��/1���" K����D�[��~��X-ɢ>�
�2�]Z�cU�"���8^��T�~�y�ʕ��?[U����Z��x��֌�+@z<�`�< C<��5YP���>+(k��L/�c�6v'p9F�n)�0F�I"�5���iY��d���t"ƓI�7#K�p�Z�Y���S�nF�R��U�<"70d�%�V��|n[[�7��I�@�̌��}�?����M�eNV�![z����3)�*����H����߸
*&���2�i��c�����|#Ϭ�3����$P��rC!���E�� ��K.N���B�-Q�Wh�K��v0ۜ�u��4�NyD����0� �c��#�7�����PY}��Q��B���(� ��qL�r�5_B�32qFv�E\O��ȶ:�)�0�"A���U'���`���iRY�aTeSj�TL�Xf�~QM���D'�%����&D���$�������Ғ�m�d	w�}��V|v|��g�(7��~,��o��s_;�(+%�r��c����[�R2���'^��[����q�\%���d�KT�E����f&��o	�ʸ*Y7�lK��G�L�/���ɯ�ˏ��i�ֵ�H1!�L2˝�t�U��z����/mn<�'����Y��5.��!���9Ů��m��v�:��A�;���Is6�2�/Y1�Z8MsR�g�t�Zq�{_�l�a=��;�}v��t�_�D5��ܟ>w#�޺g�?�1�.mt��� ^^U1��������ا���W���߹Q^Ȅ�UgB!�V�� ��3�X�=�R4J�i&h/� +#]�HvX8
��_K;�w�u�׼8i�S	�!��i~>�kGe�k�8��n��S�'�v�i9(�l���%k4�ܴ������X�����vv>�������W�g�xy`���,rz�~��"6�w�t��_�NvbA�����kk�mΘ�&�Z
�|����ܸ���q�(:�S��Fq�g�O?�/o_��[��J��t�²�0�e�1�E������1~�i;ׯ�>��x����'�%�:�>�����d$TH�	$X��!��zP(�F�N�
Xԅ,hѲ�)iI��in���s�	��q���}�<GJ����oX68s��_/�ʼL��U=��;ӽ�?�7��ջ���^��yȄ2�W��[���S��y������{_GE����w������<��T���ǐJ_��Bp_ �jN~t<&i��w% �b����[���4�v㻇�H�{<�𽧶���{T~����o~�����7�b4�L�����sT�������?~����J��$zG,Ϟ�q�a�۳�k�J��R�~K�_nK�>`�k���½�`���M�m�A�lߏXF���Y��=Jhm����۞p(h)�%�>������:+�e�va���^{����{�{﻿�T�C,�ܿ,gu�gQ�������ϫ�7������ɩ�[wd��r�)S��S�U�daǛ�8��ET2/�^�]i!Xu+i+�e,�����$-:��%S[g����>�;��G>�����m8.ϰ2��	u-ǿ�m9T��w�1��/5�wn�f�q�;��~��`���*�v��;���� ��#+�o*
V���ƀhʝD�C�S�pw@N���w�Ue�MM����!��k7 \"8�'�8��a�#�!����o/YyU C���H['�p,E���3R�R��`j�q6���r��_۽�Dy��co�ܺ�]��I��KD�7�V�������>��>�;��yj��7Pߓ���2�8��}�&/��* ���!~s�&�Xf��!K�~�����)���~�4Qi��.5F��#���-8]��}�aw3�K%�M��)�r�nb��,��H=���G��7>���c/?����On���̄���Z���U�p���w����=����u�;k��὿^q�����\i�"�0v���d��8��q��C#��4��p0j2�)>p>ǚ����p�ui��B�L�/�bђ�7)�G�,���YhRK�TO��53�������������g�u|�ƫ��(E�	Ne@�)�2�W��Q�x��]�;�r���`3�K�_���9���3���R��=ԁ�w�5�RP�,ZB]�pKkB)�����TOX S�@�L9��-����qXV��x�_�^�YUp�gN�躈���N�u�o��ON����e�Ϟ��={���B��YCc|�����9;	<��>h��e:�����x��_��?�����ɯ������=���[�:����cg����2�3�r�8�P-��� �e�� �R�0�,���	>5���c� �&�����^
S0 ����6(�0�1�G��ّ-�5~>����}��NX��L�ܯ�.G#6~y8~�����+G׾��ɍg.ƻg����V/$3�~e̦7���y�ޕ�*�_\/��&޼돢d�L'ꤑ]��� @����Q_i�.����@����Y9!y� C��]Ƒ,�i�	]ݐFƀ�	b$�淄m��jx�1	�OÒ>;�=���pPZ�����]m�b qw^M������'�b����:��O|o��o.&�,���M����P���ݽ��"7������������Dot؛x�;3Ͳ^/Is���q��X'���~R��8AK`R: e����r(u�4X���zdi
.�\Hd��q���9SP�c��1 m��Ŀ]mz{�1p2�YR�I��!�n����;X�T�gh�߾G�����<=��̧';O�oo���/�#�ܻy����O	 ��^5���m�v�F�}��}+�i>�W�wџo�ѝi$�U5.�/i5�vX1@���##W�qP�Ȉe���ڗ�j�IҐ��,Z���q���~2c�JKc���+������.��y]���o���yV<*�L
n��lzs;7��Ve�W�껮���M���s�"]-���j;��D��⽇q����,�	�Q1��5�j���7޼>������_���_t���qF�n�Nb����Hg�;F��V1��$�V9WI�e�U�	�G�JW�LI�2��j�Dne��అ��(��,xa�n�n'���NQ��"KLj�Op?e�B�O����������C'�s��O�Ԉ�0]^*ˣ�d|������>�~�o�{W^����`/SZ��v�v��5�<��r|�o���a��Ȭs�C ��=���`ŕJ�c|�ki��:��\g�=a��ʥ�IX����"U��h��9ed�*��Ov+��-��G�E^�5l�Q	��rd�_�uj���h���-S3�}�M�x(F�2�ݾ��S��M6��]���sB�AtH3�j�_�u�o����c�K��4�����譟�XF
 �m����R�*/!(PGѹ���2J���

�)��^
���e����b
j���R��hb@���Tl�a	~JX�ܛ�cW��Η®���j@+���@�@����Z��p�b�d��]@u��9+����O]�z��{�S�w��G���o}�0U�F���ߎ9Y��׊��BlM��o��<V�ݵ��:iGUe��1C,.�L�n���O����[�{��o��{Rc��g����s2�����z?;����?7��V����mWt�krw�n,u���-���U��1���Mc^��ED�������z%�{~sZ���$x8�l���%JR��p\7T5�:��>�=��-�����ɩ�;Ig:H����b^�Z5�����]n�HX`T�P0���e"�7�6�"*�"� \X�5����p�!9Y܁cϷ�$2����T�Y#� 'ŝ?	��n��<�'�WLF7�G;����]M C���0�c��ɷ�{������������׭�]������*���%���ّc���� �z��md�(0#�����ѷ r�\O��sJ���G@�?�k��.KS}��1fd��ȏ�`���.����Z���U�1��{����b��v6�X�r+�@C>e�R>>3|�K#��y]We��5��7yu=*nU��'���	Ulr�%���[4��]�v���X���m�����rq��Ue���#��T�=O5h�BƦ�����YF�Q`�]��GU���^v���o)WvA�t�G��P�;v@�=�3K�Ͷ�"����_���^����������;�u�;@BX*Um\~���ˇ���N%�g����n��� ��B��@{��:G�F9�%|�a9����>1 ������!�����m�%9 \-M09��U�0O��h �F�D>u�<���\d�,{3i%\���s-��ɲ��N_9�촑�Ğ6��_Z��d�NW���Q����äxm��_���{[zwo#ۿ�@&��Dv�-%ЋE�@�2(�o�J�Z�Ю	Gg�E�K�ƨ��o�~.f�Ep���m��E�k����9j��qnU��X��T�8K�1Z�8R����c�)�7%k\�yC���K���;wO��|��72[�.6)d���`Xä��l�@F���%��\��>UY���>r��2jt�����-h�`Qq�Q�u��@����}Ȯ���;>�HO��C��ɨ�v�N�9ƺ8�  ��*`��/?���V���k�t����ɫ&ן���N�66J�[��t�Qh��f׼��SeW<)-��Aħ�Lj��v�"� ��K|`��,��M�If�=�dǱq���م�K^�	W,Voۿ������ ��1o>$;a�쌳����[ݽ������sI��&�R	�2�-	���/�6ѭ�<����;�������^�j2|	�D�ۑC��D, &s�*��tdf�Gr�ͯ�hf�ǡ�	m���M�����������X.4�
��Qj%���� �AJN�!s�h�6y�����]��l�M	�J��+<ͽ?s�`�Q,+�u(�̐�h*ˋ�5:�|�OfHR�[w����.ز޶�k_��Ο��^�I�et�4ÉT(U��io�6.~�Z��{)6+\Mؖ7�sq��T=vV��(������D����Vz���̅����� �0����cV�DP �yd�)���R��)s>��|g:�q��u��)a��&XJZiJ�c���*u�]M�p(Ԅ�zE*Gר��%�������ӹ�E��_��C�2�?����]�]�s�/T�R��bM��w*���kB�#���RU�U�q���.���`8�\���WI�2���z�E��{�SK�^ p����ȍ$�!�'C�q3�{�x���H%���k�dT�X�T�C{ul���� ����h
luy��V:��3���\o�]�6x����Mk۾�,9�������Ls�5 |�������9�� J
n��Vơ��9�q�x`Kf�:1�u���W�jG�����J7���Z��y�Y�{{��pǔ[8	��&�=)�(8��̷��j�R��8��K��Or����<�t��*2#�?M+����}�GT��������/>�搋nR�ۯg/���K)���������V�ԉ��C쟗�����W:���5at���ں-g,�a�|�5+���=F�S�/�XM��v��k(��dQ���E`v�I�w@m������!�b��zz��Ŋ�~�����Q}|5�ٶ�a��X#`�6qԩ��@�-7v8��ߎ�����E����S༌�]P��m��qh{A��ޚ�TKn (�ޅmF�z��q���5�&�mp� �͜�PK�E�*�������L�P���K��J��"��~�GL�-V�{Ԓ���L�4��گĆ�rc:���)9s���1����dNtnL;3��s�)����l��z����?^���_ږbѬ\M���_�J�����3����v�6�֊�6�y}^Ô���q�l�Qu��/1��O�~/�$���Ф�Κ�����> ��,�5ˣp΅��`��R��ڊ���hR�s�E�h�1��%�︈ ��^������WW���I�+�]���9z��3v�im���yn�"Z�_ʦj��aS�Ԓ�T�~3������������ʆD�P��6W��3O�H���&u4s�|�J��B�͛��x�<ޭXKj�c�ca� ^�h�hj<�>��r��n�~�`.x��2wi���`�+�������~����>`�u��W�v�5C��Rf`6�6l�6We�c�$H.}ۿ��QtZRoI�l�z4*����,M��h�=.�y1�틷a�E���D`�����������=�4q�(��v�:_J��7��Ŭ-�O�&[�>��ŋ���R�0LRJ	�V��K�l�aS��+P�)�I����
t.�M�r��H[l�S��]�7os�ǁ�$��<aY�+�}��I�����/M4F�o.T��<:�z:)/f�Ӛ�%��t�1o4�u;K���Ͼ�+�ijn�������$��̜��c��qN�c4��iOd��1d���[̚�׸R�s%�U���I`�8	��(mfP��w��vЄ�{���l�HګlkiG��mٴ�7�]p�~w�6]m6��^���Dp�j��U���L3bZB��?����U}�o�-�]��͎�a^��L;AͿ�:pn��m�gP�7��`���,�_��@�QQ����.2���ϫ�JZ'{xiOG/o����ےLV�����8M�L1�J^z��cZ��+�6NT�%Bt4�l�c~b����h��a�md���cl֫�C���?��S9\͑��0��dyB�Hd���sX&��v�D���` s��p��j3���U���j>�[��"�3��Ϩ�Qp-��PjZEI`U�͚��L�����$r����8����V̕�@9�%6���+?�bF��ʝ������!( W�M�L�e�N�»q�����^��Bu8��2�/��k�*�xX�/	&�Q\����6)�K����D4i�hp����l�FRu�%�%2?i9}v, -]J'2w�T� ��br�Z?tQ�Vx�9��7g�	~�0�c�G]u�Ā��b�����h�`M�{@�V�X�	�n4h{�*v��g�,�`�!�X��p+�չ� ���x[���s��a�R=C"iv`��8�Zj�QǷ����yƙ,}]6&������P�2��L@�*:����҄]����p%���+mu��F#b3�����`Yɰ/�]��ӅJ37�h%�\i
�wz����1����������٬Fۼ��;��*'q���ڍkw��!�3�4��cJ���O��k�ّ�}�8��*����}�1I���QR�qD�ؑ 9.4�}��OK�^�����ĸ���@�L��n��T�̓;>'='���xC���-x�֍^��� id`�AX)\pJX6���,} }Ɂ�bEMx��+�Ry�T���q�P~�]��v}=!B\���ߕ�m�E��q� NQt��m{�p@�h��ɾl
�}+��� ����%�0, �T�>!d����ax�[ ���a�2X�lF���9��ӣ ��'x\0aHF�5@Z���7��n�S	D^斸F~�Ȋ<�_22*N&^�d �]����&�uw,�V[L]�g��ǑL�Jeff����`��s̉0��v�[����k1���2�+T�, �.H���~�,��K�V~H�}a�T"�TFeb'i�dbc#�i)J$X�.0���	Iw��l��'.��r�$+��)L_XW"7A��d^��h,�F�q�nBp֕�>�X
�@��"��#�Q��I�� �;�b�$xi
�(B�Bt��*�����1y��h��ҕ§��U�]B,��*�c�n?ﭟy����tw�̍~om�U �¥%1hyV�1��	��:�*ƪi�rL"�0��\D��4��@��� WҎ�������iP�K��b�.���)�8`�*) O�,BWX5�I����y=��} �� �B$V��%�;�@S���t|�x|�|1ھ���M ��r��Zk��;�e!-�Z��[_��&iw?�:���>@Ņ}Z���B���%�4��Y�
@�C�%�#�/�ێ��D;�h}�$/V��J#pT��U�����{h)�8H���X0�gx� K ����{�Z@4�v���:$�2��˫�R��RFì����t5�u��^2��_i�gn9��3����%��A�~�LGE���F����.y���$i����̃��I�o���f�s*�N+�����ΰL�p_�G[��dL��Qv����J`�Ofui>�Po
�xZ�`\�2q�@r�X� ���WY1�����EҸ���>�
,N��X�#p_s��̦��$y�ߋ�܏�m��'�b2� ��R�GQ%,����Y sՀ�%$�>%&�5ʩ��DeS� ��-��B>)��������(��(zX��2v*`U��P�
,��eZ` =ގC��؋R@9 �6���'��[�J�F��|zz�ͥa��T�;���p�~̚�X��,��Jk�*6�UnDU .E��.p�8Iʤ{������8w߇ַ.������g���0ʳ(1�4 �I�M�2�;MJ.
�QՉ�+�K2zh�����f�0�;
0�',�q�[�cY��NR�	B�}up\���$��%"�+�O��U�!��L���磊����}�����ߖ�]�66���x*�Y�x@�D�Z�(���/�S�h��_�=�h�� �Σ��sX�k%NxN��i�dub�]8�9<}��o���s�)��߳��4��*��$��J��O�JL���o+�ш��,���G{[�;�|]���w�����j���[af[ݸ����V�*3�^�u�s�w�sBv���mM�(�% �2,s��J�:`Y�� )�~pwGԖ��ci�!�� ��b�Y#Μ� ���3ueA�ߖ!<S���a�FA�)��:�(��jڂf�%�` �%������xxi�}�5��ƃ���T��J�U�'T%�F�#�f���H^9�v>u>��ʖ�zlڑv�X���&��{ �\z���`?���}��Km�ۤuN��=bwn�Ι�������y}��W���ox֋{7'٫o��ﻮ�����V���պ�����
����f��s44�&�w�җN�{�{{����w��z�;}�
���jr	����{d��u�r*1�`���N�&�8Zg�q �RQpVRw�m���!�^�uu/�y0]$b��]WH�`�C���o����+��5n�\A��p٨�����O��n��U8���G,Eb�8
����
2w�'�����78�U�>s��O.�E����q�����'ա��tQ�L�ż�!��N�P9�r�2!���B��裾N�jy��� ����!����R�߸��ذ�ъ�:U��br�J������=2�]S���L�O�����ow=D8b�2�]���_�����~��y���rP�#�E��q����e�7��L��C'��9`����9ǵ=�V�j�M��
���`����[1�X��ļ_Q�n'�;�W���Ͽv��?��<��*�;e����~�r؎�^�R�J�I��^L��?���蝛������{��3ᕌ��ꈠ�źD�ͦQ�"f
Г\�~&��
H����O�P�d"T�"qK)ٲ���7/�Ǻ[����`H4+Dr=���7��O/��:��'�8�A+3��4�i�Nja*H����_T<���~�N����0޺������ō�_��s|g�s����g%�Hi(�!M�}��&�� !�7��Z���/:�k���$h��Bf}��q�E���֮6$|v+��t�P?D�,��邂��$�����1�7P�m ����-����4��/�;�r|��Ӭq7�T)xrZ�t�Ι���̥�}����p�{�e�ԝͷ�\� �,��)�`��cVIڷ�[WM��vщa���x:/P������1��|�ܡ���>��;��F4�Zz�ڥ��hlJ�3垨���N�������LR���W�b�[XQ����	��n9Fg�������������k���5�w����/�{kq�*J����L/,��Dc��^���� �'�
���+`l0Z�`*��
������V�3V�3���19�`1�-��
�V�~�P'��҉�-Â7�J�X�`��[A����oa�@�ف�9"������go~z�y�c��ͫ7��6�7���j�ׁ��kc�s6��t���������I�����+�;����J$\�����-J���\�_�	�� �8r\�sĎGӔ ��6�jΖ��^{_P��v'^�0����lqh�
B������&Y�I�Ci�ܹ����X�{����˽���x���B���8��9���x�%YWo'�d��p�1�e�?g��O�_��C�g�u���w�GG���M���C�De�yn������Vz�:��@�9OY�H���w��1A�T���t�Đ�����{���pQ�G�Je�`$4��"��~�X�U�Ir_z�{�i��ộ�~tR�6�Fof�tv�ы���g����ŗ�Ʌ���q�փ;d_�g��J䖃FNP��)��M�F+U���eV:Q3q�[(2n�IW�s9�������v�GZz�+���:s+8�ОR5!�Y�o)�L7�}u�./u���3�۟P���SN�����5,7A�2�����,�S?�=������S�����N��i���>�l�
,�a��e�n^�X'����#1��S�6���¹f�D�'��$���9^�q��؀���4��S{�elvp�2(^.
}�쩩лwO��=�������G��U6}��t���y]du���������%��w�����;���%��k%�������E��	3hŊ���@�A��*�#W͜@�������6�;�����P�I�٧����v�-��v�Z��K�6�%�~����m~�������T���Qg�*��C[K�?���Ҏe�E�P�d�?V�&!�w�N��>�����}v����s?zK��v��i�%�A�8g�q`����IaD�^Ϻ���'ƣ�C��n��R g{_�!Z�[lE�[8�̸�*�Y'�U�ޭs���x��������]}o�w�>�".1��H�vi�?�nl�n��]�޹�~�쬿��T�ߵ|�	�+�xb�0
G;�����˹s���rr��;���]7gۺ���V���7�q���T�Cۿ�H&�r�u�N��o��3�t����rp�M�p��&/�(0�4�K�h��#kg���":w�k�7.<��;f�f)Zϊ������s����Lt�7+�ߓn�M���n�c��uo=�x˩S�F4�gk�w��h��Χ�ʽ��( �II�#�@���t}-~�z®����O�����7��ߘ��1XZ@��n�˨ <>�sJ�s��5-��IPrl�;.I�_��>�yf�U��� �v��=}ǫ~��ީO=/�<���:���N��sAx���8��J�3���J���B���M��(���`��=���?�3�'��}[.ߠ�����7b�X�` w|'�
�t�i��^;�}�x[q�m(z-�([(qw#6���*b�M��y��o}���O��������v���K�������%CF7Ez�s:9}���x�\n^ء�̹���m�Q1�|p�e�u��勼=&��5,,�V���N��l}���K�����}����Gw�<;�/��^�����d��m~�'�������C�G�~��[�*M�]�Ե~�*Y9+�����������Nf���[��g����1�v|�L�~o��O�����_~�ՖF��d�CƛW`ø�|�5�sݎ�t����ѯ���}{4�Վz�TIPfuhRv�����.j�ΟI����	.���!;s�@L��ؼx�m?�w�������W��o쌷�E�ƛ��L���n�V[ߎ����b3]�Lְ<Xx�������Q/br-�ܜ�A��=��&	�c�Uc��Ɖe���	!b={����(�3o�(<�֗0��m�}0��Ip%H�X϶zk,��ŧ�c-qR����q� �#Ђ��QZuz��h�v)�C�)H���JӨjPS�B��aq�t;��q�o�o_n=��+[�Ž^�CPK2:�y����.p*�q��8�f�������2S%/b�zeG8&xH�C]������Ë�Kͤ���J��B��ٍ��m
��p�������G>����ᶩi�chD�M)�-�
��*�S�%�T[	��*�GA�eD���bn�y��n_|��hg8��g��O�,��,�*�Ԕ1p0��XZ����*��R~�T4�D�$7;7��&k�nn��κر��L-񠜱���?/}DF̬��v�k����CR�|�a[��cN��j�lSJ+u�����	�|$F�um=����ed'[_r�ƪ��%�B3�R	��:B!�z��ǥ?�It�"�2�}�W�ؓ�b.h8]��Kjɓ�W�7��M����ynoz��v���*r0��4�K�s�39�Do���
�m��.�&fE�X����ݳwt�CX$�J*t�n�d���Zzƪ4l�7!���%��<5��������5n0��[|��o-?�}m����:�a�{P�f���MUMY�M��Ǎ{w�������O��;�}.�q�7���N������`A��p�L(�F�n"��*d��I��!�q*�T�V�{�yԭ}���-T��$+�z��.��N�s���w����K➝r����|���&�'XS�����]���X�Y��mF�ch�#�����Dk�pu�nʐ{+���\l�����`�jR�R]0+0a�Tl�e�;��^>l�7��_Y��tgW���D�[v�rx����ɞ��� u��^�����X��p�a�"���n�݈�1��2�0T�.6�1&�	��uȠV�����v�A�����{����;�Ȣ�e��M!�ft���\��5�VhKႻ+��
����?���LT34��M�PZJ-�2�%3���9
���>�c���_I�ո�w줖E'	�N&�o��$���6��(^C�D�91�?.tT�
���P�A9����_��6/�>l@����e���~�!#dW�1wឫ	��-��O��������N�>,���i��dx�1�Jn0��H\eS���u�xuIi
���˙������W����d׾x!�mTv����;:	��pIg3c/�l=�]庪�{r~�吲R0~c8�ɄO��Dv���p
���U�9,h��8���x�C����a�OY�����33�x���|d9|g0�U�{���W�Cv�ry ~* ��.��vbM�'[G����N
 viIf^m� o�N����/+�
�ۅI�L�H��P��(��� J��y9�����E#�%���F�c��K9�̑��&	��
����}��:�� W�1
3�k���"b��w���^T�̛X��$� ���.�	b\$�K,��=k9�$�eʎ�ӌXgX�8��hj�"?�Q� <p��P�4�Շg�QX�!r6������H�U.��/�,���B�8&ή�M'Muw��յ]B��5G��r~ !������
~�r�tp:��Pr�/ [�={��)r�ׄ������,�z��]$҄$M+�2�~��2A�f��"-j��Q��f6R��n!�&tS��Q����S�4g��}�$MYiU�IY���h��)Kӎ)ƙF(� @:����f�Vi�T��
���{�1�𽠁�:��f�T��RߥKD�8^N�����"��]Ӟי�L���8tN��V�s�f�-y}#i�J�R*{nfŨo����Ys;�"#u�_[�T��;��ʡ1 F�;v���i7����2��_�y�d��3��7�����&�f15�J2j���\��=�Me�1[f��Q��A��l}����1e�����i��b;~
��ϪV���7K8!�Aڟrq�,H6
��AcȤ�.��F?_�<�;e��^���Q3'�4���ف�fˇ@��Ȳ�)QQ5w��'�V�r���-�QIBB�3�z�i��X`h�l_n���NV��������۫O��[㐦L��1+5��N�>d��&,�^��G�;g�E;�Gq���0���y-�ڿsI����cn,���PV�B�=��
��T�G��?�7
���Al���>��H��j'%�Ѓ.�##�V.��cZ�!̈K�
*�^2F�ɩ��
�8�2�����%�qZW��C��..޾,D����t��~P�.�7��
�-)KĽ(gC����b�n}���p\T@���|�����4uH?�B!R�r
��DK	I&����H��W�l�fjRK�gR;�
 j�{�_��d�`+v�0t���`3�����x�!8��lXZ]9�g
٭K�#�4���ZѬ���"e,��ː/	,b�>�tcD*?��(�bͲ)1Q�Kz�g�}��i��^���H"���E���Aj�����4� �J�R�D�X�쀳��&�=��}�0ў[]�Q��\�(	T�xS�1r٣9x>M�n��� "53�;�� o@`�j�p%���Z@cNAj;K]h�pn��n yUs���OI]K�����`� ���$�R��K�&�J;N0�n��:��M�8L>��:0�g'���ۂ�w_�Z��L[��NڬQ8�X�t��gV
���j #�[F&":W�[�$�h�m�,J��
@� z��$\Dv�D��Qܲvc���+�u*AO��@8	�b��d'G���(�17�SM�:c�%��k�obF�M��L-�t��
s�Qh�]�OՋ �cDG-���E��6�	���]��]�{�%i0q��n��?b&/���3�I˔Q,����	�|���B��@?�Ru���R����ODc�1M�u����0��;3"�i�K�P�r"@@���*"S�(:�>|n�>.���Z-�W�@��n�sc-ʬ�F�#�jɝ 8R��*"L�Uk�uӍ)
�QL�)�f56ߖ�[��&��akFC�t_�d�7S�07�Nx�H�}�������x�5蹤`V n��p�S@<u�u� �	�>�:ު2ch<��\��|<�Z��{Ɍ=����Ў{���S�M�lÇ�[Z��l�0$\Q
������3�C8)�b���%JE�& 0T�g2|��]�Y��Cm��0F�hN�B,��^6�#���fuT�Y����[f�B�!@�OC?�Ԅ�*�*;&4�^��d~ X4-9����"�p,�u[L?�q j�	Ҽ|��B���j����{zs������ǿh�45�X�n�@�������7Yе$��ud��T5~ �0�
���an��.������Ba�v�f6�@�TV����V,~TMV��7O��G6�� ���h���<3�L�c�}�ɕ�\It�Y���C:�]iK3��ݰu���Y�a}�h@���$�TWh�0x�3���� U0��g����Q�툿�g��I�$�I�d�	�k�V��42n��rNR��<�^;ڬm%�R+��q��KK<��o�zh1w����g�i���.kA> �R_��ރ���m�&�fhv�P�߈eb���-b	��,����̊�Wv!��|��K�UXL
�P�]2? �kd��צW���4�X/�О=�Ƕ�v�?���n~��e����2)�@Y��i��"����Ooc$jkG�����3S G7`���_�8������^�w\�Ѽ�����^�M#�>:4�!�h� l�"�w���P�2�"]�Ǜ�Ȝ��u8<&Qm�#a�d6L�e����/ms���s�mf������ۯ�,�֭���A�"o?��A�KB È��9a��Y�v#�G���9�j2��R�FNG�LӯI���C�p��`%P�$8v�i���#�f���I��iS3h\�d�a_y(ܞS^�u� FӬ�:G�E�q������^`Z��A6eD�M jU���X�#�m���ld+O���G�����¾d��Ċ���>3���?��J�b���<ʨ�h��3�ܳ�"�1Fy�@�L�4���ߕ��юn�ԇ����"�ń��Tm��Z�Z���J/��EN�q2��o��	�塺2ǐH����
�DW2�P�C�!���jT��E[�bb��߀�M�E�P���7E��E�7�	�V�z5|	�^�v(�wIJ��PV&�:=|1h�R��S.��]�른�W@S3wR�U %�<
.��G��JpQ�Ā!w�ez	^ �U�W8s��a�>�-z�P�%�����A��Өw,�f&��*^�n>$������8q�!H����nL7��MX��XR:���oP��u�5�9X�_Z~��/�J�y>�Etl;�7�1+s� ���>�2?��i���>�+#IZ)�2�eG�(�p����O�
�)m�|9d��I��]��<r6�X�V�8�1������NmX��ξG�h�cS�F�y�&��l��V��+�Z)N�.��uM6�0hϰ*J��#�fS�����J#��� �#�#�C.�"d͖Tt]Y@^�=8Q�"��9�X�0�5TO^��W.��J�<�������_��V�j<��&�A�ڪ����Fb�x}�B���k¨�jx�#(���q�%	�0TR� :�R �-�Hs(�gxf�_�[�L�y�����ݽy���`i���pQ��ś�ڦ�yM9�o%�$
��wR �� ��[F޷�8���MF9���J�.DXZ�A�Wt���&��AlT���4����1��T��%X7M�R0������ߚW胦0�\���3��"Lp�1��ߨV�	 p�d�pyV1
`w'���MX�&�?<4K�4�Ө_�&���ȏ0�	y������d�WQd�E�3�K;u�W��� ~Tʪ\d0c�RV[JzL��%���Q��T�Ci	���qU���`�8[&�	�<�4X��ʹ�x6x��<���{������:`c�v�v5 �	8� �AȤ/>A6rm"ɟLS�#�r�r��>�'
+��	�kj�rQ�ɷf��v!PV\OT�c�1[�TJ�^S�]e�حe~l3�Wm|��m�hK_J{x!�v��Ϗ0x�V�_�Oof��в�b���k��?b��gtU޴bRE:�*y��:_�Xt)V�R��(���cNR��g.�ѽ�*�k������"O��	ǒC���@ܺ�$B����şs��5�(��F�ƨ/��NL(&�G!��P��-	��ZL�@sc��Ǣ2�%�VL4�����;�Ì�5MGm�J3�n	|��z��Ih����
"p'`�7-���C@=j#�M-SB�ZD	l���:=��~�����l�w*}B��c�ǖ���?so&�Q݉����V{w�I�$!	$��4�j`<#c<l��a��6�3����1�ޛ�g�x,l���f��f� 	���꽫k����✈�y3+�*���ԕU�7�7��9�s��`mem��J�F��[�f�<G�[��OʼS�V�u��.<eMPQov2v�S�6��{�Cq�V,�m�z����"!�g���q�(㴅s���,���bY1X�����zU1��z���z�殒n�9�U���,p� �FE[��dX�XQ7������DN���r��+�J �-�-�0����f�(!^`Ǵ|V���Z�S�%(�Ѓ�$,�;ƹ�>�U�۰ТRjN�r�S�AbÊ\��*.W5����J o�=�_2���a�
]-����ߺ����te�����T>��Z��۫��NL�@^�Qs�ĽP�j��1��x����)����g��:��_��4e�V�3�-�Iw�Q?4�8��+�,&_X��q�)+.�q���S�y�Z�#�N{��?���v=��~��Dg)�r���$w�3O4�+$���dճ�W�V-�z�V�9e��S"�z�%�c�6��>��_����!��A6ؾ�8Lj�N�c4,����a�d��z�WM�Q�EE6d��#=�[��+�9�l����w���W\������5{~9S�JC�����^�C;�.?:��������:Lj׆\��/�V����/	��ۻ���[�h0�Q�J�1(�:����$����C�jWi�|���>D3t]+�PCʭ9��!��#Ͼl�[�y9��i��7)��Å��˒$'ҳL�0�p،p��:5c�����$�;�8�
ʏ�7�S�є�*�p�&^�p��+ִ����%����ҏ>��3�m
���= ޽�jBg��k�5���Ϳ����W�[���/���k�̛�L^ZeU���:�<���i����q�	�tc�Q�
����
�a�N-ՙ��������(�Wz)a��U�!S���r�9T}'��ُ���v��}�E/��@wVT��s!�X��A�œ����;�L^�$��e!�ћ�d�U��L���N�bhy����l�T(9���\P��Ȅ�e���g�Vù`�� �)�XBrE�7��-�x��@^��+��oǳ�<
[j����Mv��n#�/�1�}��{�w��]L�-	T\M����Sm����g�~v�8�ּ�x7���q�s0�z�!����h��[�K��9���G���(��:�D=���5�$���)�	���jv�7�K+MO����"��Y@�Y��b-}�#����W��#D/�r��;�߅A]"ӏ*�@��/[G�~s*pDM%?zڙ��=��m߿�R���5��7�?��Q{�:�5�@T�D����Yu�������#^���w�S���̫^���˔�K�WE�4zOnt��x��rH��X�T��rvh����4M��� ��Ԗ,{aJ��#"|_T����h<�B�5��>K�f��߿����o���΅\o��,�����Q ^ԅc��C7?o��w��n�����[g���Zɝ�&�����a����6�M!��~e���c�h����Ms�Mp+G2Zt�	hU`�L�ϟ0h����qn��+����+����W/3v�P7]����s����_4s��߹��&�p~�T#ϥ���+��l?|�G�9y�\8z��I�%�Ʉ��f���7�.I�i��dC�mE��%v�[�p�FmP���#�NVz�h-��$)��gR]}�pZ_�hA[�R�����,t\M�<�g"�"m..�Z�s��鼪%с��S~����T��ɩ9�xW�������������k<c�cN/��M*q Y���;�N�c�ݺ{��P��t�r�p�������vi��D��I����������¼�7�g�o}YX9�+?z����Vr��x5�9�p�����\O@,�0۹.�kuH�r��{'��[�����o��`|Y��q��ņS�a��m�WJ����7_������/��\va�7}����sj�{!?7Ϣj���t��ٗ�#���9p�%���������	��֛)�#�7��q�(�����D��ֹ�#�a�z�8W��8����S�[Q��b��R�M�S^BMO���:�xϹ�?��s�c�^���o|����{����?zͥ���}��Y��C}K�5珪���Je"�Ƀ��֭�ǿ�?z:����k�,�b�|�Z� O��B����"������c���V �C���_��p$�Gő`hPʉB#ORR
�C���tg����YB)}4���"y	[��yʑG��%6�r�|ު��?�[T�/����o�Y�����G��
�"���lԊ(��i����}��T ��k3W{}��*r�Lm9���/�Ŝ x���n�wް��Wwb/@��B�Uu�7x^�}�gO<��u[��Vȗ��+U�S���m}=,2�kPe!����=����i�? $�[FS�]�[+����EY��+sJJ��4�ey��^����Ι�G����W+�ޑ˭o�Sw6m)��
�#��2x�ʛ���Cp�zq�[rA�S�.���<܀I(:�pMR�����ԐFQD�˓��;�u?�
��^�jqJ���$;o�C�dvög=�sn�1U7��}�����3U��J�:��Q3���YT��=�3S��#s�3�[�rר�<w:��w��Y�P�3«2��i�Qe-21�{�0ӧ�m����W��w�F��4k)�5E<�&Cf�B`d�,OtF�)d|k	��� �$|nrZ
cFb$��XL�!��(~drv�Gx̍����zv�O��K+T���Ua1b��ܻ�~��Z���0r�G�:YǄ������l@/O����X����O���ު����5+���VT%X�=���z!,tV�z΄�DF٧�W�{���۫�3�f�� F�;7�u��_�eCz�;z�#�`���C{3�R8��ң u�<k�r��6�b�h!�(2�q�I�Z�<o�o��M7<�})�~;8�ߍe8st9��W�A��;��.��U~�u�v��|����}L}��n~�V���fr %:W9�	�M�,��:�j5�r,�C�������p
���P3�Z�*���ϻ��[Ͽ����|s���u?���]�C������h�l�n�Ѓ�'�Ԋ[{%b��S��i��O1��L�ku�\�S�y��BDq�ڪC��=�M��n�ƈ�3ZT?����/P�"�Fh������;6z�����%̘ΆV�S蕰Q��퐭�尌�*u������'.=��&5����Oj{BVݒ�s��Vsc��R$�Z��W.��Ȗ���1x��Fq��So��b�)6E���H�#�,���;9�4h��2��D\Sd�>杨���v!+�Q��j0�D��9�� �ia�=�%r��'��3���%��N
a�C]���{2�h�s�p���q�Bm�F�8��3���~Q���A����Q`�깷z+��Rz�D���zB�a~ܯF��JX9�9U}��NE㍭ę9�D��*�����w�9\���v^�W&��Λ���:����mt+���]؍�������M� �{�c1�1�l��)4���!��"��a4�"�LT��D�c�j_y�-�4�!���?�ug���D��k�����\��^C<���X[�&l�HD���G�`�ޚ� �$$B? Wk'�r6�QN�Ą�D%��B4����S�F8fFj�|H��-t�J�.@j|����n4q�2�N*��i���h�To�r׃'꾳����4L.��g&�rQ+J�	/ ,�Q��pF���MQ[W�k��U���uU ���H�R�X%�W)�=o�m�8���%-w����)����K���k�a �� E���+z��q	��"���@vS�^ �I`���?5ÐW��u��4(-X[S�8F�zÀt�Q"`�^���.RX<沴��չ��.BJ�L댡Ǥ�2�v2$��Y�¹o6Q�������.gT40�Iϡ�Rq}�3�>���?~,>���5�3ډo��\ox���rÍ�Έ�ҝ'/mu�<����}׿�5��'�J��;��=�5~�&��������*�g��1���{J<�L�w%Q`�:V%���V��9��=�	X��[�[~������WM-�kpbJ�R�AR"�NI�S�e�Խښ60#2U�J�H�ZZ�W���F������d-b��جYW�-=\����)���S��c
+-2�e�)zH~)$�
U)�q�I�4���U)����9=C����֭��6��L�oMw����4���c���}P*�ӏ�N�)�Y��m5�)���8��8��Z J+f���p���X׸Fł�kVǄ�Ђ����ʇ�0�$~h�F����@�P��"'���nI����I�j%q�&�Ҟ��>��'��C3��kH���@g�s�>�i�V7�7���_[�ɱVC3׵�׶6G�k1nDC��1�nsu�����ݭn�A)��,�'XP�d�Ҽ23FHG��I|�B4P�vL�=.	e��^A]�=���rϨ��M9���q���m��}�bW�d�.������ʑ�_k�zbi!"r&�7v�~쑃uݧ�������bŅL+!U����˟�/�˖d]�)��|�R� i)�5�a�*��u����y N^�W���!�_@����w�Xo|���W��|�6�K���]u��G>�q�u��qy~�������:��ڦ��1--���l��d9m�p/x�8erR�p~��+�?T���o��<cYO����FĿ�S���f�~��b��j�a������D�n~�OV���_۽�_�)�g�<g��j�T�F�B!�"�tyTfb(膍ö�4����Xx��=n	�T{I�ƫR�!]�
E���T���T��C��W�z�:�«Xv�_￷�w:��O�Gn�T`�6}�rҒ�(��{2��p�K_Ã�0�Lݗ���*�@�%(@Cǃ4?]VB;�0�a��{I��Ӛ�R���������I�ř�[i���b|�G��[���Ji���i�H�����ɚ�h]{k��G��մ��g��אfA�EKm��l\��f���fn8��9��[�Ԕ�B��>��3�f�(˱?��sSk��ԍ0����r�)Y��1x�$@mb0��dlx��	���Ӹ=T�uƣ�����{��w|�Cg�J�K�+'��/����G�~J��ub���BNC��&2��l6��Tۘ|7k}���b�G5�@SS���X�T�����Xr�{�L`۫2ᝁd��c�Z�����V/���Q<5�;IK���0D٣z�8��^�&��<�ӡj�}�1���O����u����?������G�/��L0[��َ�\KoeA^9;ybW0��a�?���g=�Kר�?��嶜|�V�&��bZ3��}B4%���뵊�����zpr�&��#X�g#��fm-z�`ײַSl�PX`��)�M���k��(@FH!�+��ubDWP�2�R�����v�Ԣ�h�N��=0a˶��ܹ�Q\�kB|�D���A��y��e�vT���� ����:ʘ�!�*�����dc8�|��7�2	�6y�-���u��׼�%�ٟy�[k5�͔�<3z�����U��O!��)4�i��:�YШ�9�ג�g��Y��,��gȰa}����hC?�!�:�&)��z}ʺ��ﬦ_:���������%ݎzI�˪��[�W��`U&a��,me3��j���y1�O솢f�Z?�앨�P)�)	0���Ѯ���������_U�����?P���vs�R{ǴWw��ܹS��>tn�9�}���z�W��&n����޶?lv�KN�,Xܚ���hz�#7�!��#�|�_ 1�*�>�U�O'+;��I������&�q��)��12����q�0�9��;�$���X��;��~������9b�ښ�'[�sL�2�I5�	�2��G ��\w��������SE���&�y���↓�Fə����w:�u�`�1��#�9.l��,8�q)�$�b�Ϥ��,�4��󻇟ܙi;�Ӄ�u���0�SjTv�����T9`ڦ�InF���I5n�Z����Q����u���/���gL��*���?W/�<���L�;�H5(��k�����V`t�1����B�W^���u�����X�Ϝ�W��DD���z&q���D(�+�:w�S{]�x��{���<r%,�۪�������ؙp/�:'�=��3o������aU�ʗ�&�~>V�ǉ��\`aHk������ӌ���{�M�@G.�/j^��p_ᵑ� ���(��ڧX��@֭�O�Ց*8�O�:��rN����'2ӆHSZ�O�Z���Ϛ�+a��ĂXt\��x9�B��W�D�N��0F��l������N��Թq�S��JB�P?���2�P�d�{4�Z�-�`g�9�(�s�]bz
d;�8�������j���3�����m8%�ez�^�.΍X�p���r��9��Hմ�8ok��]3@��fw6�̼L�SL�5&7�e9�O����3�x���X]_*�K)ʸR�X8t7LSW`˥p��R
�� �Bk�RL�@�G�-��J�����������ᷮ|��ߜ���W�C-���σ���O�����6w�������~�8Zeu(�ue̾Dfa�N�$���C��־��n@�(&j��S^y�'k��b[�"� h�?gG	
Л��|�#���e����V�� b/n��V��A�Q���$�@�Թ��_��<�كh] ��D�iÂ���n �(&z��[����φ�4��Z��`�'�~R�A���׈,�`E�փ�!�:ڌ�hE>�+ޅi���<�z��# Sm"#�5�������y0�X������9	���8�a��Sq0�5"(ϻ�g�ڲi}���c��Z��Κ���3Y�	=�����6\���<�I�����b��{A��\QFȮ�5�C@�z�EG��RgG�̈l��fq�'��3'�*0�7}� �	��ʃ@�7廰Җ�4`2N�=���[�^��>��{���>�Jq��������3����~y��5�h���"@I<�VC���A|� !9��\��xP	B�^t����P�LV��8n-���fT4h���C]I.*��y)gO����{Xݽx>���/�9AV}M#��d�ذ�����iŉ�ɩ�O�h�/���k�
�i4�`e�ďW��d|�c��:EA9�@]O�,V���$�'b�+�M��n�.�	���JXB7�<O��5`+���"�)7%U�lV���W��Kt�Q�M,����2*ȡT���8m�f2��N-3>�NC������������J�^ν�$��-xaʁa�"I�G������Y�4���������dier�d�#��U�q�V�D��W�ЊQ��萨5��o�i��X������cU�m�g��s��e��������n�W���lk�5�X
��
f2
���� N�!k$�<X�d0ʹ��=��Ǒ��u�u@��T��8��e��eq	2tT��ZU��l�ęq��YZI��^���M�����D�����VT飥���I�*�l�*��3�~�߼�p�U�7 }�fܮ�rKP(�Qɹ��&7jŞf &�?�4S
8�1V�qc�LMV�����ȚtC�V*��E�ɀ�V�$�.�r�٧�a�:���P���0z�N);�w����SPL���h�#5���}*eH�h�"��\�J�R��5�5���n0�]�X�>]�lw��o{	��M�7��'g8��,��(ܕq�k��^C�8�S��
��X�*����䆪5˴�"�8�}-;SˊSA�:�Y��x�=�п��'`�}�T���{2�7�Z��gn��7�3��ϟ��c�7e�Rt�o�H��E�����u�W�����ŝ��W	��`[M�R[�n.(�l�ױ��H�J�f��L������9�����u�W�A���X��(�H%��=.�!k���I���$q�<�������FY��_:t�J{;c�u7<��ZP}��<{|��=o.�4�O���}��}鉣p�G���νy����<��]�,<��1?��epMk����|/ƲO�fj��{��hF�VC�a�uDfL�Jt��̎O���oj&��3��<K�Z�;um�Pp?�+rhB!�~�����H0��j������r-�G�,y�������5��>�	m�GL�tJYRE2gl�mj��#��S&�B�e{�2�^��^1w36���V5��+�8������>���"��w�8���7��R�{Y{/4�'�����^v��je|>s̆���ס�<ד1E�J��y|�6�_�������o��>�������p?{[^����+�3��]�m�u��c_��x���O�������^|W�`��;j�o�Z�Ǻ���Z)Q�z�A�Y�oZ����V��et��f����\Vg����J�����)�HM��o�.rz=`��n��K���3����u�v"��u��~,�鸺�@�z�>�����\�s�,H����_7���?���?��W�������E��Q~�EQ��M1oG뼉�y�O��ڷY�k,�Z��͌p�n<&�/EU��C4'�i$���p�Z�<�x�fSΧ!H�b�V��l��Ԋ�d����"���6�ߴ0IDW��$On�G���Ic��^�`�u�8zb��ʗ����ڏά���݄Ƌ:�������:\F�8��P����a!_�.�WDi�T�{\�t����B�E3��X,�~|��$H�?��ON�+7��ֹ��������ಇ��l��k�:�0�������C��<3����1�ڛ���０꽿>{�?ߤn||)��]�ϺQt�̡�8e� �6���L� �;�ւޫ5ؓ�`��D-���F�%��Ϊ|�d�ĐRdw��Np�-ED�i�&�����f�ǥ/U��}��&���^qs�3uh�68m�_}���({�Tu��s�9��G?�/>~"­�$�
WA���P[*Jn�-G�I9���7�Xz�V��I6�U2#h��m#�B��Z��4������d��6%Չ_������|{S��N�)0|Z�ӱ��S
�+��,��4%T�MӁ��\7{ �t��6v���DS���LM|��w~���^����'�d�ܥKq�Zj�z���s��1��5��Zq��&�4���f�a(���5��X�q�(�d�"ʆ+i�j��5�W�����߯-�������+��3=4 ng0]�CG%0��I�֟�:r���˷*u�������Nt�\�超���U��E)�����}�$���X�xiC� �Sa�R���p��}���p�AI���!�����U� ��I��_�������,�����+�h�Iܖ�;����q�]ڎ��4mo�{G�c�f՟~�G�RsnG��k}O�iD.��Z����Rt����>/p�Z��t�<���d��(77�i߮�:qֹ~BD<k��<ם�%�#�Y[%O*��+�:!B�պH�����ɽ�甒�4��xm~Î�d�⣠
^+ԯ�������9ʓo�k�<��cz�*
ȳ�������w��� ���v����;�J�c��;t����*I�6	�(�Q�Pq=�լ���K��%�ɕ2���V��i�GFьRΰ��5`�M���l�K���IX����m����<ڽz���Ci:��G6�7���a��E�������~�D��9�yI�����Zvx����rt��_���"L��� �3����B�f��{�y�aE'�=���(DW?�D��=�^�Z/I��&n5x
��VMa��Jh~��Cd(4�`1�v%qk��-�t��.x��Я�6L4c9�S�$Q��o]���'7�����c&M�ێ09��K��(�</�C$͛��;6��H� )!x�'��\���^��5�c����C���f�P��g8�O�3v.9GW��c'�ᅐ�c�Ej��{B��F�5h���n]��b�'�A�Y挈����,k���F}o�+z��ߟ᝻�Rї�������v�3�'AR ��vq^$�=�0/[k���� $�:5����a�lxF)|�I�`-��CM���)[h[aZ����M�a�nb|W�p����l���-W����'���S�k�|YZN�M�5@�E�����+���s�i/�W:���,���iiE,H3��~���H��4����(��Hb~\�0�-W���$Y7���d�Ś���r�q�7�a�Q�
g�)�B�BV9)褓\�b��&���h��y3�:���	L֧��G��h����sb���pq�s"sr1��ć9=֘�9
��;�?j33Zg�fj�����$�\�U��w��tT��.�2v�\7$x��(���}wm�}\���v�Q�/I�!��1��L���?�f�iT�O�7!Oi^��C46�iS�o=Yo�T���l,n����ST��C�[	}�ٷ_w�c�c@�4��N>���m��O0�OaD���L@Y����d���n�^��wb#*䁿�'ʵ0.lE�u|��f��p�ʩHy��Q�7UӃY�Z�%UR�a)�*�wj�Z��w�rR�9��3:q��g�,cq��0�eQk��f�{Gs7�E
�־*�~c��Ϡ�d��^L��L�S���q�7���N�Db�l.�U�1��ؕ�
���������`E���e�0\�*�|Ki!���(�ZX��hS�\��:9�A}�I&�����v�I��zQ\cg�ɀ��\���o��zr̈́�����y`�Qi�IOtƓ���JX�����;z2f�p�K����z��}٧�\q���7W�z[�'C
��@�B�w�0����o�<Ŧ�MB�0�q�
9����E�l�l,Y&�@#55KG�MЬi9��ɢ�4X����w��$��Z栊�P��֙0�!y�ݺ�}���r?pÓ��r�:Դ2H�<��7V8�h�ʳ�^�6޻�`GΖ��RD[��5V�����]_���I�������}'�jA���^P�xr����'��܍�W��'�r�3�:q�'���9]G�\}���F,���%��z*t�b�h3?�RbA=��}8�M��v*���S���$]�-!Z�V���s#�v;Xq�7��Q�d�VޓL��Yp�>Q�Q���"�e�! 6'�XA�o� /a<m�zl��wS�L�Z-xldݓ,�7����U���W���]Ϙ��&mh<פIvn �
^�$P����Y�z�V��Y��[X��j�n�&iMEm�1'㨺S8���Vc:P I����$8KD<�����ep`뭀EO��W�}������u��O5~�]N8
��|��U��$˵(AE�.�0IS�c�`��9�6.�̺>f�(J��dWۨxvR���"FmF܃b�p=7���|��u��P��7���0�5��P�R�!�M��'#���m��v*��t(�*k>��n���?ԋ���m�\��ݩp�~k���z�˔�
�^�)%�gCػ����Q�}k���3�z�<���ӾVΌ��X?ەQ�\G�Oۍ�(�a���f�a:4oa�]���g�Wna��T�p7�i��������[m���cjAð@��?E(tB���ģ���x��l��Ǩ��fQ;������1ގK����􃂤-�����\�G�
y�������տ}�W������Ȓ�¾�麒�¤�yT�Մ=�:Ml�����+�;	�v�t��&Kum��L@1�lAǧf6�j���IfB�:�f=��9h�v�0w��]7� R ��+Sf0%X)�jc������.PE\�E�
�X��	�0���M�ip��q�d����.8S
RQX.�<:Q���[���>9����_���޷��<�U�ʖ��ɞ��L������!Vi�z����x���@N��.F�!U�^�ZWR�7^�1�>!�{�BX��n�ڼJ��_|���>�L֧FB��GI:!�,W��y��(.�J�)YqA)�O��G���\�֪��9w�����˗�|�� �N�Y_��#[�$�L���i0�e'��UkC��ɭ'Y��;	�ɠ#�jj���~�a��澥�*�:���=/\��*�}��!ù{P�b���}��G*BZ�斳�j���-���'s��C��i���0��]����wk����Lܣ��A��������毪U&�I3=&��C_3֠o�B%�n�:Y��5��f'���b�F0�9&b��wO:��{Lo>:C�N�*��YL����o��Ȟ ���ز���E�0%��D���K-x�\:zfZ̈́���@�F>]C��1�޾{���;�A��V�>��ʕK�se&�,-��pn�,W���m�/�gZ���Æ��!�X��Ұ�bt+Ld��
b,�0~�����r����=�yD�y��_���_���3��1}�ܫ��ҭ�C�p!���"��H�����z� }3�q�<ulsu�B^�	�=T��MH����P�~��7�����8S�ȥ�.�1����������dP}x�gh{U��g+8�.�B3�����7���R����c*[ɪS��g?�����5�7���W�~E7R."hh6�pd��\*�K��3�Hn�<�	����)������lx�J�����-�P��hJ�]�Xt[��Yo�Z�ƹ�\�a:�?���s�7�h�ֹ��w�I�\�-~3����N��4҂�^�Մ��	��]�z��P9r�Rξ����Ƶ���_A�ƭ�舅To�>J�Q�Q�v#�?ki��֭5p�����Tp]�{����Ӻ�����p�@�Tn�|�`�Q�=�kEj[-E��m$��:������U��l�����s۽�fj�K�U�o�������2]�gKmV�|Q0�n��ya�J`��Ǹ�b0ny<��3�s��	�dc��(5�����-z2mܭd;��\���n��z���dW]�ܿw�}�o���<��ęW�Ի�^��R�����<_�ǫ�1�U"@K�r��d7ku�yHovAR�E^�Hh�B�G���������Nc�L+s��u��A��T���+��Z�I0��]�����.�=���[P=��<�rE��ޘ�
Ț[]r�n;/8�����0���/lu�����������fX��Fέ�T�I�����w<�#���h��|Gb3s�V�xs �@���]0]y��BM:�m$��.���eB���Wv���z34���W��U�����#\��2��F��<ޒ>}/��Y�fn�嫼�ܵē_��ͮ��RQ}V��;�A��v�C��r�������gU�	�D�6�4'>x�^xJ폒�C^}=ҕ�c��?���3vf�7�On�{�7~z������L�����]ԼD�l)t��w��tny�v=��-��_���o��᫓�A
t���{TeAD�~?׿���I�r<�!.A�H5�X�1Z�:�`�0+��D��?�^o�g>���ﳷ�ySݺ��#����?���<9{��8�%����V�:��)���ss��,�Gx��d�w���.!�����x5�;#���������xٍ�m�I���ձ*Lr������}Z�:�#�P5��rG�j�'YRX�_0c�m �_Y>�����E�"�U��ƹWI����ո�7�@y_����d�+	�Q���v/���1�L9��h�4_!�N��YZ(���|��(%��l}wq6�/7�0=��zcՏ��(�#fj�j��?�z�Y[�7~����{�z�zƚZ+���<q�J�_��NzA-H�V~���78���l{�Z<��r����fGl�'R��e\'�S(������P��rx_W�ň�n��&"�76��lC	��J�~����D��Z�,�����sm����Q0��Qw��D��3����Vs���m2f\\�PO�o��{����.�����v��8������8q��X)z��8��4߇۩�cW\F���8o��&��^)#�O����1+�Ђ$�//Խ�������O6��u߄=�Z��B�L�'nݳ��y!��;w����l�󮑰��}���/�VVR?Ͱ�&�n�eT�+��DŁ�\m�M0^C<�肉%pL����s���;�N��OEE�{n˜z����}�@\q�A�W�	'�`�3r���gP��ib���(�
���C��d�R�|����G��Ӽ���I�^���s�Vvr,zl�4Dg�sFe+��V�M�����Z��&fȖ
�_n�wƢ*P�#��b�����v�Ǡ��,�^:V᝙��\8�oϫԺ�~�؇�����������������yWI~��O��>��ZoZ��٭8sМJ	��$�� �i�½����Y��n�gz��>v#&T:�j�5�8���q���q8E����sn#��A��j��\�/� ǵ�Q���bi��e������y�T�mWN�o� �Q��=^��r�Q���c����A>�>Fr�Ø�Ƨ��'�Q��ܰI&�u[�tPWQ?Y^A�"W]��(�=�:9t?�pU�j%�?=v|�c�y�W���ˎ��_��޽��g<}��ҽ+v��g�|ڔL�)Օf�`yJ�^m��N��k���1CA+���q���$><�@��s[�MR--.�Gn�d�
�ÂEV" >�14�i��?�n��E��D�mv.���� ׅ<A>b8�L�����<U��	�B$�r�#jTX[fZ�w,��zPP96���֎�8�ĵq�Z٠ؾw�b��.^ �&��QfN��Q_��	8��dۂ���G���6/�ҽ�s߹�-Xy�����x�J�ǐ����4o0ǭ�V��K9{];�ˣj)��A�P�(GA��ˡeXJ�q}07%T}�$<��6��7ެ~������J��vKw2�8lD*mQk���e�ѤC��9==7�ٕ��UWT^v%<� \�F�����c�����:���=ߥ��,ޝzm���Ǜ�$�a�G�^A�Z�k���߇d��k�T��!k�I���u�}�*լ�!Uh�\b� gѡ'k���k��.J���f�����?x�.��D���&Rf~��W,[I*�ϼo����>��Y7]yf:��"󣧳,q�Ж��d�S!�=�)��a30�������/{��JM�bϋ�'�X���me���*�{�/	Y^J�Cឣp��uXZ�4��z�h�pQ����n��ԪQ�{��ZiT�貄F��v��;ƥ�z���0ZZ��@���c����/�%��|C� Q��7�u��'�l��bH��^��%�|;XV'5�B7W����ѥ��	��V'ySXq�Ћ�&�rLj=��u�k�>ю=|�~��i���)�G-^/ެ�`
���g�';a�|�����ӛw�M=��L����I�Z��ŵ�� �H'� ���$ve���m7�� 1O�
D.��e�vg���� {��D~�B~5OT$����l��s�أr~~���r׊N;ћ�k*I�%28�^�p|9#a��|@í�f���&+B4�4,�F�/���q���T0��\�r0��{Dw ��L�/!���͟���Y���/��._�s�E���ܵe���6�V<��I�mI�٨:��4Je�Q�02YY��.H�6�LD�値:��ı�������e�c���)�����c��,�su�׋���+�}��L{Z4f��j0at�&�_�����)jY�m�՚	Դ�2U�t��C�]{]vVz�pl)��3c���k���]g��~�0����hq����iP&%U�6�Ʊ��$�qB/�Q�L1(��i��A��̥��Sށ�}]-���O$�fe�Gj�'��8Rq�{=�(\�U�Pc���,����Z������޿�r�/�:�\�c�Qez��*�;�{��a����O>�A_�����^�x`�=���K47}��V�t"d�R�BuK2G�K��"�ß�Z�В;Mb%�̵� �V*|!�@��L�_H��0��E\r�����\�R�-�%9�wk-�^V8�n���D�����o��8
�4V�D�>D#l|W�� }*o��NP4ky�eX0��'�jM^�5&�s_zr��S�DC3�t|'@�딉.b\ E��pL���i
<��,%S'�u�{Da���ic�tR>�N1�m�=��=59�^��Տ�<��N�lH�5��+aqk�@p�9VX�M1ʔ*��E���Ot�s�\�Q���a�9�TE!���2���|W���k�����W��aq�I� ?nT�F��9ԡ��'�*����pݙ��7��Eo������I�ꑤ�J$ԉ�E�g��7�܎��i%�G:�D��k���G'�����O#lP0����Q_��?*)�W�h��B@k�N93�[���{��C>�A��+�(�8B��j&�V!	��Z�6i2}�����Jl�׏�31tf�U�p��U��(��_�N|��R�&X���wQ}��n)}��f1xu�!�J 
kɌԕVA_����5�C����@l�l�2s	�+��'77�(f��Ѓ��	y2�'lY`�j_
��6?~#�t L�E��f���S���3�?��.z�]���~q�`R�`��(ݙ�{�*��(.��>̔�S�7
sSCJ�?d�	kP�o	8��\;��6Nr�$N{E�Pf�0R��P�pJi�1�if4}�4ﰄ�jV��H�c���FJK�/�C�������V
�2J8{U�2C)�Yh��p��� Đ��Fc��Fʍ6>��FJ�Mr(h���Y϶d&��v)+5�^�YGXh;K��OA�^L��R[`�"����P��&�
)��5�g7ܾoat��������Z�?��l�@I'炳S�A*�)�ʙۘx�[;Łt�I-�֏�A;=�������0S6S��v;AYTq��t}d�f��X��̊Nk]p-	GG�Ղ�|�6��v3����s���L�"�a�`2���E���5��ױ�����fpr�,�k�~�`4s@v�B�^�gDqS�&�`�O�7��g}g ��%��f|�]�D�2�m\8*���9Z3���L	ʰ�&C8
5����V� ����:/�6!_�ܕ���)V��&����ќ�V�0��`�D�2�~���eV�
��r-59=G�۸ܺ`�4K�c��bE�\�F��"������N���޹���Ǉ����cF�f޶�(�e��fi�3!#���bl(F�G.x��J<�x������5�t#��q_�Ǐ��$h��`���6�h�k�F�C��X$��y�r�&s��PX���T	�itۤ8xR+�a̘�C'���Ǹ;w���B:],����X�	�c�+���%�������{	����f��J���B�dFh&���q3�# 6Bɋ�β�ԏ�<���:�3Hq�N�_8���CuxnW,LC14��m�D����db�	�ݫ@N{}n�4����?Y?Kx�.���Q���:��jT�U�.��+tP��,˳uǄ�J�L ��/ZE���^Xh4��U.��!��wH�%�8_R����itR�j�Ib�#�l��V����c�������4r��ٹ��c6r+w-灱Y����:���5�N�
5#P��`qq��~�b���cu2�������ZB�Ht�-�����\$�D�����)j���q�����C�c�pQ�B�]M@�V#x��1�NK���P)2
3}rw͉8r���+i��j�F���S��e6��5����(UhS%[h^����5^�D�P�eztm3�g_P��%n�eM�ߋH�w� |�{4���#c�2^9c�%���#��WC�$0Ug̯�p���a�ōXP	��(�*0k��2�l7�
g���,Bg�'�P�Ex�^�/rJ���"{���E��Eu�ЌC�܂�l���m�������[��_�a�0��8�K���`�:ɚ��V��̐F��&B.�����8E�(_��uprZ�(l�
(��y���2��f�؈��u�z �\O����*~f\4#O�,/���j��2) �r�Ox����$1^��މaD���^�d��1�Òxa�aq�<�,64Р�ED�_�Y-'�X� ����'�۰0��Rք6� ����i��jHQ@����]TX+[��(��A��Jh�(��	bή݈cn�U
Ņg�!²��4��1.�V;U�k�˼)�5���������x���S���q��X�~=ԉ.e�۔}�d|ƎpKɊQ}b<��`&��YI$���WɌ��5��kT٠ [�x(r
�o�%�3d�Iș�k=b,�z��d��q��ߥ�F���:9�f�ta����������o�HB[X-_i���hpS��,�P��}Dh�p�ͧ�k�)�h�jO)���h�?73�^��G"�y��4�i���Z��0Ho�s��&�a^F7�͘R���
���R�1�J����]v���v�b�� �_��5k��C��9
�!�8z"�]ţ08}���2h�Qmd%��$]��Wh
K�3a8>h�I����)*H����f��c�0��;땩+��bGȥ���OO�򁍮��7� 6B G)�La� �L�^�-*��%��&T���Z`a�.(t�T2������ȁL�n��(v}&��MHr�{�F�7�F���G��ƃ_R6��G��y_5V�uB���u���/���c���Ɨ�!�Pf��UJts�0�<���;M�9C��M�����`'��0�;&y�BC3�`���`� ���B��|�}��`�'C�������ǭ*Ō,��
C]��+�����+ث���8�]��o'v!cze�}��Ӡ6�߸I��\��3��h����44_1P]qW*�NԴ;+61sS�j��C_\��Q����&�	��[,�0����qq2$%Ja�V1�VA�B2�B+���"W�)�f�)"QF��Hi���1�]����a�o��_%hJy�G�I�NЌ�����s�� ��]����#�Y��NqbbM)T��ꑇ����D0
a�^h#X���;YKd<�Γ���$S}�ص�O��V?R��Jڶdo��V߿7��u:{�ae{����܅	�
N����ٻ1��Np���q���SO
fh~���O�r�����Go����BE E	Uz���$�h�9��9��	���&d�Z1o����d�}��9��f��6���
�]tς��։(��`�Pu]hR2��HD�j(�b-�ur�Q­'�m�&I���i�0��������*���s2�x;"��^�;���K8$*���B���`�'����{�%�C�^������z���כ�SH��h!��1Lb�:d�j�����,K]w<ѽ)Q4k��fP�|�$��+��-�����q��8�^�mP�s�%m���]a��G��$�Кz��4&2@?��T��[�u�rYi�g�����`4h�8�סSr6(�XzJ����� ��L�X��	|Z]F71�Wc����\�2�S%q��(ܙ��s'}��~��prH�v����0V�wj4SX���m��npLI�۝cȋb.���iv�\�V�k�o��<���X���]�p���Z
�"�0��!��?�!�v���H�,� �`�w��R���@�OSa�b��B-ܼR�����X���1�c�}�`�����Ƿ��VN�a��/a���M�2��{@%��|�+uu#IZQV<?ZM��X7;����˵ʐ�L��K�����Q ���/E7�a�*���l�*J[D���q�Q�����*��𫰖���~Ͱ�����aԷ6ר)���87�Q�QH����������m��oV�$f���N�"�j��N����*���<KPaW�$eBkd�;�+���>i3	�r)�(��i���p�BiѬ�T�S��HOf��c�o�5�J�V�ҫM��������_l6��ŌQ�C��
Z��ZXc��y�*7a^6��ݷlq ���$u�YαD�2B�K;���&��;���i	(&���^o6Dh�7�{�{.�_GC�h9����h<�ck[�Do�� !��D< � �n�ޑY2����r�m�L�T%q�U� lx�S[O�G�-?��+*�vA0S��[%e%H�U��3i�ނ[����JYk��G��V@�ՇN�5
�����ds��ۆB2�S&�;�7/�t��T
-d�ēyZreq�E0�OC�,�f�U�X#5&M����A� �ۈ���Y��s�[|��@���+szUH E�;`�l��ǟ�+� ����4���'X۽��Ud'W�G$���HZ*,�{�'Q����f������K�,M&R獿����O<�J⎨�j.N#���Pi�N�8�>�!f�!z���ͫ�vn%r�1I%�9"|빂{�Č�Ҁ�/j?���K���~�|��~���i�ję�����%�z���/����av���T��n�D�N�E1�Z䘼
����$���$�ঈQ/�]����<��z�r@Д�sJfey#�Ÿ��{�}����E���}$ux)��ӌ�n�3\P�L��UCu
���D�\9L{t3�d��!g�5m5xya��Tk��$�	i̼bo`f$QY��l����<jf��Ɂ�,���08 �P��}A>>�ʔ�����q�)���oL�����w�x����+�t�EW��wb�1\�����|s�8�1tSIG�hEUŎHT�ˌ�/�y%�,�s0���Y�l���"!^�4�2� V��+�Ŋ6�׆��,5��?n�������lt��!�b�8̑��D.�	�s�yZ�D���҆�j'�9ց�%�iSŝ��`%�p��4mW����чf���^mvYF�l慬�9�K�j5���O��!z�Ņ��5[��j���K��!�T/�vT+��"Zt�)H�uCb�)�+�<kr"vm��
�2c$�zUH�F3VK�,;~�}wE�'�+��WD���P/d*ٚN���q�|TI�"��h��	�|eF�$-�Ȝ��X�~ٓ�xmي�j�I\0|����b3�A���C!���
��C9�	Gq�c�[�{�z��N�Ͳ��?�Q���#�Ja�v����2���.PM�w���D�P�V<��<��
*c�hM����Ke���Ŀ�6ә����X��x�_�_OL(0�Wq���JZ~/z���Q�L*)IF��!��p>S,^K���\�͏/˒N&�S~���Ź�J�R!j��E����Ó>o9[���՗5���b��6q��C&g�:�`�q0OozI9�0���m<Y>_�M�������?��z����$��L���*�A�B�W'Z�-��m����j��s
y'��ɥ�Ƿ��_��|�ܱ%8��U�K3�!���:dI�Qa4X�͢\k��'�%sl\-:��ȔѢ��"/=�Dɞ�o�=��%��\��Zl�����a�j�,��ð��F���P��	����Vk�_���l�O~z�̓:�'�l�$�D6��ڻ���X��L<S������\/DՋ�P��\WfRb�R�UϜ��串0AZ(6��R�Bq|�I[j�4�������(}�7���yQޛ�"�5��#��a�f��T��}�����关�V�2������K����^x�{����C�E,XVA�>9��IR�*�ʬE��e"��� ���&�`������PJ�1_83�����U�b�����d�}ֻN�y�<�8^DȬW?�����s55��+�Ç��r��ݓiOA1���L��\��,=+K�{O���α�%���3��F�jtV�g�O��rO,ĥ���J�QMm�~�D�u�dx�,�uZ�1[���[�=/zpS}/YcJ����Y��׾������vw��.����z��1�h��q��4~䛶�����4kć��;���ŕ�/9�����/�t���+&XB8'������.���g9a�Y��L5�i ��	�W��q�"
�C�F��`h��	��R�s��[�;'�jY,%�l!��l�c�بU��EG�!_�V޲����>�����a|�:�f��'v�'�m]�?����t��+op8LyH-`&���s��dڣA���s�����Z1��7�����-�h��$����ݬ��a�c�k�����������n&�<9�F�>�t����}o�//-/>Gk�U��Z�H���Y>�S���\f���~�ox�Y啰�!d���Z������u8�<��V�b���-Z5���|�W"J̬:��J9���%�� 8,[c����8��s���L:It�y�i�>x���h��5XZEG���"���(zU3��<����o�s[���غͫL�\���v���*r���8hH��3p�	묓χ�%�6m�+�����R�������M�m;�:ѯj�{8�cn�KF�` A@@�&@@��T��F���sx�_ԟ-<�)<@p@�A�	*2xA0�l�@�D�{s���XU����Z{�}���E���u��k��U����K3�}w���1 V��zq���w�����`�۬߼��Yn��r��Ӳ����l�0�v�mu`�N����Z�"T����G����>y��;][|d!�3�^V��~J��5g�6W�J+�+�Sx�v��&��]t�����l��b�[G��9�.��ۘv�e\߿���1^|FL��|m���6n4Ҋ�PJ�Y��B�&�9T�"Z���'E�����{���t��v����l���T��g?z���#�Y�Yx~�ѻ��Z�߬��'��{��^>��/��&��Y���La[�h��	]�B3ơ��_��
��Ic��fb�L#WK�=B�� #\e]"'�+QQښ��e�~%�.l���i���/];{���N�*�j�wI�!��x��_�Ǐ=��%W��?�v_�)��5��Lv�B>�L5D�]Ͱ30�%�/���(LQ���.��[�i�(����g[]_��1W`Џ��"kwW+�i'k'�g�r�����|����fQ�J*ƙ YL9�D�<
n+͞u�������3S���3��O�~.��[8��
�$��b)R[�;��eI�dB�u^�@!��	�|B��r���O{T�U�8�x����i.�\ڎ�b�9'cF�tqɧFD4�hh��ȓ%��di���Ҕ�u���0����_�����?�����r��<T��}��TU�1�Bt۾1���H����2�#e�sFC�4�D�:���G����"\����w}6��͓��TY��=�q��sζ(�+�7�2*!V�pAF�i3y��"!�ܹ�Ӫ=��˲�^\L�]g�P	����kl��ʄO��ޖv�Z��t�A�@�ư�?���
{�T�r�_^z�w�K�+g���/_x��υ^k��T�T�b�'���kC���ڧ�?9�+J�)��sl�ĭVR�	�����!�%a�JS<��"e�q��x���l�*�C� �Nr3i�<e��b(>+�R�y
��j�&���as���҄">ux^��p����+z�j���rZ�i�m%��읹�U���T�{��%RSع�^*�+�ً��G�e�y��������w���;{�����ǽz�	�N
m&s�h��%�ޔ�m9dfs]�h;������㍝Ʃ�3<#�Q��h
�[�Yr���y��]�G ���G)L�� ����3���8�K�ΥT�&���E
5��\!��b��2t�S�6��q\陸�|Gw��/�O�s�w���㿴�w
^�H�M-��]��Zx�V3&�+��'��CO���'.}�͟��W������P�P��:�)�1��J�jڴ'U����ʗ��"���I��\�7+�^�� hc)q��|�2�����ڪ�=4�O�U��!�G~�L��1F�Ŧ�2�]+ȣ�tȦzs�ME��Eh;��J�����T�ݻ޹~1J���*��]1[u��+�em4�W!��i�9�->۵����=pS�L�*ry<���|�UGO>��N��������<�Ԝ���SQ�5K��\�|��^7|/:f����5�\/�5��|��O6����`IO���{�[�m������kfd�i��q/y��������:�O��%�X2|a{���dw�$�Ė���5�X����Ie�d��3W�}2X=�����~7Da��,�5�6e��+l�����}�r{�=2�����=���]�=�^�����QD=Gky?�7;>=t��x��a�1�`��}ᓟv�������y�+��ҏ@֟���d���W�f-�DG�����Ϻ����k~�ƹC�~%\����yG?�ڮ�YAlS�`�'�2H/�"���P�l�T�L�ܶ����B�l"�СH�2`��*��/-�H�-i���T6����U�c\u� ��¤�1��5�#R�)i�t��iۄe[=W����bmL��:ʲ��R�����tN,N�a&�=���dey=�,����k���ޫ:K�µ��a�0b�7�cp��2��_z�G?q�$|�����z�K��#ߡ��g+׬�Y$��|7�o[��\��� ��}��^�p{�g�����~|��!�j�w)�v0�u����MV .=�RJ�#�Z/C��� �~왻o?��'����sw��E�
W�o����f]..,p��d��	R�5a,y(�F�1����m�xs��"��*B�<��K�+���J�O�[L�չF��O,�yqg�� 9�eOg/�Y~���wY�&�#-�w�m��7�P������C����z�A�>a�(��(��R�2����l�����蒸�z�K���L��%�O[���H�c�z�Ep	C�G�Aj��v'�P��R���i�25J�_��f*�8=�/s՘�N(�$�ѵ���h�	��$1����k5��7���D�`-ɑl����@GR�m�����W[�A_��p�)�S��qQ{J��7���0���y�ŧ��U���[揟��dy����#��-w��,��.�,B�Q�K��rp���&�W�t���2������7q����>�˳�w�*EI��!gR��~I�O�y9���Ga	�y�1f 2Ҍ�(T2#ܻ��}Of���+�ж=0.g�ձ�~Y?:�m->����{�g�/�+�(�\�M6��߬�����+��G�!��7�Ο���;��ZM%I���͛�%"J�az��d��
ԋF3�L��,|� ˆ��\O.�W%g�/ί\���4)PT(���L��=f5��������S[\�'E.���A �ߢ���d�YՎ[�h���&�P���4��)<���ʕ���j���2�,���C8�3,][ӖY'�i$ʌ2� YE;��S���W>R{��	�cPx���y�bM�R�����\��f��%(����cD���㨨ߧ�ST�(�I[���5C�BB�P5	p�:n��k�)��γ���yډ�	Z�{���y�Z;�W?-�.ga��X�d2��VB�W,���Y:H����藱/�2���凬�ke��;uP�Q@���1���c�l �9�5�����}$	l%�>R��dQ0㳐'|VU�P�M�v�&�<j5����£�4ff���@|l�F�+�D��2��[�xS�sf&��D��Grh��"�D���^&���9��ɺ�Aq��dZ�Q�miӈ���/x�����pT�j�f�YSv~����S��1�Iru~�b~GSI�5'��4h�%�!�>���#���l=�g��>cmq�ɍ�����P��#S&�2���(6^�$1��lx�6y����w�E��xO�R����� ��Ā~T�&|��$ΜH)W��r��	��H�pV��)�4fmK�i;bzb�''�=q���s�>ng+�/L8� ��NTq�������u��
��Ҷ'/��uO��(��iOH��*o���[�"֊��Mw��n��	O�felpUhQ�\t�������@(qH	��CG0�OQI�6ٙ3��)$��F�j2\=c��o���I�4�l`2���-��6��421HB���$2���ڲ�_o���Һ�����+b�M���j0�b�*C�y�m����\��v[g�<�	�tG)��HuʃFM(��T��ybF�a^f!RTgmt�}#�U����ɛ�Bp�2������s3����9���k��Hr��(펆��a����٠7��l#
����%��s1S�rA��#����fO�j��wS���Κj[ۮ}_m�Zv�*��O�2���b��q�DsbG7��2���9���ϵ MⲘƠ8�]:~�V����W�pvwd��+����>゗�FȑD�(�to��sQ�MQlJS	A��,���c��4�2	�:��� I�b���Y��7f��W��h��թm�������/�ķk�c� Y�ة�ù$�KiF�����~hʡp�<��<�A�뫀���!i���/!N"�d��4�?/�E�����6� ���<��i8�lOm�G�uԘs 6(h�J�#�U�`����'ay/Z�Q��j����\��ܼi����.�7���Yl�����rS-���DkPL���zYn}`�4T�p��b���
.X}L&����򈘚"2�L��#�N��D���kt�P3 ����P. Z���h"�qR�	���|����+U�*(��/=Mӊ�������κU�A�OD��.@��^>��F�&�r�.h��aj��-.�&��Y����9�����=.ϥ8#��_h�zI��N���1f:����4z&i��V��y�ʠ�����b��=��h�%,���.�����C��l�.�՗;h��h�9�R����y�
ށ�� �*Lhon��E�䨱�o��ep_S@�Ti�ݰO��C�n���w�
�R��&?e����23/z�"�-9�|��̅b�w:��z[	ޗpn��2'IR�޸�������x�v���L5,U���Ht� 6�I�r��g����ᐋ��N�,�\3$���E�P}Ʉ�S�X^�|�N^�1lb(�@�\��4DR�W��E��Ѝ��(%�eI�_^�����&6��3���'o�Sb�ށ�%�;-]3S1�����5k熰��f�M����yp�)�8�����h1?�k���`L�ʖ��?̝a�M;�T��!1xf#'�zN�몯fp�&��}_F�g��������aPP�!T���H�[���_� YX��+k�t�ч����&�[�'蔁"�`��[Ǟm4zH�>f�f[-`��[����<e0F�h"G�+aLy/Z��@�ұ3y�X!$H�s�J��%��k㌣���S��2*��9��ȉ��<BX}	��5�كr�2�J_�9�#��=J�0,�W[�A�A�X��]�{Ax�L�+�o]���'oc��4��f���hv��@	����[��z��B�F��.�3�p��]+���%�Q2G�;F:�nԜȳ}���3�M4�\�!*l_CEW\�h�1?I�\���w�3��i�d�F㎶x��[_��Y,"�Kx^q�$��W�kR�*��m��=���~�0�ȳV����gUm�D���912����T��l��TQ�����.5z�|3�����J�r"?ԍы�FU|]�R�*��Z(�y�G׬�?���.�m������3J`��w��������|���}����6�/��h�� 3�{EhS�V[�(W9�y0����d��H�ҙvlw�l-A�5�k���3��JՋ�9�/��ţ��%��<��`Z�Y�j�͏��B)��;.��*���5/�6�l;ά-��F(-������7�2�䐔9��-,�{\΍n�����ͼPŹ�M���;>�۶-�I7��GO�եT�?%�*Ƞd�����ʢ�C��c�<6�G�����E�5�ذf�Vz�m($}�v`p���ӇV[a,�a��Ԉ%�J��D�GGU� F�9�Z�u���FUį~<j�z����p��u���(�`^�J�� U>�<<�bE96�v̭
s|u�K�S�˭
��F��K���o�~�ߏ6U��T��Ԇ�(+Ε��!ݫ�����PU�!�Qh׶q;������Nn^�c�gΔPV�)���EI�[lk������� `������|����k�V��fD���0H�:y��3���&M�*"tٙ��g����|��e��ѣ���>�c�����g\+B�
SW�(Y�Ύ!`�UqN��z������61a쪝C�oA�Md���8;G�
�H6�WH�U&8�h]��т�\�����7�;�{-]ZX�Y%2k�fo�$s��a~G?H��:@�/25K�_iE�@��FlZ*�[���_AAm�e5KU�n�b�#���wQ��r���?f�Ä�J��y��h���丙z�^>8������g��V��7n�}�2�A_��ɣ�bm<jF[%)���@A�?����<dj�ɩ�fz9��S��X^!���g0��];hI~��8�G�)�mR�U�@�:��=�~z�嵴9S�/�Z��y��b�`B�LEui<Օ��[΄ۮQ��PD�����*�6h�]���I�א�7t_d�K�v0	Vz�Ȇ�b���o�OMnE�}�رG[�S�r�͞������xdW����?���Q�3R���<f-�u�����z#[9��&�%��=����JT�Di["_T�8�g���T!�&���oA%Կ��IcS*V:����B2͙]A�����X�[=�@l����Qqc\'��k��m��xj�Jٸ�ܼ��  ]T�b��lQ:��5-�Hie
�c)�7�|e�y*�@A�G�F��Lb_ w"i�Uf�.!�Q�K����F�����7'қ����񗕋�[�F��Ӟ�nl&.�`H|Pj��$���&!�� #T��[��]��f=U�Yw�}"q�`/�4V�I
�W�V0�Ơt�����#��u;:��'�4�ʀ'1���4�c��7�B8<wP�j(�-`<���\λܶ�&�pe��y��I1�Xu�}�������7���ɺ�&���E3Q����چ� �OM�l��ڪ�t�ɘ��"������W����GF�pP[s!��L����Q�;���,�#<;JXB��G�̲�٣��S;�,;jB�ņ7W�^m5�8X�si˘�����.^�'�S��O���y�%�J��h��d;V�jb��W��swIW��aњ������L�=�+J�c&��������x�c��h)e�ZЏ�]i�4�Z���(F~�@%��}�{����:�y�"��V�׮HZKW�Is*�r�����rU(}��-�B�g�<��O.������G@s2W`-il�f�����LR�UM�0�T�� �G�� �Z�(-[�p:5�XGl�R(��Y��8���W8��+�T������#�4ڌ�߉�T:&�|+LgB��~W�,ȋC�S/B����R�Y�]8Z�}mʵo�s��]����G
e�K9KAP2�ejjX��X��B�,kþ�*�Z�1�:���_�Mӑ�^=I���xln=��%O�q����,�!Ѳ��lf��*Ϩy�%�����%�l����@1_�n�E8t���~z�k<t���i�r����n��,5�61�&s;Ͱ�������_C,����]k��m1͵�U]�S����෤{�����e�	\�W�\�����e�-�%e@/��'׸w�����̜8�7���מa���ǚ
��7>t��{���y��0�v��/��?s5�A�K.W�~��W��M7�V�+�e˛K|;]�������Խ�a��|���S��y��o��3���C��:Rn?֜��d�ܫ\���(vD�vc�>���Q=�T-9�+7S4ѕ�I�o�~m���8�ė�=�x,�rd�>2��{�[���X7��Tlj��D9��;�V���� �)W����Dd#ʈ�sY!$J�c�]�Kӣ}\�������p�5I�"+)���`E���)L�x�s:�V��q���9ϻ�X]đ�U�)��:LE�/haN�f�n��WU,>�u;����i����|��wP�Ztj�Ne��/��Z��8evB�q�ȗ���e:�z��׶^񊸸�9T�n}ޥ�^�*��[�J���L�!��zl#���#AН�c!Iv�RQ�,��~����	UG�*C����Ycl5�M�l�3N��4��}���k�(��F�$Wϓ�?yz�J�O���R-�4�%�ӕ=)m�ۀU�"!���'��4[Y��gf]�{�ķk�O£ݙ�b�6�G�z9�lAPTG�5f�,]�
	�L]���*[U�{7�H5�t:
��]���=���U�jӵ"KKD�m(���w���. �y,�5.zEp%�Yv��ǎ��r�:�ˢ4^]h�����_6�ǋ���~䎟�����9P]��4̿,
��^�4|��q��?u�_��&�/@��Ci��4p{~�O�b"D��Ե�[̓�H�G���O����OeVa�U0���Y��"(����)�A����`��H�S�����r+�qq��R��c}���ܨ��Ư8Չ�i+��*�F�F9�|.k��Y���E5�_ܘ��cj��!K]5	�ad�5S*�"- (']hUH�B�U��8��=�Q"]ݳ���T?,5�q����7ߧbù�1��/<3fV��+[LM�{�f��}뽕:�/�J8�����em�ؠ����
~P�G�$���f<Mcy�e�}���������˾�^$���Qz!	���]--�5	�x^9%�{��������)l�=dH\�2a�="���9r��"�� a/�q���������3"If����ĵ&�Cr�*Jۖ�@m�v>���;�/M]z�c&�\���:����	�>�3�\����+PL�'����ܛ�2�b엛��Pi�-���	�.!B2]���)z�[�x���P�c�ۇ��6���|�����K��JԄ��c�>3;�����f�t��bb��{�I��Y������{u�����lZ�{�ds�z���<�I�V�d!(�#�"u�3�K�p���5������Y�m1���guc�W�)�L}�!W�-4�*�oޕ}�%����l�Ѹ��׻u"l�>
DY�K_�lf\�edo(��2t��bg.��o��woy\�9t�w~uN�/�vJ��9AY#�O�¨�*6).�D�g�Rq���������#���։Fxr{:��>?y���R�C���R��ͶWl�5�����(�Ww������!�A��4p��;lB��=P�����1,�~G��Ԑ4����eƑ��u�.o����t~�--դ�1� ټV�uF�"��3{K��������G��W�t��R�Mޑ���������GKn~?��UI���[���'���o���Ca7��{�l	�1�d	C1�dN��L���C�<���˟���E�	�7SO�5��"�����&�=���%��:�m9�Whĸ4�i�gB��T+_�V���� V�Sп^RTӘC �����ӓ�ə��vӉ�ٛ��W}��� � ^��yZ{�ZO_0���f𹫛S����KK��q��i_��!�Ұ3��t!>S!���� Z��yh�]j�a�H7�XE�t�u�v���V�p\�����g�ob��������z�^Ŵ�5G��a��&���;�S���	���\�E��.k�ğA�+D!UA;������M�L,�G�W�M��7�/�07�����0�����y�M���W��T*�a����Su�U����=-�|��2r��BQY�i���vŕ��7�й.y�68��:�qN5�M[�ʱ��˚�,�����a�n��Q$Z ��5S�m�A��HX6L������H���i9Y�n���G�VJƖ.X�����K�����d�Vd���/� ���V^�&��Y�>�u�>�N͝�iO?e��m�Y��X@�o@H�9����"����u�}9��P����ۢپ�!JD�v����{@uz�UB#��Sa���į�����$P�CKeL������_�Y~�#7��O�}拟ug���H�7�_�r�y$�������Fm�Z�:�Kk���^Z�����ߓT��6���MI�62Sli|��l�B���S�҉8z���vݥ6ԎN�j�������Q��ӳ�}�Oq<)ѾU��)���ϱº��:����Y���Ņ@.,�C�+{HڻY	���H��+��겑�!���l�W�����`Þ���ٜ^�08����b��eެ��_6���'�������ݯ��?~i�ߛ�M�_�/�k<x��#an�lS�RfT���'k����g{�]�?9m�Oʥ�\ ����9�!!�MΩm��f���$��k�u���8�=��f=��c�hӳ��\�J����E�;��gAD�+�XmnS4B�k6O�3�h4.�2����D ���hP�8�;��k}2uY(I�JE [�h��2��Vq����{q]w7�@��I�5�xMv`׶��MtE,
x� �>o2p����;)x\c2�^5s���x�{-�v�r�����N}z� Q�Y��g�7ü�)`O�e�^?a�RWw���:ɵiL�Х؄#�D�2�������W	�VIc���R��0�}{+-h5W�ff�9c�?r(��c�W%��F9�����\�߯�&��3=e�O�H9)�����k
#*QVR3D\���3��Q�:&6�v�o�<�����_�`��P]�Cx�h-/�4}�z��o�i��t��r�l���_��������-�������VM�[ 	�cu�A���W�ʺ��_sY�]éBb�C�lڥ5��H�Z�S����R���q�+T�3�j$�,M�r �+��Ѓ��;�Fݏ�A�.#,�,�a��e�۶��nԆ0.��C�h��KK������q:�ْ�8W!����(�~d�R�!��q�.�6�L�9AU�2L�����u�]eB�[�
m4k3�v?�f��MW!J��y�s�P�s2[��~�"%wz��HP��H]v�`V-��̞v�jQ��{G���v�k�S��kiv�Jzs�92\w�Ⱦ"߀�y�
�2mE������[�����r��W�T�pVB�Q���)D��L��*̝8��'��ϝ��/,=zV��6&��,Dm*���pu��5��L�M��y�����3��)�%Scr��q��!b����XCi��tǌ:��Z�U(��Z�����2v�y2F�G���I�3��=fG"�"��A�W�oW��6o��� l��ύz����}��Z<���Y�8pG��΍���ցyzq��j�����%I�z��zP�����n٪]���l�lY�>*^��ڐ��2�ָ��XU^g����}��Q;c��1����	�ŏxbdn�"I7�k[�!��[�7m�a'3��,�p�5� �4�EFC!}�&�$Λ@���&,;�.�E�U9��:�Ɇ���%��\QE*eC-��ȫrl�� ӟSZ=u��]-]�,s�:���F���N*�Y�"&�e�L|0 �>U&<'@u�,���u�z}��A� ��,�H�2�\��F�G��;��<�֬�r�!�T($;#�����&.6�؟���:xMi�4@��7�8���8����O�3\܉I/f�t����>5���|.։9sѕ�d�|�܄/�A��g�����q<I4m24R��)�%�ϲ���|,�h��AE���wN_��kE	���(d� �+�w*�ȡ�̒����WhW���iJmgB̡9��w�k�´D*�Ą"��ky���"^ދ�ףϒ��^�����ۆ�P�U���>���Ԣ9-8����vi������-��KbZE�ϗ��bqVV��m�e&μ`�1��M��:d�n���Nty{\ $�#���$f�2>�h�<|�b��,� a�ɷ���-7�8���$N?	��S�`�xXRc{��&�C�і���h,����4���}}�A&&�&l8	��5�(�~�ﶕʸ����A��y��P��Q\��D;��83�#�B��h��=���ݶ����0]����y?������Cw�Y�:�#���S���������*��
���̦~�����{Җ%[���j�*S�@�"��Bb��L�5�O)~W�D�N�5�o�{5s�yH���A���p��r��w��C{��R��6�B���t��V�i�T��A�^]m%�������� M4j�}�v��QM�训1r��rm��N�<w6�BZ+T�a�i0 M�I�*%		Y���OdP.��v�S�є��f�"o�����@yN����� a8e�f��L�����ra�,�w��x^�I��U��\��Q|�Y��{L�,�h>�)�����<��ި�� 1LK�>��	�9x�� �°q�**�!������td�!dUi=ϝߔ�I�y�T3Rldio0����//�Ѯ�엁2�W��lC�YFА�F�������玎�OҼ���EF��.a��E�(��B���)�MON�_���a_��_g"I�6ii�;y�-����Qr��fP����[��!�msZ��窱��F	TI��^z�B?��B+5�,�9�P�̡&�8�P�"i�d2P�h�����w  ��IDATUL=��ޑ�T�sJ���t{W�"E�W�yH�*^���u�֯ު�d#�6��e·�j#l}K��Ѧ+�n�-�r
�zr��c_ҚA�`�L��6H$3s`��
����M�.i�I�X�c[��_vٴ3���%U�[[LZ�����Yz�풖ҝxYV���~�k��Q�๞%��$Z&5Y����9;�R��v;(�cQ9[���`�P����NL@��J���Ü��]#��jӌV�rCmD	��B)�XJ�K��9#�E��6;�.�v+H��F�]X�I�/L0���\�g�
_��-�8L��V�e�-@��|q�A�#���w��J���������
�'�c/���g�M���
T��A��GdQ��e��)ej�%��j��
��������:���!�z��z�Y�^��o�:�M�ˆ̎�_�����f,������j�����We��K}���iԲt��������q�`'�K��؁k��J��m�ж�D��e�}�&-�PAe�T<J���u�exJ��䥱S�l�D��mD�u6$���"�_���tG'�SeP�e�Y~�f~|'��!mMȕ����̄��6�P.�@4B�<$�����Z�lg�(�4���ɚmC*�"�����G��v�y���ǫ��~g���;6��9�mȠ�8��/3��<��,�H�j�8�L�?���%�خM��L�{��!w��@�ȞIQC�Q�\q.�S%͋�GO��(V�.�W׾j����H���ER�g:�	*�Kµ5X? ?Zٷ���kC�T���u}fgg�?=	��^�B�8D�ya{� �i�4�U���Bم
=,�Q��V�E�8�s�
��_#�&�e��`��o;]bD`�r���Z��J�j�J5M��Ut�a:J�M���]gj��l�Yb�\I$&���W<]��A��������@�e%��xh�r"ӡ���j�_߽~��|˒?�V�:T��͵3�t���g�L�tkyi���#��K���-3�8�mp]��x�VKB��'l4YQ��)\2�Ȗ�j�l�
!Jv�30�hZ��p
Һ)�Mƕ,�r�V���J��عd|�O��έ�� l�(�s��{����w��	N���' ������칅r�!�*9phq�J	�3����z�k�����`�""|u#Ƙ�5�W �Ho�����!�a�+�m���1�৉��q��H��j�@�q���8݀:0���LK�N��G�'�����H�'������M��E���1���X��	[�zz[��|G���<�^��7o���{/_g7-���P�F\��k���f�{���D��t�)9Y"��%|���I�{�R��%������
!.�auoJom�Wj�6:���M�m�R�]&�����7�P��s�5&�������g�+��{I��\�ձ!�t�)h^JG�RK��(ځ��-����v�xxUz L�6�v��r�"�JU�@��e�������l`�F�"Ş(��U�p(�q�-
�l�)����5��Ŏ$�_�*!Vi��&��w�8W�q|�#S�F�4�?eӚ8�A_͘���`��(��J4c�y�,Ȳ\�c�;o�-n�W�d#T\Vn�I�h���
E�۶Y��Ʀ@z�r��7���ըc`��*�ix]�����w�~���~��E��U� �Ef��ۅ��x��gë�D�s�s̈́���p n��w���CoۆT�v%(��f�BGјP?(+�V���u���w�̔�v{��4���HL���d	�����@�� wc$5\��#	�47�8�s=��5��:
x7DڅlSE>k����?30���kR�l*]��z�]��q�
��'oh�׃7�����"��:�]P���H�]>�NVв;g���4e�&��^`,�1.���^�&��>k��4e4M�|��*����h�fij�+l�$�E=��Y9l���M���#�S��Y:��.*�ИL�L'�4F�
�tjF���7~/�+N+Y���pK�%-<��F�L�<(��8�^]���3�T��/��5�e��eE��!߃�j\���1�T��!�ґ��E���]W9�d����N�M6l�R"�E�X��E�-��ʛ1��	��ŝ.xsu��l�&J�bF׿�~�O���-$�іe�L,�R��*����p'7 �!�5��%ԛ&�xuH���=�Cz���5vSb'����|&Q
u$�)��g�-C�Z��06�GA��������\��܇�PP���$lS&�O�L�_�2$�>Ԑ�X��Y0�\\%Iƚ��H~�2Ok1�l�HY%dz9�w�/�Wc5��幱�Im��c�j�d�����"P�ޭ�-��#3�*e0����p#ِ��$iy��s#U�m�#w�b��I�;]#�HGB���3� k(^F���,��LY�F���5�4R%�~��N/��x��/EѤ���f��-�՛�
�ߥF��<e:C4�#��u��	>���9�~Uv��5tî�Fm�7'@vB=/5�rvsJ%VVr�s��s�m��s �Z�G���r��5-Ê����2��H6&~�9��UFN6A-�h�:�|�4&®����Oy Q����d����$����)$���a��.m2���>.l��>32L����6xF`��O�~���Λ��F��w�����E�����o��ۆl7��/ �
z���%���uZ$�6�ْ�U��C�+Krp�ӐuִTk���l�t2�A��7^m��yFƳ�l�:bF�MW�!��P����9��wB�C-��S0;����"��
E&V�j�5,;N���q���9�M���麞kZZ��uz:c[���:�KS7֙����8 ?������U����1BM��1��� �8��5!����[y@(�'�g�Z=B��4�p��	6�x�4��"��R2��-N�Ҿ��n�c4һ�N@L�xN�#�t��&�gp������a1�\ڜ�ܲ%r�Ҳ�ܢ�\EM����L1Y��G��8�,�$�҃Y�0��]���˴��}����`��LNԂ��gX`���h��Q���1�KH�yJ��vʦJ��h�$���GInx�NN:�a�[6ZP�n�>����z���h3��R)�\V����>����t�}f�ݎ59��z��7;�[}.ZL'��pqԉܣx���wnՌ�f�`��N/P&XG�3D*���B�al�)�E�ó�).ֿ53�me�{o�ڀ߇��yG��۫+�u�I��W�����!��:��<Co8�+�%�����8�8��}#��ự$����+_u�|�����Σ=��5(��%,�X���Q~G����Y��L�OB�����5�i;̮5 �j\#��*%���|hLz�3G�g�C�I�'�� zDܡQ��a
W�������(���$��D��8��r���hjFrO��((Kd�ؔut~�׃Ϩ��0�&�	w��{��{��.������$�j��I��s�֬���S�\����hpֹp��C�%���v����G�t�.�v۽pe�u�X<�S����UC���F� >+���2�Mu�'��5�[�ΡN&��u�92e�(m��)�l�>ӬТ��Q4M^�g��Wl76����Q���^x<�HD�P��8�)�EY��Vݕ�ѧ^p�Gam��꫍��&��p
7zt�����u_=]�~����g�P Zp�>�YH[*�T_E�p>��V��S�q�H��7A��~�}��Nm{^���yߌ�_CJ��s���H`�qT�];�:��tN%B���zgQ��|�s�#���/�:��ؤ
r��Xf�'<LLE}��"4�Po]^ux��X*θL� �'�-Z��\5�D�� ̸ ,�h� ���Y~$��Cvc�WR!������O�i�e���R^��5�O\y��G�G��_�	Vs~Z�z=��	���^K�q�����'s���Yk=ޅ��_����rs��bu]�rx-�B�2o��h���J�b�H�~���<��u�����oV$��MҵX;�P}>�&����ΐ�+�{2�������c���z��� ����f����#ZڢdB�>AE#�>�UX�M[%~y�sK�xG�B2�I�2W�0Y�R�%w5l����)�����1yݍʺ����ث[^�o���)\.���������i�s��5Q�'<�3n잶�^"k1�d|�_�e�b"�����<U�au}������U+cn��Ø�&�=�B�\��zmh�I�C��*c��h�c���J�'�S����3�����a)<�
���/݅��mМ��4.)v���fA�ކ������}��c7����K�����Ws�ާ�8�#1��d�6A�i�?
ҩʒ@%���~���u�����_� �`^��ک��!<��~q���a��y��X�A棦��T�sp���bq��A!��?���=ԍ7���;~��ڡ�ω~xy�?�gk/�O�s�R�I����$�ƃ�1�m��p���+��b��~�?v���K�5���˪�k♉��-4&MѪV�Q[Dag��ny%'U��Jʵ��$���v����N/���������}qݔ��N��M�����Ճg3r�z�I��a(փr�jdb^T�غa��b���O�}���s��;�O֡��DO��-.U����t����:�sbJ9/���/j���XL��_ʬ���_����+�����/|��h+����,)݀��v�'���VT�8霍�e*�"l�i2F���Q%�w���u��N���,�/�*�i.�?�m��@�7��p�g��NO�9��wR�'H,���Y�k�*Nc���}$z��ޝ��n����w���x�%��5e�H�[x�t:|~~>y�M7i�/���W���W���f�KK���nHO�$�OkqQN4�*��,��T���h{��ލoq"Awʽ�����\K��G-���
����^�����r����@!S2��l�������M7-��k��]ׂ7��[o���Ň��Y^���f�q~凬��%�^@&0��6xf��Fn�k�vM�u�]�v	>B	>��RE�p�cFY�r8��1�eoL�}=��Ķ�zP	T/Yj�y��4G�XsCyT	FTu�R"$��	����p)H̓�^Ӂxa��j�-��~�N!q_���j�T�'�>�@�HU4	�UO=���n����D��7�,w.����M%83Q�
��XQC�a�7�hX.�A17��%�2S.�E�	L۴�զI�I|ɫ�;%Y۲�-�l���Cܩ�M��K�d��妜YI��"�kr�ST�ȠΡ?]c���%s����Ϋߥ�{��~P�������vx�%�f&��Q�H?��:��'����/�<������lO�PG�nBw��aχ���s;R���v��H��Ɇ����hӏ�O��8�j��,4"c)D�j�1ݾ�_������V�����c�;e�ٳ���x���]4����]�;=���~w�s4�������`}]��կ��յ�1W�����������
	���_�4�?���n������4�wsC��m*�!k��:�	LL6���:��o�������j�w�$N�#c�ujq�pz�#���O|�+_�������ǿ�g���O/��k���;����̖;�U��%�F��t�_����,�~l�ps>pC(cs�FH����ȫb�{?�R>S;
����!adȕ�s_�;�h ;��@P�Y��x�2X�x��J4=���k����tV�4��n隙��ɨ�ז��� o9�<^c�H �3]8�1�1xG`��YH�T��d�y��X>������YI��u��*�4� BCs�y�mɨFBHz/��Va��;��V�,���IJ]��1�E��g�v0�,d#������nz��]X��	༾
^���u����Ҙ�uυvl_�������so���7�~�/���_��1��(��e\1�6ſ�e�BS��v��@��S4r���1�~������?�یS�h��s�������CGv� %E�!��Cqu�F<#��T��y��c:}5�|Μ��c����/��2�#Ox�:���n�g?�q���ή~ε�����P7��?��o��t�yVWR�C[g!}K�˸���f9��Z�\ش����R�S�l�7	F27ˌ��J���LŸ�3Wd��+H�N�y<��Kv�9���F���ϯ���6��i����y����&����N�b����,~Ҭ?wzm��-���'?�>��[ٵ��Q��Z�K_������|����Å�C1N���ح�����BojU��a&�\ߎ4�-	<�C�	~�F�t{/a�D_��W�O�����FՈP�s-ߨm0.�k�(����q�ց,z5*2�\>q�&��g��\k��˵���^;6y(��,��q����n;ԑr�8*]yuV�L���<Ƿ�{�ء����G�i�4d��٧�#J
Rn���A��$����"
�9���-��dՄ=��N��Efw!sU�7�&'��[>:?w���3q����N_�Ǟ��ޭ1T�j�ob����P;�������6Y��~���B���:B��	5KE"n	
�5�L����A� zf`��,QB����x�.�7��?�q5�G�����$}f��׾�ŧ������P)e�oq�z��J۴��|��������##x����bg�x��Ǣ���
4�>�8������i8<]��w���_�&>�{�w�N�Y���j�-T�v;LZR�gݐ�}�x��,zb���~���a�,xb(���9���i�Yq76x�3��$�`\4��fڥ��9L�6�>$��V��./�L �5���$���9:�aޔ7�_]i�G��v8���O�+u��>��+������#g�)�p��DR�+f&o���Ӣ܊ ���}!m�}�੩��<��L5�H���X�Q��$d�Z�(ik��7X<��)H�X\����Ignx�G��[��߮5z�>�31y]�ܺ�~���.F�i��*	�)&A�H����K����7=��CO��}F{��Q��3<�f ����0���f���:1;�ؐ2^����I�����Ù	ET[�a����`�����m��
�w)gj���7��Ö]{R��<��(muP�vmW��C�֣ZYxɚ�����^y5ķ���g!R�)�2�m����Lj�l՝z|
3aA�=J,�B�I�f�R�b�벝 �9TL	�-�=�����Q�>�Pg;��*���䬁���٬��w�c����cI�T{m�W�J}RH}��
��H�D�ӧoz`e�A[�c��� �[g�-�� \��~3�pa�Q�BǳY"�.
�lԑ|8��T����h�F�XF3I����%�S�`>�U[p�M.�h����	z5m6'0e�4�"ͅ'NVΠTe��m�.�B.L��B��#�YV,碳kϻ��tj��~u���o�o�����C?++ϕQjT`g|rj��8�&����<U�;�f�6���M���Bx*����6��V�MA��S�2���UdC�Z��[R6}7���'�x�O��^��X}�ƿ����yϤ\�vg�?Vt���w�Z�v!Y�Y�Q�����������i���^ii1�hw��PM��%7�I���U�tɲ�:�R�όTRE\�JH�����"��)q*hsU�;[�:�h����J�m]�����[�`*��Np\Yyb��?�:^�����f��K�[�r�j����ję����"!>�J���Ժ�ۏ"qѱ-�*KY�i/���aU�:,�6v�D@�q�{�@�`�mE��jB��;r�¦@S���(�v;��Ԋ���n���%-�9a4L;<{�~�v��E�Y��H�擐���6a�>�fQv��o� �\;s�Z�0w$�Y�a�ZG������nf���Ku���U�q���D?���l@vMt2�fk�0I�
]�W�5��6�$J��C"bS�����!���ՍTsr~��ptRd�t��'�n�֮=��o�����K����{��O���d����=���$(�/��N��U�y���������%�ӷ���:%��jh	���r�⧙"Ӱ�&y��Mh�<f������q����_}׵�~��tx�Vk������H�����b���Ux_[=s�-O Q�;(i�g(��j���h啶q���B��R������:� ��a��w(k)s��It/p㩗6W� ��t=�tV��7q���+ֺ}or�g�!�Q"�h�l�tb8	u�N��������P\JT���5�5"�J܋�h&�(0�|O��!<a$y�&�`F!�'<�m'"ݧ$�P��tc��)WH���(��:�]p�_G5揫����ך	�|���e������s򑀣|�dw���7�w͏y��u��U�g}H��tQ�Ei\�!&�o���t��u���P�sf���N�����F6xة�W).�t�<K�Hg/ZF���ɪ/�A�e�:(( �"8
��0�f�FS�,��1����Ձ��Ӽv��Ǌ��sn���O m��
�~��Kwf�;ꄩg1
���}���c����=
˪[U��'��������Ifff���w�g���]��"����˶�ٔڏ�d��H�����Ws��������m}��.�c/n�j�'�N��`	[=%�R���\{�����#�N��Y�+���-����� ��A��9-lʹ�՘c(s!��/��re������Np�|0���3VR4� ��i���ͬ|�Zؔ4?���3qp����2�HX��5_Zl�C�#H�L3��:�9���i���<	��7�2���Q����5����H���%�C����I�R���uh�!J�	<��#�+�s����V�}�h��d�0�)�j�&3���i���!�ѭ۬+�����3_�s��ן����]ui)�@t��!bI��BNޑ7� C�]�d����)P
�eB��t8��@\Zy���j�=�: �0��T��+1���67�ࡌ��f,�qλC6xK��O��L�8v�P=o@����"dP�K����RH
�'	a����NX���Ռ����#W�x�u_��մ��ݮ�����eԶ&'<��E�u<7��s-�?~�Q4{wT�D1�y%@�٢�e��J��)�G�/GF���p7w�HG�?p�ؑ���a�^u�>��2���_�ڷwx�;�G��Z�g�k���{*�.Iөxi�� 6TVc�#8�C͝A�:Z�2h��m{BfS�Q �*c��1����J��B'��Y��m����rԙ�pǒ=[�v]�wΚ]`Wc��̉Ss2����\C	��Y��FpŽ���$�&]z�L���>�.xu+M�u!e��(��F��93/_C� D�:嚥l;\]�׉o}�C"�v�3��'�Z�3- [���#���A����s����$�|jy6k���Mȯp�2)�U	T���ȠX�ao��@Y�'}���A��rKfͳ��Z8焗NX�*@"��2U�ϊ�]|G���%x
��)-�gR�J 0��*��M#�R	�J������M4�LQ�LcB	|��=bV���B��t(�v�Z��`S��k����p���O�Y�>������n��{�u�=�~�:PK}z�3�	Ɇ�iJK�R���E�<�x�9���d�6xSc5�l4��!�Q<xc�<
�t�֧?E�t_��P��$3���CB�ǎ�Ɠ53Z[���Wo����s�?]u�翥n�q���W�m��ڭ���X�z�7��n���x!k4�:/ٺ�o���㘆�!���c�[���YJ�����8��=��\#_d�� �^p�6�Pz��f��������W�Us���tF�/BK������G�G�R�&�#_�&�$x�]�b�iu�O�VP�����9�� �R��>�$��>ǿ�s[_���;�]+��Lsv��z�;i;ڙ
U���a�*m5�u4�UH���Ǳ��~���, fWl��H��t8�����8"4�L��4��+�놉1Ӱ�x�Y4E��56���x�k%��i�V?v�����I^G�Ħ"�,w ��92w�r&<�R��g�:{52�l����Տ��!	�����N�������u�u q���A66b}���f��;xm�ǿ���cώ�x��1��Şa%cs�BB�`��MK��������"�UVUVVU�$����|�^�xq|���cF>�ˎ�Ǹ `�1�<xd�Maj?Cжn;r�l�w/��A�_L���C�i$o{LȘ*#�����8Y#nXG`��LpĊǭ}b}TyAFG����e�Rf:/���'p�š\8^A�,�A� �X�69����3yڿ�U��ާa�glz=옝%sqJ���&�9uF�, �@4n����`W^�Wuυ%�^&�y��[��/������|���Ŏ��?��P���ĭ����V���bO�j��;�_㰯���3K?Nʍ���ʤ;w���S��詓Q۝uzq�kǌXZ8�8{��Z�#�Ѳ"���sN����+�usBjM�Mc1:�֊ԫ~+~�5yh�2��l��L{��9��5+�L���G8d�q}Z���p��L�Y��'����76qk�ԫJ�i��Ѵ�%�.��: ,�t��c=>l�8@��f4�i �q��V*t;�[`J��$�� e�N���k��5Ҝo�Ȋ.y�6�Z��򩗽1%_��G�@�Z��:2�M͐�]$)p��x�o/�����_��h�z����Eğ���"��E�r�u��S�n:��t0<w3�yNa��$���-��p�Ӽ�*�@�SQ��Nu:�D�R`66��3�Y,�$B�5T��Û����D�*���э��a�Z��5^�ˉ�\}�\��I�y9�y�'�W`�, ��(��Dy:cTb��	�Yg�� ��)��f�l��°�x�ٙ�G�������z�=�x�W�� ��_o�:��G�c�ħ?}���E�4}��2�g�5z�y�f�gϽ����3U֫��m+�YNT+�ʻ��X��Q?J�^T?k��v�~�l��x�4l,�$���t;c;~ 2ë��gz*�[���ǏBh_��b�i>�4q$�^7)�*Ff-�Oh
�5�E:�i1M�SO�}@��",�ڱ���ʵ�ǠkmP��KQ��ӝ0%u���������\�7�*���FZV��i�Q4al�t���$�"Dݣ��4QӔ��eI�Ԣ�Pz��,�ݣ1Q��HRkJ�җ܊���v�{w���06�u�Ԟ����x��JGRH�C4Mw#0�N�ĪZ��Qj���J��,�z��i'bT#�`1ZG%<�*Pk��j���LG�G@�%�mZ���lL�^�A�����Œ���
�B`LK$Iƥ�)����\E���L�ע��R�T�S��-婝t�$?4D�J0�u����:��E��n�q�kX	�Iy��Ҏv�4<$mf�ê[ü����w����}仏?��o��[���6~ç?mU7����ݠbj*k-,�_����6Oi'�9���*Z�W�铱���]q��K�])�Uտ��S���=U:C����vUHz҂�����|�<���W�T6������e� �Z�p��#��;+n�*���i��%|��������b��p�-��
J��bs�I@N_��� �*7��b�Ͷ�8���ʒ[�~	��\}O*��e�� �C��.(94* �C3��&�y������lַ�8��W[4�*�J�{��6u�j�>:�l��ٳ$vY�Y�k�6� �^���8}2s��ä����0�fw��M:-�9� d=T��Z�x�]�H�-�s�y�-����87?�ַY�����DG��Ӝ�<N�,L#RAMNN�������oH-T�	{/o�`*iL���W��m�+:;��$��͍E�l"��{��� "� 1���E;vNe�Sі2�_��|�e�>˘^����\;o���*���׃u`X�4̴o;�/1��#Y7l�9�(��!q3�!�aS���RV�Չ��.�˽W�c�L����׽�fy�Yw���8Q��M�2����.�?D�>��ԭ�?3�V}��=H�G9�}ό�B�I$��t��3����J����0[���"���:�!5���J�c1�2
���׸:�f+��Gm����-��_�m+s�����X,�FS��F���L�V���G�}�+>y�����o�A3O��	��[������qnݨ�ޟ��g=z�Wf����'GE������������-�(�S��u�)��}��E噑�Q8������+��p��(�g󷭡��PѾlt�l|A�����{ܨi�4���a.%<�t�Z�w�~k\ ��x,z��X��4E�"���S:K��)�zj�*k�%���4=��ݓx�
�>5żvL|'֨��9�A�I� �F�Q�@����]�4F�h�}�s�nГ}�(4x���&oz�����p�C帾�'i�j���k�A<�oԲ��h܎���eS'4j:�;��R���Z�@�����fרh��Iȇ?�[�ڗ~ڹzz��~���v�q��� r�Y)ϫ�����~x�������`����x��~�,�rǿ�M��.3��P��o�X2�
�I�\�骬���Q+56�P�4�/�@ZX�.��p\�r��@�&��y.d�YR𓒈�4Bm/�s?��^6���,Ϭ~��4N4MOƪ�Ӝ�GK,{u;�~_�I�5qC3��O��Ϻ��T�=����w��f�/:�i�9�V����=,9$��}:+}�����6}�$��]vi޾�'�	�c�4���u֟�t,,�j��4�((:�Ғw3�	����'���P'ؔ�T�P� U�&岯:�!�:e�4�:�
�[t‑i��������d�A�iK�}���9k��P&���j�g$�B�����$�K�3���-�hJ���Uxr�]���G�dg����K�(�W��D�HYD��n�'��/�}�-� N�lv���2�٫.7��3~�����5?хw_���_�?�����c�JJU�DU����E���8�̶�{vr��w(�g\�̧�G�,�6��!�i�y��l��+C�mk�o�o�l�Ȫ�:���hs�0��������!��R�uM��2��(�L:Bo
W�	�'R�U9�?�V��G�㢔��SG��x�V�����d��]Q���"�!�*Q��j�l5	X;���hv:�-N�qOG�	��q���NM��D���q�|畯{��W��Ӵ��X�߿߻�}��KU�K��Ɖ������ga��s���Z9�뉈]&g���8�O�%W�7���~���i4t4.���h�6q�u�#V��������Sk���Ys/j_1Z��1���֞d<�ۺ��%�n��2��Y)�zq�h3v��#�� ��DŤ�:n���I"xb��%N5ֿ��]mH]���q�����$@�W��B�<hc�glӷ���\��ܼ.��	���\��x��\T	z�1�」ޓ:ʗ�r�E����2��������K/%���|�V���VՋS7q#&p9��E�?����و����ͯ�7�Y��z/��mv���d*�Q?�S�p�ѻQ�Q��Wi����#U/0=V�C �P%BDPW#YVP�mI����L�Ѱ�ݷ_ݦjCJ����S4SL��%�r�.w�Ա̫J��0�?�� �{�	sjN�R�6�e�\r��79�gt�UP��G��/l�	$T�ecM؉@!T�����:�wXǉ5��K�`�c$k<�H�)��نZ.o0��jn$?ꀅV��GF8R��K;��w2
��3;��7���[�N�W������K���f��{�[.W���K/����8��-q9����IB�DQ+pyg�ƛZ��\�2Ȕ�c�D���9��KN�w�S�#�R�r��>㆗D�r��"��hdŗA=6�h^A�q7zI'�FJ#V�ˬ���3�LZ����	<��O�t������P%I�G9���*5�2e8v��D������2�o� ��x��a��@*�Q��v�`)�j�7l/vٔ�������h��3/j%=��@Q��E�V��E 7��^x��ޙ�RY�IS���N�����v�hV�}���Cq�#��/�S��K�:�W���U f�J��T=�t!��m�8�����F���|R��-eD��Z+�d�i��N�<#ݥ�!�8�O�Љ����7i�̜� '��(�:zt�&p ��>�X]h��ei @R��f���FB�g&(&��H���@�ą>�Ja3a��Ѳ�����&�L`�E@"�n`yN cW��t�w�'�E�����Z�Q�y�g<�zT��}W�y"�F��UO3F�{�.��Of��~;1����r�FV���5�z��֝�R��7��H7}��KF�V["��8jAqZt[0�{=sޛ���]p�qE�.gw=t���^q�5�0J��s����E��sOe,�_q���ԉ4�n�{$�˼ݪ�y����S�+!�^�Ȋ;#r��TNK�6����+7)X�DD���O��
0�ֺg�)jh�Z.�&�HR��]�n�x���&*�PBMh}N��;�`ҡc�zKp9�@��;!)���]���.�t��qN�J_�6�� ��`�"��|cI*�G�1fרB��c�`za�����?yw8�"+V���V���-���e]l3*y�6`.`�HTS��8���9 F�ԟ��p���Z��?%��I���-@�:)�J�Z+
'�m*�c'J%9�u]+�M�S/���ҟJC-fwʷ�a�M]��R�ɮ)�?x�"��UE�4衇T�F$���#d�� i`4ʣB&�7-������y�k{�$+U~�%�ᳳ=�����s�L��sӅ�)�nr�6~��N��<��{T���q�{&�
4#ƊQ�cXX(V��
�&A(*c����x��!���y˴ܮ\���n��;.��<��oy�{O�:��tD����9p��lS�ۉ�_��[����7̠�7��P��V%̪�%ԍ2�Hl"�˺z����d�o�v�nE�/��v�LS��(�j��*fE��Z��nC�vwDv�C�ҕ^���S��@��r~2�'I�5��i�1����S3�=�<M�P~Eu���'4���;;ERu$�.k?�Sܭ{��	ĪEd�t�,^$��������9��|�M+����,�Al�>�@��
�3Ld�dgM}����)ͷ�)8m俕�˳�͸���I�N1�:Z�,� ��r�8�H�+�1�[x��@U�Sʄ�ls��"�* ���O:��;��J�k2�渊�/b�A�4N�O�`tH��ia5�|�&k�\9{�+�|��Mr�}�e~�P����S�C��`<H����.0NJֻ��Jj��m�}��JN���`��z����W.��DǄo#gƝ�$q�y% =� Z���z���^��o\�h�_�{������6���=�M��w��4;mtƯ�4��uT.�S*=���]�O\�I�@ ;ڃ]iU®�<�Dl9��G��Ӣ�5A��a�Ep(��Y���U�{P�C�4�=L���J��*]�����]�9YX���<��X�9�F��(���<�d�t�E���ǏgY�8>��7�+���#e;Q3D
�@���Ӄ�7c2U�I�R"a�H��2�/�鯩��f��V�K�Y�����U+�He�UW���������c�V��=&E(��~�*V?��B@aċ������|�uS�.ll��T[ڡ�N���`�ĸ��t)Bs��x@�Qc�����dL�Llx'�vM=!���hoz��}��O���r��\,D��֠<:��)�I��$�(ZϘ��y�j/�B���'U�=nP�	7ɑј�=D�3��5�T�(�m�ܡ�1Y�cu�F'�ę/������F�����z擷��[v���8~yujO�CT�B���N�9K�����:?+�o51ׁҠ^��2)3"$-�vrdo�f�&�t:�؞w�ד���F:P�nۊz
i�2��A
1�a�T䥽��?C.��=kw�ѓ����5���z� �,Cu���$�%B����{Wrom��6����we�DT�a)�`��27�u�>g�O@���������+w���HV`�<��A��@�hOK��%5�^�9��"0c@e��6�O�O���Q�5�"H����y�;�n:�d�[*��d	�V�Y?x��s���K�D�ԏu��- Ī5N��$�o^Do���]��s�̝�W�9r�s�?���v;��~���.����i�x�w��FA�@�ې��)��B,(E)=e���[�ڐ��窷����0�9�p�EJb�K�\a�d�B]��=�)�=и ����<L���|��pɢ���~п�ػ7��|��)��p��8��c��q�Y����z���a`�� ~�؎��ۑk��(�Zɐ����F�����׆6�3*&���4$-�#t�Fm�!����e��=ԫQ�a���_(=�Ww�_<��7����i �z�":w�'���Cj�8�ڏ���=�(����<2���;r���J���z$n�%�l\��3C%����o|#��-�H�7B�#U@
�9[+E���S�y�bU"e���qO=FX��"g:��鹣���`M�@���HԹp��X	.�:D�!Q�prp��/��9MT>eV�2۠h,�\ń7�5ݔD�@�J���:���&сr����34U�"t�f��~�W�x�����?&�=T�/g/�a��qv�:�+��7�x���~������zf���tʾ-���CB�1���Pb�W#dPC�z"U�;�Ū�v�/���o] ;���y�������쒓����F?�8w��k���)^�TVyF����w�K|�o?~<)��KS�^���zcJ@JW��ے{��	��Dڋ��(e���ϙ�{p��M�G��"�D���+�=�N�3��w^���ԯ��F��o?x��}�`�92�����BO%�8T��Ih:����ԃX��'��'�+Za�7p��X�������0�.C���7é#]4h"�pɳ����bK����P�-<x:ڏ: �~�u=۳������4�L�ʖ��d�Z�Nƀ��ɄpK�"��Wz��UaT�:ˁ�.m�D��K1��ZQH�"E���7�_���9��)Z
9w�@�f��6F��YTeD��#�;RU���$yH���k�Ͼ��o8��`O��K~���G�p��;w���=f��%b<�f�b<pM�>l��O%�TIٷ	~Uh{peD	 Q���\U�1E��T��
�	��V� ����IZ&�%�)-v.���{��CO}׵�G��µ;;�o4�/Ȳ�;gH��rQP{��)�+�(f��@�:�3��
߻h�.��k�'1(v�����W�{��w�]��Ǯ�Ĩ�:x��ʌ9x$���sȌ�3lf���v�o������ h�w���b/�>�𿲛�U:O��_�������v�|�R�_}���l�g���ׂ�hx!N ƨ�'�$$�.1i�]�nvȋ_�Ju�>�\wc��d��>�U��p�I�u�\�V*�8��^ú�^��W���<h�࢓"	�p)^R�t�]w|��x28;�$Ij���c�5���@���I��SLl���f��&9U}����)y���O:��M� �FFU!�
�1�Y���C';�7�j��O{��(ݿ������w��/v�����̫��k�+���'��M�]T�3�����c$����5��CDC�-��p�e�����@'��v;�����/?���$"i��t���]�&i\�F����b�W'��=���zOe_��A��G\S�!���3� 'nv��3�#���ˠrs�̽��9����:U�ۦt@_C:���j2`k/���3N���"��K�Q�CvEbh6HD�4���d�ÖM�m�?�`-�Op��4��|hW�`�ig<�*7����i=�Z���zi��c�V�漐��N˗�a*C�9�y�WK�����;/�p>�7~��i�^J��oJRQ��FG���
̻	�2��a��q���"�w�*=���U��Gԟb�!����f�m��g^�r7�,MG���Ut�K
ˡ�Yݓ'�)}�����B��@��F>�q�>Lȑ�,�,\"<�<>��ы��Z%O�(����H?=�$zѰ!���1��b�,N�Y�2��.9���ɞ��%���Y�Ơ���S�����':�����lp^VKÔ'���'�Z��R�v\�w���t�����r��Ou�����6կ�<�\�x]	���S���������0�iF0��5J�a���#�[�����������(���0\�8"d�^'���@����(L�-T��.�́mcҾ�����{2:NJ�i�+ܹ�Ř�ZVQ0��5�����<Ijӌ�͔.=~����]�G|�]w��]��Cӥ`^����N�q!����r��#u�#-�/~^?"��-�WB���7P�DC�J��`�^${ά�e�ً~�/�x�{.8�1J��=ן��w��+U�R�g�sww?�'?�;���~�����fZ{[[:;���� ;y�T���6gjk'�+�G�*�s���;���8J����k��:� <�yAg��6�A�Ьv��4���~@ϫ�T���i����]ic�'��-`D�{^��̨�uhn\<V�E3f�9�b"�wT?e�UьC�bDW���a�v$)+N�i���Ȃڿ��O|��n\���ܜ��;İ�~�s�'�g�3�ꡃo=�W~>�k��0�5%�����l�L�����,c*X"��~�Y'�_RL���k3`k�����E{рl�|�=��zdf�'���Zs]푘�C�iL�W�RpĲj`�g�AQ^��@�}����,qȎ=w.�T�w?�ҫ�����>�9)��I��ʋj�Nn(oz���Qo�I��cVc���?�_L�Q�;W4 �#Ydr4n{@X���e����c�/U���K19J�޹��������?ybgF���NR��fJv!�)`="��������%r�V�e���>�Є��m��Ɛs��jU�k��J��B�XsW��-D��%xB��q�C�ڢ`lwj�FFt7�:R1�0�$�S�3���G���M����pG�-�nz�d��m��+�	DJ�'=��/���"�������04�~����o]�z�����O���óϯ�|Q����0~�5�܁گ.�/<���,WL�h���!��M�fg,����-���Cg~�U9��^�Θ$�N٧2��J@�>'K��� u��D�ޫU,Z+��.�cQ�=^��_��+�+{X0�d@�+I� $�':�=�"��tv�}�2�}���_�����#�De�c��!�.ٸnV9�!��T����$䃢�b¿s�y��G3y���űI��rX���+V���_~�ʺ���o>u��k~l����~��E~�/[���S��򞬽<����@�C3�� *a3ӮrZ/��m��H�Z���Dq44!O<�Є�~�`�#��$�ht{�:r!1�8��}�A��J5Ȧ�LEL�� ��(C��Z�zme
�|Yu�T`�M��Q��LCx T�h�~�����N5a�y���0*U��c�E����)Y�	�����/a�xJ=�����rN�DR�qE��(eƋ,dc؅�qs��3cq�)�Ӷa$+	}͒e�m��_�@$�����VK}��'?�d*c�YX�8���3�!i����\�R/���rε�8!	F��Ą��!l �$�Kz��gw��'�Y�=t��-���w��W�֗�����T�u��K�ob�
Y�&4�i�uS�m�8��u�X,�����၍n0�*���m����πC�QRΤ��r�r�S':?�&�'����q�R#i�p�(�:�sfN4;�ͬSq��&_�5��G@��XWgrἕ8*$�ߪH~N]c���d�t�E���x��D����۟�b�HhLd+�Z�_L�VB �d��`��x1Cj�I�M�;.%fr������ƢQğ6�oI����z��R�,���Q���{�#T��i"A���9r�SrU�I���-v��^�b������!�l;��Q����iv�)������Z��9e�$5!����In��k4�7��.�?�3�Iiˍ�D�vX��f�I�F��mpWv��A<�����%|�}��V�;#.��'�L�~�{�{֓��NS�����=��E�ɒ��\g''3$��CP�嚶S@ౌ���E��qN��ɪ4��9�5��T#F��{H� T��S$�R��/���Dg|Z�}���T�����8�����(I���h��P�Wu�����X�3"�.���&���Q�#����q�-�F\2���,�h�?���"��'���{�,��3tO23'ya@W���4�5\<��:��rʮ��ԫh6*�y&@֢~B{����1n	1T��8^:�k�(#C��jRjT��1x����%��CR�����������C?�s�,g�V�1��ܕ!%&m��5���룳�o�E(:,�mek���y�q��Jå��"D�i�2 h���9wXA<1�LC	d&_�Gh@G�|�h8��Z 1���8PVU��2G��$�)u$���4�����N@b`t֩<�yT��V'�h��h2��=�/�+���J�WCFV\�ex
j�;C��=�VA��z�Xk$ �m���%SJ�]l#��(�xR'��� �t́�}F��}�P=��F��I�a<25��Z��6�A���@���]�!�U���.B�w��L
�f�Bݼ�J"`���l�n�V�^@<�u[/�*ӕ�OY�gC��h,*������D_ŕ�s`\��=��&Ф<m��"�$iJd�dG����4� ͹	'��&�Di����[f6*��o��0}R�z]I!�\��y�l��<,�� �P��+ύ&�L
"�PcѠ����D�0ƬK8f�O;C*�|��!��h"�B�f���՞YD�V�Maƴ��{?p���F���EH� )��)"Y��Cz�\%���q�,��q��%e�GT+im ��	�n��Q�˂���u5sb�j$Y��:�������&���M����6��5�D���d��2"vbBt����1e@�*�I��쓩�������|S�$"�,4L[��׺E�1��".<�b}G�����MA/�8��r���nB�E�fZ�T�o�\�į��g���-����(v��r�Fwi�|�:��|��GG䪚lP���Z�K����6w�{1'+-(��|��[��iH]h�XJ���
\w���0@i*�A�v�Iõ�HUhօD��\�]����I��v��u���E������j Z����k���-�ҶR(8y�*l�1T3bP?�yUx�ܽ�D�$1u�Õ�݄1��zde1����Cs`-�Ar���ɟ����@�2Lig񫁂d*ԤfX�'>��.��ѿ;���F�
whqL#��^�=�j?�x��Tk�I(7�I�&�$�r��e�C��3Lw\dkۘs���x�M���ψ�~��B�W�g���]Z��	u"(ӪON���OԾ6�:x��U8�099ܡ�ʂ_N�S�2އ}��A.����e���#<jR��c��vV%��`H�̉;�~��<�G���VO\j�~���d�m�?��aܑO����9y����ԃ�� {�F�ˊu�h�����zR�iF[��x��3��#���v���ER�I'�Th������P�<�9���5ƌ�G���2s}�C^h&��Vow<�S��I��#2�ȧ�N<<�\�e�D3�3O�_�SL&�-D�X��&:��G�|�ϲ����P�V�����ի�lXm�=��K��sr��,_1(�ߖ�?�Y�X�R�jhj���oHr�0�n����+���E8���뎷@�
*4S�L�W��j�R�*D����yzz":�qs�YB����~�� %*�ʚT�:|)O��ZUc��Rk:ܵQ1��1�OkiB�5B��:׎k��Kq��h!/Q=V�y����S�1��J�|��y�Do�t�_aĂ��g��Z'��c�Ȋ��H�כ�:�F�����z�-���n��z���K���(n�J&G�)�SuI��yjz�_#.z#��.��Z
��4�"z�a��_��B��A���j���]���ښ�ѩ�D��1�������ۥu���:���H���?���vA����86�*�3-��l�@��E~I!���lV�Z�3�{���R�Se$����%_��M_3(L��¼w��1�ZP
t���9��]��{��η�G2��}R8`�Y&�E��2�/7�E�<OH�?=�hܮ�,Wﴰ ���DO����܆��d�,[jJ#	�3#�� 3��0��h�����J����ApE" �-�2fNn@Ȇ15"5�5�_MlѠgr5�}�o�'-!y���s�B�%ªW��:k�&���]��'L�oh��Y�.i�z��F)%%W�����/�������	�K;��U�щ_�TS,�sV�ˑ��V��>��q���d�t��)ۍBe��I���v~�ɕ�Y�!��81˓�b��u!:�Ǆ#�krdє��ES='u�"ۭUgV�$�t�T���ד���߀K��٭��]�M�C��a�2&a�o�O樚�>/����=���l�/�����,W�L�$9��v�#�;W�] �B��7q,Tq�L�<�m��c�g��wL�E�c���B"l�	k-e$P�:��?I"�a��c�M�i�9��c�� ���Z仏�����Y�<�np��}���Ln�h,\�扔�+J�20�I�X����`:�i�됋.D����:[[���5蟶���܂ie.
_�J[��g�q"�rق�a���&��.Neq�R}���:'s�1�3�!&<�*fr"�ThG)H$4'�V=���~���u�?f�3X�'ﵗ��z]�C.Z$�̓�o���noc���j��M$�V�.�
� K���b�*�2K�
ENC����~�����dr���շ�|���9��1�QQ�v@�-���r��TS2m�2ēi�_b�s̾~7:Q4��M��bŃc����(�+�]3͊{����}d%�/��u>μ�����W�US�e���U�>����P��huP�Uy��<�K��t�L�X���x8��"��Uy��>3Ku��gS��;���Z��<AݺV��Pj�3o�$Wأ��1G2Ǒ���Jc�~��9��Q�Z��b�|��u�����q�ϵ��.��N�Z-�hB�
��N���q�'u�Ϙ�F3YtMv}�^1�6F\ZVf��Jo'0��'�>U�]���sK�7{$CϢ[8�m<��QV�Zǩw�X#t����-��zC*��5����Da�nvF�Pq^���o�eX�>|4�[�:o�*y.����}�@o��GR�=fY�S�,L{Wo4�鞄QJ�8$A��h��3�V���a���:Y&'�0��U[���J����X�ڔn�TO^K���U�a{|���'Q��>Ւ�X�RG9[_n�{�r� �1\�<c�3���+�3�s�ź^K5����r��`g�ʺ{.�:��;#��� � Ú/3�F�rQ��cm![E�73�cM�I���j�#7�@9w@�U�?]��#T� 9q94� 7u�Ί\�}��l�Ml�fo�l}q��c}��	ƌ�<'k�&-�X�'��r.��W���F�<��NN1B=��gn�9G��DbYn(�պ�v��������ߍGXޛ*�Px��9��J��n9�U�X��	�2�&H�D���ۈ{~�Q��߄.�r�YH�Fs�J+�~�oΘC�z����ld}�P>R�^�[o�瑈m�`f1�7{�~��n�D8":��h�|�%̞�������R'$`T{�A?�I�Fd��A��ps��l��7M��#!ۀ��e;�G�D>#i9��U�~�^�hzӾ�CQ\��a�:eb:���Ȋ�6�=�6�W���H�p&R�B�0�(6����0�0����=rZ<[6�f���(6d$�8�j�~1����3��gd��@\V���8*�;:[8I��p+&5�9���N�~��I�����4��ba��9��c���V�+]��ub���h�M���h���|��w�򩌻֫�CB��8F��鉛H��S���T]�s�ly�y������.}퍣0v��Z�rs#�g�="y��V��r�w��1o�ڼţ0c����V2�M�"t���xJ��n�:H(�F���M5�ʋ��z�I�W�`���ڸ�����n!��Lhoun��@K�rlEL��Ѿ5������M�+!&�M�*c�hFK����Q\��6L��_,�P�T�=J��S.pH'ě'[aD�w̐h�I&yg6
�>���Y�'+/�>\*���6;����q��}T��f�c@~�i����s}��Y"�4�B*��#(�}g�>Ee�3�Ǐ�[�TJ �q�YEV]�G�蜙�� ,��a���
� �U�~NH�*َ4Ji�=0U��~e(�ӡ ���Zug0�p�+�b�.R}b�c�H�wH��aVvj�~t��\����SlƑ��7�����N�GI�<��Vd�_2Y��ʤ�K��<-.�1�j.	R�y�z'�
󝪯6$�lg�����٨�Y����D��Si��ԟ�%8\��%*�j�]�)�i+�ʉ3z��Lwn�OHF��P,)�R�ꂖ`LzK}m�8՝'���1���)� u�j-��5X��;�c��k�8��Z�t��{V/`�	2�c��ݗI��I��T�u�/{�Z�(&xe�r@�pX����:x�̹I涓!�N�󷓵8iq�1����ǳ$;���3��;��Z{�(ieҞ_4Q��ЀD���V|`��Gb�*|$�������w;�P��]�K\��T .��%iC*B�0ժ�z�֗���s��M�q����b��I�JR� o��!ˡ�#�.s+s��0wmè=���m�.��@��u�IB�#.����=vg ���4�,N��Ё�=\0[S�0�G�êB��0Q$J��h����YEr6W-?ND�9��O�lS�f���̋�ӧ�i�^���p����))O��Pj�yi�u���d�#S��9U��b���RV�M��i+G�?� י�*[1_I�/�.N|
ҩ��n����N���K^&��·j5Z�z��MV՞��.Iͧ�k���r��f"$��
p�1�u�t�����~;���O������j���럵���;��y��C����Zꆏ� ��)?�(9�]_�<�\K���Mڥ���h�Zo�o����RD�Q\H�	Q1R��w�%�ݾ��+K^QrA�����D�^'���P��Z��]Š�5���a`S��LX?kĵ+������I�8��nɝ[P��D8Q��6�L�,�"^�y ��;b9�j-�9�x�[�]���R圖��
	Qk����*�8�.,(���=j�4��0ٶ@"}�Pe&�����f�M��yEEne�����z���F����k6D�3n"h��!k W�<��uD7�{'o9����~��Qtv��*{2Z5(��$2��f��d:_o�v�G�)R�5�L��(���P),N\ ְ�Ɵ�3���ZG�WWL��뼤�@0k���?���~PU�0g��#�RB�=u��Ż~x�q6�p�Ҝ��ҖI|�Ut��7���D+����W�(M�ܯz/o;�%��F�$}�����̙1pk�e�P��#�句`!c�J�
�mT)��u�k6I�G�H٨?�R��w��}�c1��ɴ"�93�}+b�v�<������e)5MS%V�ﵚ�������^t��޴��ݠ�ϞQ��Yz~���uR�(����"ub^�p���w�ڶ��<n�XW�q]Z�~��62�0��ӛ'�O�:�	��8�����"�@sv�v%����ţ^�������ݲ���y���f{��L&�V*��aó�,��kJŤ���c>T����R(J�q6���E�2��M�㯔r����-�T��:lG��-O�E�S�>��ʸxڣ�]��������?�؄�~����v��>q`��s2I=�<���2����_��+;��+��+;��:鋔�$M/l�ݝ��ۏ,{�n���~1]8�󋴴�'Y/���d�_��'D��v�c��H�QG,Q���l��qţS5��3 fh�����w-����F'�w��!�j(�c�}��u\,�:��r)�y��Lb!c_j���'7>��p�L������={�%�o�ز��y�L�!a7��圉�^Rz��\��`����"r��y=��Fח�|N��%���ƻB�
3j�m�H��1�I6�X^pٗ��z	ɋ���`���\��6'�V�	��c�S�I����p7l��eG�;�ސ�?sK��+�kGc�������1o�XJ1� ��M��a.�I-.$#+�1V�����<�F����(�Ċ߬�����Q�qŃ`q9�.f񷞌o��܂�h7���=��de������r��DǳY�������3���'�����w�䟋+��=V.׳��J� `�zI�Su/p�6	�t�iU�`�*�����3����V�d�y�eY��p��-�Df�!T1#5 =8:����|��Qץ�L�� ������F)I�J�ɖ�e���(ĐR�ρt'��
;lN���{܉i�3��H�<�i������3���ۋ�{i��c�[4w�2Gg臤FM�g���H���T0��{?���wSz�wƮ��{,K#&y`����Ƹ=UH�Z������>����#�4�Q忓�y�e�
+6�LH�l���|�d�X�t�������0�>aCg �:��Z���m����\EN)�+��6w����O$�r�D~�_&q�֭,�5暖T)����vɿf�3%������ܵ�me�\ҍc��!��7DNиƩ���@&���j~���7��Q��:���h#P9˼*����[�~��Y$]q^�Ӈ�) m`P�"1�ɒ�����KI4���W-'_������y�b/yS�S�0���3��с�M~;&�gV�NQJ�T��/�4����eI�Q���"��c�{�ǯ��R�bڪAx���q������1G/�Օ�S�}�b�[��Jvdn�"�a�AtW���}�>�:�\\�D����y���/,����:�&B#D�1
�۹Op� ��[<O��X������ι�sk����<��˧�@K�3����Aν��ng!w�qӌ'�������MW��.4߽��{�+~�J�EB�a�6%`�J�E�,�:�>Z�$�(p�@m8�P/�)�b�����0�p-p/�u� �0��B)XIi���8�}�}w�JF&�t���g�Ev�vpRR�CE�0���}_��-:nܼf��#�'���i��mh�\hK�] h��_��d�n/��O^|勿v����>���ʍ�i��b&�<��Ԡ�P�@#.� i�Ra�sLA��ϨM��R��J��G�-�tc?�hS%㊖%Nth�$t�#���09���`:D��Y�a�w✣��c�P�z�5;4e:J�~|֖,�A�.��	r<�����:�e;�˿~���T"5��{҇0V��bIjKy���߭����~-�:���/���q� �����;b��B���b_����m�ב��E�8b��!5#�*|�Gd�R!*�ɷ��^g1J���6H?�z��'�Q��:)V�5P��s�!�(2F�$�_ɱ\&��Ez�NZ�����xd�����A#�]�7]��O�*��a(~��T����q��2U& %	�:�X���9M�z����S8�R����՟�h�]��z�E�y�|��ds��]�4�r���DL^l�l$�P����fD�Z�!��t��>~�Y�Ņ�W��s}/�s^��� @ܽ����zV0�fffH.<������]ǿF�����,\����Y�=�\��*�%(�Ib© ~�G�C��3���KopQ�`����?��zf2��r����;�h�y����S�Ϋ���<�b���iճ�])�5�Y|���B�v��f��-U��3[�;眙���X���̩�%�Fm=nI덯l�n��0�`����Ku�����RW)�>�8��s�c�˵�8��Z�ͯ��`GP�ʤ�����(��P��(�ɲ���,N|��x*�]m�M��1&t;2&��,�DS=g/X��w
�7��ը4�Kp���r��<P&�ҠX.*��0�ܖ�B�ן��:�������-�����1X�%�l9W	�u����%|���g\7����,����Q�f������y|+<g��,؆Η�^`�9��/3?�#�|�y��,|�� �t2#/Y���[p��`"z�V�����ܐ_�<�:xe�Ef�~��?�Ȧ��:���$���te3�S���]�{�g��P(�Q��A��n� ��A�4X����u+#�,a��#�q��yl��g@l1c\����$:4A�q�f�Z��i�wd�`��灊�{���;|fX7E�e�$�a�{@���vPg��3g��2��i�=o9%u�+2A�T㭠�g��;�:$�69����q�`��.L?p�x��o��k�1��@(?�z?5S����I�Z#I��,Xl���?�w;��T`���m�aנ�v�\��o��F�b"�&|��~�Eo�~R[k�tr߷�G=δ�(�����ч�������8�]������V]�uU���rJ���fv��� ��Z�ŏ�;3sKͳ�:t�+G��X�/iLi����R�o�D(5��1.��D��W(�+��S�<`n&.����l�HC���0ש�	<�%���9`��˃t�2�{��j�ԁ���n�"$Z��8��RX�-����ZG���A )��8��g2(`��db��X�<�V^{<Lވ�%+�А��U��(�P7MCŧۼ�������_Y��M�HD�s}�y
W!�$aa�[�f���K2���¸�|15��F�b)�Ѱ���G�,T
�s7Y��e 4��$����#����H��΃8�4�����U/�9�h,Ph��9�9q�ƽ0����tb-k�2�������=�����f���B��j�D��60�N�lH�7Jki�E$Ƚ���u��*����1nG�|1�_*�g!9���{���Һ�f\���p���S�~x���6ћZ�
*�O���,�0+c�ԩ3�&�«��v�� }ɵ}y/�=ʍ��K?G�� ��.����SQ��]{1�+�5D_n+2��i ��6�r�e��%�n~c+��'�4k�˦����A��Sryy��rkQCe!y�q�֬d!T������%��}�%����&�g-&:�:j�f�69Ɩ'u)��*���}��(='!�m�=�����A��q:��Z�� \�=13"�a~��`�5Vl�&k�[���`�W߼���/<�.���"АgJ�~���/d<0�Lɼ]��j/I�9�M�ABڙaC��2Rm��ME�U.�)qN�-�YG_���F���J@�_��I�Ô�򠸾}��a���<��mk����ϳ�hϛ|0h[�Rk�$&�B��+�c�Z!���7�9�[5	-�X�I�M��ETj��S�$i���ah��ٵ���b��So��Ru��Kٗ_Ƕ���.(��E�����;1v��Vˠ�u���ڿ�������y�A{�t���Q��P�k�����Oő�eD�~��~������w��4��G�~*�C���Xs�P�w	i�2�"���f}�6�5\V��(c�s.n]�;� ot�Zm3��=QS���<L5�5hR�xAq�ן��R=�Ԅ"�5l�������6˰�bwn~ϊ�dv��R�Ѝh]Q�ڒ�@�	?�6��8v��8�L����|�S�l��gl�ͫ�J����!�������7k�.�JB�.���\Y��dNt�L4��uݨ5G����㔵:��S���D�׸(�˅nr?��`�i|������97�Qkܲ�:��3�K'6�5o���3Y�vb�V���l��8]V�S��~�����0��\���v�*b�̩X8�_�c^�l��[��oik��FpN�����rT�>��տï3�����\{��$��ؘr-�����o������QO/��;��('I�e���L�O������֗�W�j�md݄]{2��:g�x6���?*���g[��\{�0�驶=�6��\�Ne����̣���l��GGUXZo�7��fY��Is?"��D��^4���=矿����']�m_����sp�mT��m���J%E�I�$�*便�%�8fk����|X�dM�~��q3h�k	��_������=]N���t��R��#qǂD�����s��P� �����EMC�	�����
jL&��odA�/��{��D��F	��5k% 9]N�g������),�@s�C 现@��>��x����nW����L�l�Ȋ��nשV�u'�����S �D���X���r��.��WA&�;vK� A�<x0����{h)��o�r�2!7I9���@�)�*�<U<���yE%�ڊN���t9]~�%�V��y�ُ�\*\V��zU����Gw2��f\~]"�гa"�Xt������u�]7��n�i�[�bF���t9]N��h0E�x�ή]����?�������v�9�(7Ѐ���r�#�3��]���i��_v����_;7�p�x���}�? /xQ� ����tyN�gۉ��.�W�-Ä�,�Gfgg��x�{��}����.�H�{6����1�h��5P'���_���<��?M)�&��
��%���r��.��
w��lV��$I�AP���P�5@ܫ�N�R�8��j=�~=.^��m���G�L�⺓��P������>xٻ���c����O}�S�={�|s�پ+ᵰc�32�Ȣw)x�c�Q|)��6�$�CX"�*���*���:eq�b�`�/Ѝj�Ƴ�v��R��5��x�������#k��ߵ�<�B�	�O������q@SW�X�H�q܌�T��t���ao�ﭼ���al/�yZ*�Ѣj���H� ;| ;E���:E�	��xG�\��{��^8�4�}������|�OB'�FQ|�Ȳ>7�ƻ�!ib0L�/6��*�5�zqP�Ͼ��%�8!6"�v3�}hэ*՛����`c����q#����|���덀}i!�gq�]o#�N��}�Rp�������v���8�E�?I⾙��.��V�!q�yR���)C⎙i8w� wdB���7��뮻��p��t��9���� ��gO$e_���lX	p�D�B�H��<��k^����������Ї>�۷�k����G�-�+�T���t������Sz�c坴����ěX�c_X����^�����F����z���n
	އ?��F�W$��7	�����a�1֌=�#^��7��Nt0����e뙀�x.H���Il��h�oE�kT��T*znXw:<�� ���g���f�{�%��ŧ7�AYk�#�J�u麾�d�`�e�91�~X*u3��"����6\fYi.}����u�� ��Hlf͍�.�6]�4粀x���'����o��믿��������Ç�����Ý�2{���E�zmU�v,'��|���Z�X�66�f��F�r��� �A�w;==�4���hl����e�~jj���m]׎;h���}5�|�vj�&�+��sjsx�������%�z�_�P�G$��N9�J����n�F}k�M߀��)PL:����yek�a�xX�Z�B�=5�������׾k�9܈�?���^���V\c�^k=�:�n8�׺�XN��6�S��oI�ڨ��L�n`�R���A����):Ề�����L"�X&�I/�zF��6k6�����;��{W�ǷB.�qu�}l��O
.x� �$�E�(�>w��8eo������w���Ǯ��j��ѵ�^{�/x��?��?}�����B$��.�L�&/b5���&��'r�|�����V^0��3Ū�x!!3��;�]�{H���:��w��m+��	%��*O�i�c�;��;8+��ĥk��G�[�mx�qKl��g��(��%@E_�1�o��@�ժ�vqS�~�x Z�ӯ��K�VJVf�˳���W%i��0�{T#c`d����dy��7#�3�_�6�Ĥ��o[�4�09��QC(P:;��uy}ۛ�t�~H�Ի�I��`ԏlk�*]/o��z=�1C+��^���U��=��O�����q��K
A���'�u��7�BԽ��"��e�&��	�٨X=�^�%q����/>��?�?�o��ozӛbt���4��c�]�$�����OUWW���43 f����K��?��b mXA��!����^;�4�#�0�:�v��CY�wm2��l�+�2)ٴesVZR�#һ�\`�`�3�ӟ��|�{_f�򽬮�|��
�]Y��2����=��o�X_�|��n�ʉg�=������+Wزڲ�;��+K����?���
[��~b���ߵ����/~����쏂�{f�U49(�cs�1�v�]���ğ*�,(Y  ��^��ܧ>���~�����~����ɑ�H4�XcKa�P�U������S��?O��q�r<��U�y�f^��P���KOׄe����(��翑��O�ğ��������˗/㋚Nc�5vRM\�tI<��#ɯ�گ�8��$Ap�0��1�B_2��%�9��<�}��gkP𫫫*�:���`"Z��Ye��;�x�1�O�9ئ1�O~�w~�y���p�������?��}��� ���=޼�n�n� Km��}�wy���Ǝ�N�Ō�F�ʯ��ʵkۧ���/��{��{6>��y� C�4���l0���q�'>�P��)��������
0�&�{���q9���x�p�����[��ex\SJ��}��Ȱ���2�6-)�Y)���y����V��s;+�)���1~�&S��rn��0�;�QM5Ƨ����0Ƕ��g��粄��yѻ{�|�t�ó��V���Ső�?�G��-�/�P�11�nwM^�~|�֚��0���\�L�+�?��v){���N��'�|r&���7/;H��+2������j��w���I���Ղ�w1����S9�)  �wȘy�w���o�fn�<��u^G��eQ̻=w��m���3��͹sX�s��m�\�����v?a�޸��v�����KW�b �tU��@ ���x1���.��~����ذ/^|^�{ �[�6���-��M,���s:a1h�#��G�ۧ����WVʠ��Nڻ�P�v�w�-�������N>,{�����ϟ`�c�$ݹ�c(�'�����#��1����[p�o�c�0Ǜ'6fΜ9��:8��c�&xZN�ܾ�Y͹?�!>�����ϳۮ����nz}�������v����ޟyu6�p�0|"%w�@�z>�>��fY2������I��n�������|�3v�۲�7Z+�?0�<���z{�����Fǥ�1y��a�� v�v�=��x��y�N���]����v��6�W��C�%`�эY-���(��(qr�]w������n�~�ӟ��[��[�06���ի����r�O�����H�O�I���&�;�n���6=�;m�z��_ߝ�;��}��;m��ENHp���{>�x:{�y�-E
Q���{�e/^�[]]��s����O}�S��!^c?�я^��������si�>t�ԩ.x�)����>��nĻ B_��{|����k�̺n��_7O]�pL0y�`B�M��L�[�@3��p,���?Ը=s�h�x�iF����?��̾|��Y��O^ӻ�����ޖ�ox�R;���S�<�pd)"��?^�}��/����/��/���/�⡏u(Al�3ǵ���?R|o���̲�n��=�rP��i���{�[{��IF�C)�-�s&0�V�u	 ����Ё�#i�� Sf�b\�����ȭ�/J����q"x^��Z��a�r����FpA�398:���q,�����/R�T^$�r&�$ڠ���7S
/�@��AI5)-ɵ���u_�B��]��IT�.Ǐӡ�,öx�(�KVVYv�?�wHW�������m�Jqq��s?�3�pߴB�����E�0�I,����q"������s�����=Q�ñG,����kc^c��Gx��螖�GZ�h�����x��q|o'���}V˽���۔���X��)/c.\ �cR����{����eߵk���,�H����8�}��ۨ����Xeekcw�ʥ!~�DJX_Ծv�����_��@',�e��~/4�s�U~�]M"B�H�{�s�A� t����=�Q���R��>j^���}�>�N��-Hd�F�yt�xЬdX�h��m����%O8֭tpR��U ���&%w���0����O� pǉ1Y鱷��39�߀��َ� 0ւc�z��_������J3h2�s�=ʌ�g�e���h��l��b|z��"��l��^�����,���p��C������6�<\�xc�;�_�������˿���_����d�W�^=��~��>�8O����b�<�ϸF
|Q�w���,p��ˊ�� �$����2�%�`��*��E0��!P�0��z�ILhM���£Վ�`�G���fK�(c�<�L�!Q��~�h��Kc@�|@XC@/��E;�o%�������+(@�8'��N��u$r�Gm��2�h �)qr�5���0E�m;�K9�S¤���h�=� *�f������Za{Ĕp�J�����ɀ�-\XMJ����� VG=3dD�=�rV���Iø	���br������X=.�5N���ۄ���Mx�1��ϭhғ��g�e��[5
�MFJ@:�w�N������R�l�2�AJ%�( ��w�ԩS���	V��	���s�����C�ffm��/��� @���ׯ��~5w��n�������eٮ꽾�{���d	�y^=R��hx[[q���=&S��q�x�����e��"��K�ӝsr&1R����9�+�qE�?U�T.�P��F�ǅ ��b����'����ϸ�z����!�"�����]�L���SO��s&a|�G�R����5��:<�����IT�� �Xm���pŢ(����}���F;w�n�d|�
nDD�=NJ0y�}V^B+�\9pO|3��E�,'������d�����;������]-���z�\�� ,s�\��:��{�to
�r���'�]�z7�$�L6n)�w!A`���r�� �> �+�y��������.6M:��x4���~� �|��_ޅ�a�׻ ��f�����c΢w��S�a�;���a��w�n�hg���~�9`��'�.�n��<��\��_����C�y���Ƀ�S��Ws0�3.�A(��Z,��#
��ܧkk��/I)�s�WP `�t��=���Sq��RIъDǱ���G�g�A݁\��gE�&e1���Lc��Ȧ�i���0d��bhY���"��^�F8��\ܵ����M"�)rr�i"���y��9Z�{��vZ��or%Ϝ^�;O�,��k�h8�|����P�`�9�1LpH�ޑm8Y��@$py�&E�%3p�a8y���߸y�W�+p~m��A'�<m��t;n�&���s��"�9�j�d��p�̞q$-��b���qG�<����ʸ	BªG�F�����6��c�(+�$����Mn"XY�����e�oR���l5�[��-7��?<v����Y]]}p���a�7�;����ٟ}��qd;����;�������>_��_������)��{���9jeU0m�17�h���� �Q��I�|;Y�NH�O�&ar�Q��N��׸����>�K�v�]�~ྏƉz��J x;0!�g(`^���׿�ҿܾ������I��(р���̙���s��璟��iD+ ���ko|�ׯ�x���GW�l�ٕ�`�׺�����<���q��\�p.�E N�w_��֕W߸��¶�}m��$3C��"V�>���=�6>�鬜�/�OH�~0�x�[_�z��w�\��=0iz7�Ol��[++�^���VZ�48�q᪣�s��7�n�}�?۽��؈k��u﹍G/^<���Xl��� ��0���b���u�O�|���`��^�E���@e�k���>���/~$��ݭ4��$d�=�o_y���|�]��m�l-�=�B�k�����d��w��8γ>k�6���zk��+�}�����x���������Az�=g>t�}g��G�T+�iFD�h+������o����n�<Z�����7o�<�}��Y����4���vwwEm�9,�]�!���Taw���t'��8���3�9��!�s��K�-k}}[���o����օv^z�=���\�:;2���aNB�&| ^�|����ÿ���ܹs����"<*����x�_��k�GI��o��a���v�_}��������om}������{��+=|�#�l?Ny����dC������G��}�<��W�����w���ߕ+��������G?��յ�@���%6��2����~�ŷ.?���b�]X@���:{���Ӻ{C�?�������i�HH8����㯼���޽����?���o~�K����_�>�����<����W�m!bjG����9�������{�٣�~���sK��Λo����[����?�m����V&�ܼ��֗���7�����փ���v��M��y�ů��<|���m����@�[+��������_�������ȟ�䭻�ڴ4Tx���������>���ܷ���oL{���P�����~�+�����?�ۆqb{>8!�W��Oc��~�#��hue�J`��Ip�̗������׾����я���n����.]ߗ��'I�����Ǿ�K�Zm��jJ
����ܸ~��W����9{��ޭ<�_��7����~㡽���鍍?zࡇ�����O��O�>K���k׮�gri����Ⱦ��/Pg��￟�.]�h�3�<�e�Ǝ��*v��Ǝ�~������o1�D��\=}�?�#7p���;Ϟz��Ir��˭I`M?�7��6׺�k���k7>󙟚J���/�D�{������� o26R�$Nٰ��R����Ц$����L���_���C�=�����7uaoC�����:c�_zS���'�ݩ���g�=���w�����X�Vn4� �#�*�~��G�w����z�S{��}�s���#�'�gm�ӎڰ�p���n�Hl��ɟ�k�'���_�k�G8=������� [�x�+������፿��r{r�����h������^[��4�O�g��tW�����������OMi�|�s��_�w�_9��P&2'�+ˈ�"�6�	�y�S���/��_M�{S������&Ġ�į`+��r}m��v>��W���3�O�����ށ��-�N�����}����t�t{{�`z�CL��u?�-���,���m1l���4M�N�3
H�s�t0-��Y���@J�	k����w���~���3�٩c��?�X�v��~�(��EǤdG��sg�v�]�$>{����=g��4B�G:�����\nn�]8�(c=����}��b���0Q�i��Y+^��7V�V��*q����~\|�+��t��OI3���4��/�;&=�y����~��S?�7����O���W��nmoE0�10�y�ju�����c�����aj�Ng]��ͻ9�:p9�}ֆj���n���؅�T���	��q�,7q��tD���8�W��y�}�Uv{衇��t��������V��|6�c+��S��C��_�p�ʋ/��j�Q
����2X�'��4���Yg�#66�Md>��X\��2���4 (�3��:	�ƒ���㝅��L;��E0��>G:��2~��ߨ �=�
o��-i���5e.%5��\�Ջ7+ ��]eI*�p>qc��+�Y�?�+�N�����$��^I�B�k6����$R�5V�ۧ�$M[pi5��rQpdG��(�d����j%	�8����@lu�M,#�������#��ʿjI�s�^��Ɉ�ã��䔨L��oZv:�D�P91͍��s
���S�K��C���I�%Ȇ����k�P��9k ����-��&�9r��D4�18� ('*��R& �?��Y�c{�a���$鏕�9��J�G�^\������(���)�6N����vt��y��0
���b"b6 L��p���iv���\P:w m���Ա5Q�X�Z�o}5֑H3f��hmy��)$	����j���|��a+�/��ĕX�E �m�6�����xK�#!4ǢTa��k/���4�U*أ����k1\��6'](C�a������F�EQnw"`>�Ƽ��1���?���i+u�=�١����/{�J���@ }��Z�=�ֲYpVGA�c�������''Ef����e��U���`B1��*섃шH�R7�ֆ6��P�[�U���%�y��5T�䊢`��Hs�����["�[$eJ*s� �*A���(�a}��$��z<F�r
FZec��� �;�o��P��U�b=�!I�u\��cX�n��EU3k�T��m�(e�Q�����h<�%��O��\�� ��c��i��0�!H�<�B8�I���}l�E�q�+��-�"b�XZWT�Ӫk���u+��%ƚ-��J�u+;yKsҲ!��p]����(4i�Z�xl��r)��4n�UY�	&-n������ڿ��p��c�-'-9- �_��X�j�c���ص��i����A	����+v�"Y�b�26g�����J+�΍�q�F�K`��`����X���^�8���mo�X��)��иprNL+pл�i|Kg�g��0��ib ��}ӧ���nF��Z����x��K��+��Ʉw��Xw��JM�Mb��"l���̑�d�h
y����W�T�r]��U3x�x}X=�DۨZ
���{���,��iR2�dsx2H9������pU����z+d�bP�w0ض����y�;;&����dF7��`�;\Հ��X�'ؐE��A�;ǲ�	����S]@�"�k L0B�9
����V��y��XjaLF�p�К�I�#�>�F���y����1�hq� �*�����1aI2P�N�+'���?�Vj�E�fȢ��=�A6M C���,'־}n��D9\V���p*�qR�:���}EdH��/TVEF�0��5X*|��]��
.�;!1L�ʜ��_�&oil_h�7Q!�Ʃr�O�0���,��}XG�2�����?�$)���(�}��p��}Y�
��^��y��O!���8o ��ʯ96FA+��p�#������ᒏT�N(eAMn} /o�ܴHD�	&�<qQii����x�K��e��;]4z�� #�=�+�9N#�1�a�r�!R����ÉOZ�ZgE��s��Ƀ߮�v��j���	����4d�ː������}�ؿ"��Fo?.�7e(J�ۣ�,Ƀ���NXcKa��`���D�W:�	͋��)�\���� �I��b0,!� ����e�4�^x�Fl8T���c/�
��(�� E�F�<2�y�8쏡T	�*3�h�F-@dJ��"y� �1��ϕt�6�`�$�`�,%,-���{�������{��U_	I��I�5�Q�E�[,h9ji&��I6#Q6iQ!!�8��vy�����u��b��yS��%Zk���k\!O	�:�	#�1�"J��j��ϩ��(�^�ʞ9�f�K`��pCm�sxLҵDb8xu�OjM.�T:k#b�M3�HUHE�_�GQ�8IH3�jN��p�di+Aa�Y�p��WJ�2"tZ!�Wml)�K�X<j��r��4����vΟ�;��`|f�1#��n�"0�1&�e�M��K�2q6K�����E�,n��n����|��=�"�\*�+(�$o�UƉTQ�Ɩ��?�F�- Ѵhk�WM�ɋC&5+t���7�=����d�\y`�
��Fړ۠$�18�B�|z�Vp��;��z�!�g�@FV�b�R��HQԚ�� �\��vQǾqK(����oظq��(��j2�/'�qx��ޗ��?��1#��O�&�K6�"��������g���f���'Ym�(uL��CO�� ������%	v�����PD">���D�we[b�øJ#�θ{�
*n�(1��Z_�@�Qhk��Yx���[��%wt���/���������� �I��D4�t�q�	�7	l�y��^�hH���c�ZIO��_�&-��f-�4�]����R�������q��O2�vQ)�pނ&7�xr&�A.r?���7&��/N���\��d� �	7�5��uNpk�����`|@��	�ցU��,��G�OdJ��v6+ȃޤp=��Ű��sZ���1�8�0C��Ҫ�����Z'�U$#g׌���̜R��R�eq�N���:������=2��?����͵�(81�?��Xc'��?�F�?�8��Z)�x|�$e�S�`dL�]��M�����;�ܠ��T�,��(Q:��9��cyg7���c�8�2�k0�ON�8k�
k�ݦ��&�~O�k�7wz��G��7_��l"��o��p�P��"�OoI9����(�,�D]Ч�نx��GݡG�����ʰ^f]c�Y(�0����Ź\�W�R�!��	ܢR&S�s�x���sv� Hx��9ֱf�����o{Y!\���on���nlD�����s�Yk ���-��2u��I1�iS!~�Բ�`��Q[7L�aRSFIz���K��ދ�;>IY�4�(��//�/;EO\�G-^�U�D:�pU�eo�r@8n��dU<&P].����k!�Jc󷶪B�!�cw/��f��)x7�V}tw/#*�pyq��[5K��q�w��B6*���^.�������E2��qMO[k ~�K�KЏÅ����Tg<�9�R�ӮX�oJ�I��y�A�A$|����yeo��BhLERf�P��ST�d���'J)�f��s�w66x2�%�p�n��7vr���n�;,�]hYnx�YM ����M�ڪV��{F�%=���E��q��cA��E�M�t��f�G߯:Y�w �]�ޞe�qZf��fB!�NM���Q��o�^ށ�uokc'��?�f�(0Ec}�s>��͘��-�!��c/T���F�y(�����$kllRHV�ɥQ��5n���x��{�H�9)T�L�e�}#w�E�9c�uN�vymc��Xd�WDotx�����R�1&i��t�
��{K*����ϳ�N�5 ��u� �����*(k\=�
c����}����E=�F����}4�8��Q1���$�T���'�-x����ac��O���؈J�~��1�wY����M��E[���*�*�\�ʄ���ܙ})^�&!7�.�ݾ���JptK7~I��nDi	2þ��j	��X>���K���U�*���X%f�y�@uZ5�d�7Y��c�(�@��~>'�al���
júh���%$�?���)�2�M!gGR�����/M;�(�D5��4<�e��O���n%Q��C/�������";
fb�I_�p�)1]�򅆅r�$f����q���r��`_��4����?7�S /f�f��)��%��O�I��G�f�vG��p���6��eG���������jǧ/p
���^���&b�{��I
g7
�����S�~�}<<4IҢ�L����M��`�+)�]�	��t�u��e���1ʣ�$�z����O�I��J�VoFʼd�.B�b�=tL��,▓w�w�]~{�7�!���æy���gt+�)Z���Y�$7\�/ F�Z�!QiP��Z lM�ǳv���[�#8�"�v�iG��i�w��0�o����� #�Fwx9��H=�f�Q��M��ډA��� ���?��W;��g%��X��^�j�4�^�������uZ4��g7����Z4;�Y��M�sO���&�*sJ/|�@\���?��@m��8�ts
��,Q�q�9xI�~���T�I��6V0a��$�6nΏ!BB̞�8�^0��+|�>ˎg�Ɩ��?�&����� g�xr�@�[V�X�t��G��G���w��c{̲��/�>�<jф�^�9��^�Q����?w�z��Vfm���4�&~�UZ&��9�]��������"�lǆ��i�� W�TA��*�5�fy�ƍ�I�� �	7ɂE�T�N�=x�}�bG�*�`B�
ۺ|�2�t*�N1�	U2�x�>|;V�\ؚ]�5O�m���=)�
�Вhdu�-�I0V���X���*M�x��a�X���a���|���ע븸�o���R���Y�'�J0~<Z���>" 2���[ t1���cR��+��y$W�,(���9�U�h�'6m=^>��fGp�1V-�.%�����a�f���}�fYU�<x���ǹH&m����/��/H�߱�����O�	)���UZ�\�9��
�����wW�gi:���le7@�P^��͘%V,�&Y�i��[pƌT2�v��M�k�BVL�Ċ/N{A
i�BW{{�X���a>kDh���_*����#$�nF)ga��v��qa��ڎ��{f�)���p��)�͡s"G,��$��l80�ذ$IX>���u��h8�i�r��?���-_�gui�'�u��ƃ_"k ~i��~Z��8���c���WW�<�F'i�f�����g�EіTkb��z
[ŭ�� ���ߐl��0�
�����Bc��ڲe|���7 �$� �	7��S�AT��΀|Ѱ�p�jB-K
���2v,���l���S��� /��_�g+&��n���me"&]�>#�;�c>�U�(E�Z�����)
 Dy�sl�4�T�I�Y&��p�F.���˓�Ȏ
/x��GxJh�$'�]Eք����o�g��R��0��Ӣ�.[<�=���6�-�(DÙ��d���*�e�*�'�<��^po�U��� 㠚��qb��[�Vi�,^��N����(y��ޛ� ��q�X�^�Z0���Wخ �Y=�{�F�X0���}%̪����U���X�[4	���ϓ�~Z��l�+n�@)}1x{:�v�)<S�a�Ež;F,�c���N
w��<x:�1��{oY�Kb�oۗ�<�k��
����Q��E#+��a��w��aj�vǃV�b+=2�f���p���L�~�a�����������X�'ܤx{��2	U:qM��P�|�����í(�|R�ѩ�^��VC����G�H��p�T��+i���x��D4jKc�7v��>��G�8�ad�D�%�q�Q�"�yz��em��(� ���z�w��<��H*g*?�B��������]�ػ��_b��/<e-��WY4���/D�$�e��z;16RM�2�9���|����
Xx��C��\X�+��R�a�NWG6�1�@X4��و�b&'�95 �l� ��2�-?�����a[W�|?WMڲ'ka[˗dE�꜐��j��W����z�)s����ǽL-�4lu�+P��M��e��O�Q�#+XUU�6tI���@!Q.��\���&d�S��ǻ8uy)��Ul��E�-"�FC9/a��LQ줋 ���a�p͑1�{債>�T���\�Ȉ�6w"����t����n��Ԏ�oȍ�IKm~6�Y��A`'~4fǔ�)<�rC��-����S�)f�-�5 ��B&�/
�Ȩ��ӻ��9�9Mj����g�$k;^Ӓo9jQ�/�Xs1I��c����崊Ŷ��JV���"� _�N��`��:Q�4��ll���%���:�ᇥ�Q�fɽ��Ib�;��te�S.�M����c�x!�&Y�k��^���V��ES7xQ/(4ԘOq[���l��/���Y�KbU�?�2]�n�_��c.<��e=y!����4�8�a����Љ��h�c���9��{a�8��I��׆�Kj�(t�G�tXÆj���
�W]�8&�1���s�axI�����?�&�����p��}��e1Dc��)�I��c��#�;~�Q�p�S�����F�*7C�y�y�
�ЩH^����$��$�EVp9�\���G�(ÐYq_^Y]�l/��Zm=Ac'��?�f'<�(��_n��G���Q�Q&�!2�dvc���4G.�R�&�[ܘ]T��!�fx�z]�w^�V��*��(f�;���X���{��x���j5�*l�Fl~uj�}�g�T���;�� ��)�b]|s]0�FR�<�	J�&��W��:B�ҟ,��+qzM��-���K�"]�*��P�ɪ��x�ȼDG�XN�x_ʦ�M!��X��j�{	5ۃ�&::�ԯ1,��b��uDC�&6m��vV�h���7c����,*i_�s���J���*Y��I����k�����:M;|��&��� �I��㉽MrBC4�(���j���ݨ d)L�NUFc"�v�n�H��~KZ�nBV:��[�e�;��2=�`r�,�/�����Q2E�h�جۣ&is�t1S�NL�f����*Ģq\{��G��Ф����֣bV|m�77vr��%0CMT�w����#�g *�&��4���Ӌ��0�E��r�r �T
�O� �
A���(p���0�<޽%�^kW����`���sb��{�a6vN��a�Tl���B�Y�z�\嬱�����,�`�Ԛ�=d��uV�X,c���s��}�B�N^�A�`�Lfg
~J����lA���ã��<xn���LT���
����~��J.�1��E�7\=vA\�{'	�1�4g;je�{{Y��n���W˸ ���샧tr�â�#6�����hd��]x?���˞���E �&���%u���˞��ͤ��!�Ҿ�E�]���㩅���G��38�9F�"o�|�Śwz	�	�2���Q5�����s��dMx�J�O}^�>��K�jձ1�i�)�k�'�t�F�-����MZ�-\���N�"k����6$�0��cє|9��(t4���Y�b���7��h���_b�k�vX~�"C&����y��'T��&,O;[�
�췔��y8h�t�S`TϢ��k�E���?�K�V�	���s���g�^Ǵ��8�;sK��l���M�Yv3y��()����X��y�1��+��!�0S٥K_\B�`��w�r��A$n���&��8�`˾��YFfYUg9�XI#T�Yc���q����m�����c�`���j2z��y������o��+��l=R��>��X?SJ@�rΟ]AGs_�c�`�+�E��n�,Ii��� �&Lg�G�đ�&�k�Hkgj,���@;U��qݏȃ�^hl��\"���E��&<^Q��:��v�̛ocW���)k ���H�  �Z:j���D���J�K�0ɊTI�5S�M7<��Y��	�R7��܁�0��#��#&(�s7������h�د����d�z��xF�'Y�IV>Z`������ܙp&�v�8�Q0}V^)���PLQh��J���6atG���s06Sl����?F�7v���e�"�&t}�]�T�I��d9�S�ג~��._~���3���<��Ǣ��Bv%� TUe����u����
��2o˾�Ի��16��
����S����I�YY�Zl�ӕ��d����y�.D#�ͲX�K`�-V�t���Q%+�ڊ(�<�˾Xy��ֆH�ݚ1���Ym�a��i��RA�:=����3����B/n�YmWc�V0�������v��m�'D���X���7y��|9Xn̨�Sc�c�7�0bL�W4x���1�@�de�y<xX`ĭN�Es�sJwV{G�[L��v�����A��j���]��A^b�����m�h�gÐ������ӔI3�h>˶أ8�#��4�޵�X�;c�9i�ПXw3�t�� ����>�*��H�?�
Q���Tc���<�r��Q�[�����������4�8M�Z5I?�t���$k_JޤJ�Ƒ_k ����H�bC" ���_�a��̑�Wݯo�8"ˤh���X�	�S�W�Y4����s�L_�>���w��cֵ�H R����m�p�δoI��7c���� |c>"�>׷�1�P)~�˩Z���Ld�ԝ��5�Q�&��U��p��>�`�0 b*Ի�X4�@�w>D,{���G�{���=��D�?;�de"o~i��%5W���W,��9&D]�>g$���4l���E3w<�EM���ix�"�^�:8�Y�J(i�E�'G�P�6�8J���fE�&ML�z��*`�o��q�|-�h�m�Z6�^����f+U+Ր�(:v	��%R`�&�7��Z4���Ȏ`C��2�G9�T��J򝂥 ���5�x��*ש��D#\����B4��bo{��22pKhN��@�3���!�$�b�UCu����4� |c>�Ƌe�-��#�:�撇EC6�����ǏS��[@/���Up��tjx��M;^[�V������f^9!� ��wMl�Z[��:<klI��%0���n�5�h���˹ oQ��4ʘ�E#�6g5<x8P�{�X4̶�4vR�r0i��|���@�ۄ`Sp�f5�"�d=��{���7Sj��01��|�m���+�8C�l���rX�'�Jdǉ;�r�\b$EkQ�G���-U��b�K�Q�$-f#�1V����a��h+���M�,d���&_�>��Lu��)w�Z}ӖʓM�uy��%5ˎ�3��'�H�)c�������Q΋��3��.̂�qc��z�w"D��ˬ���&Z��Zz���7�4� ���r∋�	~�d%6u��ܣ�/� >���~W�������͑h!�<6��H	��$�I�����jR�Nѷ�(���Ȗ	�&�<� �	���%��qJ�(U���˛��
��M�c��h.XF�S3/�c�;��GqI��$�}@6���B������-� }0��s�p_&k ~	�P�N'�::���+$�V	,���V幺ti+t^���"Ģ,���K�V���!A��/m�b��<��!���-w)Z�ڒ�Ω�K�V�s�m���4�X�K`��U�0F3��7�aj��H��J4#\�E���Ң��р�,�iWp��m^$g��lE]�\�L��%ʃ�ȹ��ab���@ei0|��\rT�;->�±R1�#ܛ��Q��N��z�V��9ϒ�/�n��s�	A���4]�����5<���O��� Yķ�yG?%
����5�$�c��&I�Y���?x�F�������b;��0��<� 7��,OD]\��Y�*W��V�Rw�E3=B(U�T�ƤlT�<��TV�ƈ�?�}�!�B�Y4�9�Mv��yD��&B�\� �	7��
T;���Lĭ2�ʳ\'��&�P�8}�L-�l��D���E���:4�e����my��+6f�B������d0�S��i�BL��-'��'緻�9v5�eI�4=Y���_��>����Z-�b�f�;�?a���ь�c�p��(�uv�1/ˬ����hX`�t1��g�xN(� :�q�6��Րƚg�͇9˕*�9���X��`���<�)S'�52��3v1j!�ڇ�c�X�R�a��m����:5n�Ft{�縦�6k�8�����"!�Y��\��B[������p2ċ7���U�<r1�8I80
�Pa���Ao�X���-�%�y����*c�Q�Yn��/T�-<��������3��*��p9��?4"j��">Ը#�#���&���Q��3E�[�X44x�WLD��ǆ��,q�4jܛ$�X�Kj��|q�`��Y����w�]���|@�x�^�p��V �<��@�4ِ{p8����u
�.��aS'�����z�d�2���[�<��Q�u?l�E������D^��H��{����d5y��h%�����[��U�όX-�d�C��+|wvkgGֳh�x�Ģa7�$x�F1�N����I�#�4����Mi��^�����d�q�dݧ0��}j���ϳ�N�5 ���3�{�Q��B�H.xe���z,iwDG-���6 8�s����o)�h�������+���pE���' �p<��ON6���E��;�d<�dь���Um���X�9��d}���s�=�;�� |c��m␳j�+<88���p����hd�^[�ʽ1x�x\'U��	����p0�xV�̤����#
#�)[M�
q~�vIuZ4��C��8}1xw?l�8��z�g`r}�G�'ݐ���_I�����J8�h��I;5�8M 8�ξq�㸭���&��R��	��ifJ��6���'CP�5���BgG�j�m�=oߙFYՊ���E�����fW�"n ~i����� �L����'J���|[D��yΞ~���>f�,���o�Gm��Y&�Nϻ6�ѢѰq`��&��Є&F�t��腿7uR΃�O���|A��>Fm
<{��R.lٛ�����[�Р���2a*�X"�͹���x�5�1iᤴ����ΦA|�Q4�[ѐ\0,8|�n���;��_�mN �:5�Z4�p�����X�K`~v���H��[E���Qk�f�ܲ0��_*6�K�j�p��1��qҍ���'�$��K�q>-d�p&2����?���R���3�8��cBڑ���[�S�ԤMԄh���o�l�ѳ!`��::!�ˢt#��1�i�9L,̌;�E]R���O��$�_����O�ގ�P�_A䲒�ԃ�ĉ_��`n�
���_��&��b�R0I��a����v},��&ɜv�g,���âYD�'5�<EI01&ﵪ�W�$qc_^��h�q;$�Y:�&�h��`""�˙���ߣ�3�a{�6�,���d���uw��`�\7��%��O��V��RLg)c�g
�F�"r©�GP�=tH���g�wC���I�YIϏE��/%6��ش�e��a��`s5�& �����Ӳ/33�	��c�_�U�Ou�r@��K����$�<�G?���8���t��җ����p��}s�7�H�,�5 ��m�$�Q|Wlr��3 3��w��n	����M�N�blq��eh������WZ����x��Q=xC�TC�XT4�q��?�l��n�����n��16 M�tar�}	V� M2Ҩ��{~��g�׮�����B'��~<��{B4�d�s�ʕ��vL�b\���'�=��c�G�0����&�m.�>�'z������ػ��o춬,���!9x�m�F�s+Y�g����E����ڢ�=~�C��,�ݍ	X���c�+8����b��oG��q�b�}461�e��O��q�e
���(�"_G'�V��!l�()mk�Ǡa&Y�qv��!v���V���rc��M�k
��l �z��d˅���4�f��M�Y�{�qG�wa��I�.�5 ��B&d�^j��hG����a	�:���?�9���9�s��޺\<��d�5e���{�ǜ3~��;ךa:����΋���<`y�������
���q�T�<� |c�m��&����ڧ�p䗧��̱HGK����L�Y�Q�P�~�4ݞ�������<�8V�CU���;F��K�1Ԣa��_�I�s��rX�Kj���zd!�2:��M��B��e��� L�'��i��38�`8��r�dt
�B�w<�l����,�eUc���אŅ�b���~'<xԾɔ��X2c�e<x�:7�x�o��[J���M~y��%0a=���/.U���1�5=�\b�S8 y^a[YS %ŋ�������Ֆ}��\'�T1-���#�\2R���עI|<x�c�3rq�
��C�ؔ2ݶ�}s��=fRDR���-�F���-5t_���'���$
����X�K`�Mh��MG�����D�b2�,�V ���"UPk��&_�?D3���15
��$�͡3ah��D�L�����Z4�*��w>��ػ��?�V��BY���o��\KX�,�N��%9Z$G�:]��{_5y�4�a����6*��<GW}���V�[ V^{�ă���-��~A�@*��ڷ@��B�h��a�F�
4�߁(Rc�^k �1��b�ĢqB
���,N#j��s�.o����#෗E��Sze�e<�G�ٱ��GMaUz!�Vר���_`����17QD���5���X��-n\�2DSJ�F�Z�� %�.-�Gd�Dq�N�jkmhc����=<x!��Y�{�z���w��հ���OT5����}+]�ؗ��o�k�e�`7���'�ob)�hB�������]�)�~Lt���xX�V{~���mp���?�̘ф�;*�âh�G�(<:V�˟�/}3Eɇ����ola�Y�^���D	!yw��>�hZ����:	���yTQbs`�� '���p�>욤}?h��\��z񸚐�*���9�q�kՎ���5��%���-#�5,�3��#%�/_vz��
���)��/2¶|IV
���)��ƅ��e0�xY4�K:O�ؔ��\�mą:~��Rb
Y4��:�#[�_,��.�ă�U�R�`�l(U0ۭ˱���e��������XfĦ��\�3�q>`L�X���{	 s�O�Sh�h��t���iKd�j!/_O<z����my�ƶ)F-,��<F�5'|�=eY����ȥ�޽ F"�1�c�Xu���)����4��墌�!�J�
<��g�#(����
W򻂏I�O�����X�K`�ݹ%9&X29�3W1�ؓ�ۙ���:����ۊw2�P�s�-���{�Yp���-QӅ��9<���&=xwel�s|r�=�
����2Ex�xg8��t��+���Z�$L5�����[��D~LvfO�ҥ�
�!��<(J�ʛ{�w�n>"��ɳ*�ڢ]��93�Dv��m�Q���D�2O'����~�ʑ�6��&~$G.�"ǂ���i۷<� ����aq�1/e��+�	��>W�+�G�)��U�h\�F�0@i�n3O�P\H���?<s������q��]iM��!^F<%�M����a�8��sT�����w蘜@Q��5�� �	7Y~�}_iL
����Y�I!k��eJ/��*Y�"�������-�����;����aê�;�U �?'��ԍ�
|qgS�7R�Vw/��	kB4G��d#.c�8����)���Ч��l�/�Ej��!U��+�{�rmu,��c���+L�&�%�U���?5K��4��H��TDU�b��&�!&��Xx�v��+�Ҫ<�h�~�c���� ���|�A�������f�J$� ��J�[~-�Z�σ�p{�Ig��e�c���E��b�>-L�Zl���eV�<x)��֓ZƎ��ܯ�]I� �z�ׄZfgGw��e���-C��s�O"��F����|<�����Uo�f�MP�������Z��mB���T<��v9��c�@�{$cBte���<x{��y�������M��ii���nR�����>����+����Ie��b����+8�Pe�'>zWAtַ".:R̞�SN��_��TJ�|��}e��Em������e^t��0L�F< )���)��Xw������r�{�8��3������'��/�#� �#��
�F��;�>��=b�o��Mq�Ɠ_k ���L��7��Q��8aA����$q�~la���h�FE���}�*���	6̌Q����4Ib�p+	I�xY4�f�:]CJ��a�:�$��S��	S6��d� ���|�,�-�6� ���)ɚ�����\g�e�o�Y��I���3�s��X4�������Mwޱ�G��cF��/%q܃=Y�.�P���� =�x;���U���c�ώ��x���`a�;{�%�{���%��Dj��D0͑������gElh� �:�re�S�h�'DS&E��Q{I.��	�&$�����(�+U��ĺ��������=bcX��*�-�%O��U�o��*#�ES�Ӡ�vaSk<�����Z��x]��6�����I�C����]�<��y���'k��Zp1
2���-���dѐF��/�X46T��4�5����)��k.�HcO�m��m8E���p�)%���ƍ'~	��Ƽ��5�z�QG��� D�'����Ƀ���~��Yvc�R(���N���5�ˠǊӃ���#h��>��f�����
�m��g�q��:�҃/�SM˾��O�U�|���<|���F����Q�����]��xi�`��ictl�i[r\��7�ÐP�ok9��;=��L$��'=��<�/�5 �-��.Eک�Ҩ��Q ��?賨ݲ���ixV� d����al��$V��t&�-����V9�ܦ><�h�'��~�����z�hʽ��rR9w�0!����+m�Ɩ��?�,���|������{�hȤI�*�
���F��Y�VU���os����6�h:Fq��H��Bf�q1M=[���㐎fEW�Wr��)�x,��� _iCqv�H����=Y97U�pM�r�;�����Cd�k�&"q�0�)�S��B/�B�Ɩ��ol!�j͖P%pRC�K��V�e��LOz��߆���D�>HƯ�L��#��D�J]n^�3�)iI�\�l\m�'�
�Ca�`渜t�1���N�T��^����T��x�-�(/P5>=~Aɦ�u٬�%1Si�4#i5c�nOR$�f�!�2��h�7:<�7��l�Ӣ��n�(>_2@��6!7�r�m�_c����<r�9s��>θ%:�߃�F*��V�79[y͍ɷ�*��������>3�J�Ɩ��_#L���)mk�{�T΅!v�~>-�������g��b�nCVg��qeՠu�Ç��Za�1xǢa�΢7]���H�wɢy��Ż7lÃ_>k ~)��{�3.S�ҩJ��>���j�%z�q�(��N��~R'A�,�BVK(_q��e���a�����s1��g�`n"nIo�j�:�$��hj ~٬������6b��:0��p	������lu?˂�4����6�1h^�mG	T��\Afc��/Z��b��G��3�a붳���$�ͲY�'�j3��� ?�4)� ��>��){�J��B4[�s�~>�1�����ɋ��{������x����j�L����»`�@�o�m4jD���y�����7m0�؉����!~���E��t-�Q]y�Ϣ��g!�iw#ɵ�fW�hdMX���*�-T��{���BH��2Ë[���ȃo/�g�\�2����/�5 ��J#�[N�A���PJ;�Eإ�P�u�.����i�r��Xý�ϗ�o+��b\_+���y�rZj��w�D0��s�ny�	�f0p:�{b�rK���*�ds�x�UŤ(��H���q��m���ӫg�Юw���C��;�G�֦�uI��n��#ĝ���}����+=���rb 7�Ï�!��Ł��>����M��~�A�c�\5��]�1x��p�% �$%�g���FX6Jx�WW�J8>�ECO�J֥��O��w+����M�X�A���[]�`t�3f6�@ޤ�Zi����
>J;<g[��?8�-���Q6��
y��طw��4@x���I����E#�,���i�ܰ�[�
�M��"��&��RX�'�п-c���+l{}f���w��afzRJ�du�fFZ�,,���:eR�t�Q�;����^iۜMP3��cyk6�*�n�:�"�LF�|T/(&��&Y�͎d5y��e\�^:�3��1� ��Y�K`�[2��*����swla�B%�m��O"p.ưLx�?�[p�=���׏(��Ϣa���(_��ҕ���mj�'��g/ݓ8��P�S�;�aH���1!ؙ3gF�X�'ܤ����̟p�o��b��_K�B�ݓ��J��I�1i6����[uAހv��k�Q�Of'�����|�����G�>��4K}��~=x���������#�<6�(�á�)$����c��/�5 �4��\��~���-X��<
7�E ��(�ɋG1�P�Ng���:0jw:���;Q�N�NM�}�<$�Ω�Vtz[��1&Yki�,��hx��c��T��{;�tU�3�*����n`Q�?"VW���G���g?����T���RY�K`�fΧ]����!�!�v܅0!1ձ~(g��qI�<l�d#��q�
��Ö}<�Ɍk,�a.C �{�N���0b¤�9�!G_�b_M+�p�_�e���O��g�J�H��`��
S�mkS��
oK	͸��*�J������F
��R��T<gF���sI�bݽ�n�K�0^����I��iգ�L4�v�4X3��z������E�,� �	7�����\�S[���� & �1̂��B��4���69ü�6�%-��]���Mne����J<[��& ����9P��R�[n/SDD)W�6o��p�u �ȦW�s�1\�fu�7�"ð���k�~I`i��
��&���؎��'-p� '�/����5��?M�FX��9]����ۆ�s��w���o,�u�%��.��]7��������
��e��b6([��"���;�b���ݟD��~Y�y�O�q�H�9Tv8����q=TT�D���:Ya.��'���r���#�Qä�HD���T�����V�ԚN����O|^u?�h�Y4�A�T���vx���%/O���EY�D|G���< ?g��(W�̭2���X�<�;B�_��$&m]� �����W��:���Ը8!>O��v�h��P���ul}�#Q���r��8N,2���bc�a��p����_l�N�h�����ϴ��`cʮC�q�����>�Aq1*�Č�������+��@�	��
�`d�I�����>C _A%��S�m-x.�X�3'����[��sO+5�?bǲ��� 9�k����$�㗬�/?G����%������޼�)l��+"8��p��ip_��8�F�,��q�w�Լ�b4�y�赛"L��d$��Z4����m"� ��A�$� �	�4���l�^��CY6�����<y��-��!��u�+���J�o�6S(Q����V�b��$��0X"�e�F8��/v���e� Ԏ�2:�		��j��~�JS -��\�>�r��7MQ���=U�-��u��� ��`����R�&�9K���ʇu/5'�6i�y�#�8�gK�fl5\�<x3��@qs�3��)<{�A{tNXt�+�� �Ա�9{wZ�'ܶw��ҶZ�ٟ����E}л�Mn X�^��Vk�����<��B�,a�:C!�$I0�`̞�`���4r��(8F��/\9׫�K|R����n�z��@>�l�\۵]u⍆��ʴ�c���:Q���
�r�Z��b8�VlE8��D��4�
@��6L4j��d�i�p*)�?6�}�c��sk���C%L
ث�"���j��,׷�� Ql,�$���.��f�ULE,뗂p�o���U6P�C��2W�^m��%��O��ij���2�ޞ���/������u��3Fڡ�Ќ�Bx���sR���f(rf&ǖC �1�`��A���_x����K����s���j�{}�
pv��+����%�:��&�2����*�Z-�:��0���r1t7$p�1�� ����W�iL��t$1c��i�+�8�C����� �,�H�&J��?1Ӑg���Q�@Y�� WEZX��a6��r�<3	2��e���SRƫ����q���A��'���5��X�'�vvvl��[��� ��~�(~SS��k�t�LN�2Y�2���1�߳C9ȳ46-�t��X_��@���۹<�7�5�p�����f������3����]%t����������`Kg��� ? �5R!]RP��&�Z��~���	ꡅ��N����-���*���۾�ӧ��n|	$1Ʉ$���d2#�H0<$� ��i�'�2�(�F�B	((`��0��2���`�1�;vb��۷���sٗ�V5���u���9��3���ڽ�����gkժU����̌?�_4�!�ycw�`��U9�NI,49&$��^���5i���E�����rZg�/���v.�W�z��.�Y��T�!VB*�)�"4H�m&$/^���Ҭ���S�[�n�o������O�)�x��y�����<Mj{�j�j۴��>t�V�J.�{���_�bt�˜h2��5K�i�X�L�i3F�n�t�k�J����CŅ־�}��S">�67��Ez��B�����s=Y�v�,���vJ��ȿUI�y.�&0S$ֈ5�-8zo}�SeԦD�<�n?z���$Idۮ�6Ѭ���	��5Ֆk�,^�B��^���:u�Wۼ�Ҹ8�I���X�FNs���^Ow�p�-��e#�ȮI�@XT�~W^��H��]'j��&���ٳ��	>`�?����btss��tk�n�I�,R��l�4>�	�e����k7�'�
��Ћ���dst��)b%��EJB���5i���|��O�:�c{{]Uu�y�l�dDԤZ�4-p\O�h{��v3|u�M�uߑ�l{e&s�k�tE�I.���|e�غ���rr׉�̇C��b���s6O��)F����/m���F9>u�L�x��3Y�c��>�D��X�k��z4ڐ7'[�c�j�M�Y/���'=5�*b��$�֕����]��sV���Q�M=f�Hĸn�T�B2���n?��Yڣ��4t�9�˳���]U
�=2�I��l.��"�����ɩS���33����dT���������~��iV�N^|��cJm�8}��UI2�j�Mg������[��r5���ܙ��ԧ�T���!�9��3OG�EO��+G���
�����'[�+�^����w6O�����X,����ʗ��'۪�o��ۚ�4�
�d��R��֥��˗������������͑#\<��߬ݷu�omO_=v��@��63ץ�ku��W�%����ħ~��JH�h���?�㢝^'�V�~d�K�)[�IB�6P*y�������7N���|JV�T6�%�_��Ym
R�/���zÜMŔ&�T^��+�$���M��cLܘ��_��~?�LUŮ�ujm�6Չ,++�|{�y�;�^m/\��I�7��b�(
�S{���O��a��������DW�h,�_����¥����?����4�++[�k_����P��5�S�H��x"Z<��ͭ�	�{>�_�X����?>O���CN���K'~��~��#�<2�ζ"�A$��@������n�?�=�)���[5=;ޞ�����?��ϕ'׆�p59����l�X���'D�U5����؞��������8�n�D��X�8��:��w���'�"�ۄgZ˕JT��ܤ��ͫ[���g.�SH�N�k���w��ʻ����ͦA`5�p�ܚ�ſ�ru�#�_y~�9�Y���}U.�v�����{�a�%y�`1��5�V���ի7'��[	��m��6�qlm���={�,e�#�<aB��9��#��:���^[���my{�*:�ioE�~O�����4�ɓ���#���+Wo��Ѥ~�hD��E�B3O���Jq׋�_�g�+�)	0��J�T����V����S����'�s�֩�����W������'�<O	"KE���_�DO���7�{o��omO���V����M�̉����7$��i�b;-+�A�����v5ښ4���ѱͭ�w�,�Oc��7_�"n\��|��_��_y����6"ч�H�����_>=��B���B+۳��zP��o�8�~��{���c�AoR�\׉r�S�Dz�7`��MT�2�j�Ɔ�s��L�e�h8"�#�^Wl�J��{˖�x�"��=��Ʉ����R}Y�x%�}w%�l0H�]���oV>蔈R������l�� m ��7����~V
&S��Jmqi����H��N0�ԈoN-D�(� ����D�O�B�'�ɒ�����Kح�������Q'��|c�,Ѯ�m�j�{��M��a�;!��Y+�K���n@�"qV�S��d�u�/���xɼ("��@�c�Sh{��'�P�i4z��uJ � <,��+L�s�r�j���3R"�H!D�L�����k �ޓ'O^�������7��駟~���"�G|/"|`�)?Y��~�ڽ��~�i�i;���,î��x�	��{�q���%�q"w�X ˮ,���J",�vt���go+����%G�p1�Um����Q����5�m��s)��i��" ����a�0�X���7��jSv�ô� �@J�;t��?<����L�4&,�>寚`+k.��6�@[�N�m�4T�7E�6`�4KZD8c��/u^.L��&���y�` w��L�iiz�RU���2��-γ���f�ia�Q���p��m�3�+$��H���|���.P��5��6+�#�e](�T�Q&U����!�������3g^`���C$���yksu:��K���L�:�Abu-MP1fB�N4טx&�"�Z#�e���K X�$y�kDt�C���ly�i�F�%�Ъ�ZY�CD�L����wK~�!fMc����C�(ȷڻ\k�`{*3�q.D"hɈ��Hf����4qGgH� ��/�E#M��yLba�P*�Vl�qMDw+f;v���NT^�zm\&�}Iڻ!�[�ji�?�J�����f�҂��]�g	�&\π��q�V��;؜���:�ݔ�I����׎;C���,�b�� 	>0�!�[�xY��<��Y2�;3�3.p�'H �֖I�n]8 aM�o��-bn���&"��+��͆<��\MF�	U��ZC�B�*�"[��2J���8T��lmh�y�C���YΒ�/��:�q�m$3s���o���Uض�<���-_��v�'��趤Z�����ˤ�1���҈�4������9P&��pJ��1�"-ߝm!��JuH<φ4[W��5�0=�q"h���L�D�S�qK��UU�]�7n܈^5"|`W㶬�!n�֨kء
�D��1+8Į��B�1��S^EbXV_�s-�5�(�I���%�mC���ڻ`VggD()�@��ā�3Ң]�a	31�Υr�lX!`k����������
�ś�����־�kM��������y7�J3��k�Ԛ���I�Շ���3�L[7�K����&�Hc�
�om�F�z62?%qo�Lƾ�j)�s3
��^�&�Q/ئ��YH}����s�Znꕕ�������^E$���Uݖ��s7tlF����:��:��_z;�U=ϣgVî�Կ��=�Wּ>m��Ě��*׎ֻ����u���i+i;��~�z}��������IU~���� ��7J���O�;�k����U���&m����Y��v�
}���\j5��],�g�َ�бy�F���������R����A�G�fx���="J����;��A8����n��0�䮛K�A	�7YY\���7�H�a"N�#�b�G��p	>0ؓ��6b)H���^BE$�0�������7 "�D �/q p`�W�e�M2@D���#��F�ި���H���~��ˈ��E�s�α��	>0��68�mЉ�X���B�J)��ׯGM����u�o���Mz�"|x�?ֈ�@��"�D$��`��>b)��Kbg}"|x��Q��88"�*"|`P&(z��G,|�E."�����<bYp㇍N,"HD��q(���,"HD�.T��X�7Ѷm\�	���C\d�XD�v?�Pa"|`�&�����G��H��!ƃ�8`�CĂM2LD�����@YMM4a"|`�q��"E$��M4� ��1.`D�q�SĲ�&R
$"�g����#�F����h����D��F,(�����C�8`���
�E$�0�3K���-��Cq ���#"���h�,���E$��m�o��E$�0���"*#|`��
"�x�v؈&"�G,�h�	�����G�戥@/�[�/�"|x�,�+�8�7�<(��>␈��F$����oD�^���M5��E,�� `D��DqHD?��	>0$I�ÿ�Eֈ���m�A#|`�m��F0�D���x&k��@�{	����w�F,���8"�,�څֈ�� �=z]�H��6xk�����>G$���X��"�BZ�B���">���X�X��ݰ� 	>0`�/����g��4��(��{6��;>�v�?/�v�g��mA�{���ui������r�}�{�X��t�w���E���,����n[�_�g��w�h��ōq#|` ��UR��~��a�$��A�g&l!�"}���u|�;���Ed��	���WW�2d���_s�[$@�i��|�ؽ��	i�B��tn,�g��]����=wͥ���W\���Cw��#�,�v�DUU.�RD��?w�}��|��~^��v�u�Y¢v �"�^?�+ӵ���%�.�v��k���������� ݙ�+����EY���&�p	>0 T�� ��9���&v�����ZD�y���<(����`�ԝ�� _�|���}�up����t��,u>��-+�P�כ��4H�0��_YYџ1ή��.��qZ�q-��ө����g�fK~>'����(�=W^h�]�Gd�|���v��={���ُ}2���ׯ�۷o�" ��o����ĉluuU�d��o����]ڬ�ٿ�r��>v��q������F���˳� ����>1�9sfFή>��ʕ+����eЗ�'O���@��������u�]w�>a\�c�r�|��_�p���y���w��[[[������}fhөS�عs�f�������͛3����dnA#"8D������s�����~���رc�H^{�5��㏳g�yf_m���A�(�C��&��K/��{�1M��������q����1��|@�, ����^��ĝYb���L�gV�����W��	�k��b�x�;���������o���k_�{��g���0���w�x@�cz����/|�mll,4����������(�������?�nݺ���	[7>��p�g?��=�y������|������i�=�hE$���(�ӂ��B˄��q��a췈
"�f�4w�}�l���s�-m�v )���-�	���Iז��A���>A�F��~�i}�O��i�)"/�:-z?�:�F@��ْ3�`����"�O�ȇrP�3e]�zuG�n�~ ��0����S��z]E>PD�]?xG���k��t��;�ue�e��Z�tvx���e�EF�q�A�L�v��uķ3�u8Rs$�T����N���{������#�En������W�^/~���7c�1�=�������&PD� O�����*��*�T�'�E.�NKt��w_S��G���E���^.^(��.1v}��"�>CӅ�u,ʷ���_��t��e��uc���g�� �i�垏~(�����ܸ:���{&H���W:3�a��H���k��58���%���/`�D�Q_8t��Z��Ev���x����Ϣ�D�]�?^�h�n@� PG�~��u��g:��^]�~�MZ�ӷ�����p�px�u��3��$�۷��d��	ܑ�������3M���N,Y�#/����e۴h�P�Ce���r%vWF�=���������8�J�b���	>0,�E���}B[NC�m�Ε� �q���};�����٭+8��i����/Z3���]���m����S�]�ݟit�:ݲ\:?��	�G��~�K:��+c/3B�Ⱥ���/*ן�U���e��i�NX��,��u�)�/�0B����ٙ|�����}��]y��^�����#|`��w�`�;m��ؗ���ҵ�d�u�s�pd�� 2���P�|��cQrY��&���j�6tw�v�2��c<0Yd^Y�޽���ǵS�>��{��"�B$�01��EU�m��	����N{t^3�,�{!��l\�]-����X��8�t�Q��;��xxA��D���y�76������Ej�������	tgNc|�8D~9v�a��~��"|`�?����������l��~�&��e�<��.M|v�rWS�K�tBă���ru��aO�Ʌ+peFP8�~�E�1^n�v���v�:������n�tQ?�������շW9]���`l�B��B#)�'��H����������꫚ �������讁h���'�d/���l!$�݈�P7v����o����d9���ȏ6��/��� ��v�".�a<XP� �}!�ߵk��Ȋ���׿��qAϰ�!��n\��Ǖ���SO�Pnf���ᢽn|P/�}��U<s�{����'[�d��`	>0t������Z!�l� ���,ҺQ����� �-������pD�� ��9�Mh�~̖E��i�O<���f�:p�,K�t�.]���q�������Dz(��8��������c���/�c��?;Y�=�tPg��2\�P�=L4q�S��8����j�- v}�A4 ��L�]���)��!݀`nwk��~��f�f�~�%p�����n_����5i�n9�2���!}�����g�q�x9��(D�ꁮ�ú�F|� |`�ƃw?z��X�����]s��`?���'�E�J�u�EξYĕ�%����տ�@Z]7EG��~��J��Q�����~=��&����P�2����d����H�ab��K~�����ny{aWkt׀.�uObګ�E��B��㰮����]�X��[��0~��l�w�]D��U	i4ф�H�����kjXd����ȯ{��$_�\�ȹ(f��ձ�M��.�D��^�����}�Op-�������y2��������TVE��0"�x��߻���t}�g?�"x����}B������o��ۏE��5����D{;���][]���͆�=���o���F�@	>0���{-�u5n]_��/w/�w�Y�^��~:_tw��eZ48���K��!�)ŏm�6^�UF���`/o_(�c��]B��7v,�N�l,PD���V���bY�!/��׽��܋�z/�w�����%�ED��澌�l��B�(�E.�{��M��3:�/��w|����b��	>0pW$n\�X�`�5�@��60(� �T#�L4��d���C$�������8v�&"@D��M2�h"�i�q�0"�k��~��"�hF$�� ��ud_D�>�,j��"|h0������m��]����m��v�ڳ!���S�ԾV!_�X��N
��H�v��}ʑ�ەu{���jϢrv�]���������~u�����u-�G�a���+�\u��,�"��H���g��I4�h�n��~� r�	Z��'��ɥ�ƙݼD�Z��2�)ĖE:N/�\��u����������)1/���%�u]�$�L�Xv3����jFLh�df��K���kf$�21u�v(��V�6L�,'��W�{ǔݜ��]�  eIDAT���[Ru�_���f��2-p�u�zC|�w��i_uSOjG�D.��7}��''����='�3Q�Ċ��'P����3kYM��e�&�i[�u4��H���i%EbB�*C�>�M����f�h���5I�&�!$����2_#m)E�ә�&���|W��y.!���U���ۤ7�p˯j^��͈�y�fAU�S�iEB'aM[�2��"�u}�o�8�պN%��6�Znڜ�����7�	 �\A�����*O0$���[25����n;�-1��t��`�g��8W��H5�%D�Y4��H����IJu������b���|����1��0���i}=�G%�S��Z�k��kۦc6������AH���C����М�m��h�A
ڿ���iX�D�-�;[��a��\�O�A�t��_�CJ}�N�q+��� j��p�u�z��e��s�(�����&uy�͍bN�9]ߌ��)�X�f<6 ��z)>�0�&�0	><*�Э-q~�s�&o����H��5�m�7�qb�P�WY������z�<7s"T�am@0��M���l��JA�k6g��>����m�+�Zs��͊�d��[[P���t#���l23^͚c�����u֚yR��YϔX��cq�Ml�n���c��H�5�O�v�8���e>8Q����m<����H������۲�9��!��[��=�� ��R���ϥ5D��W�����sk*!�ɵf.�&��S6�	�}fqz�i���3�N�������n'3C��!(����8�u���ފ1�4KV�t�(�|n���X�|��%�����n�c��[ImK�6d���sj��+���Ӓ�p-(Z�Ϭg���Or�Bϼ�zk'te������Kr��l��*���`sf5Kz�8h��ق�g��d�[��Z�����I�Yc�`J�J*D8eF����Ѽ��f�-xOY���$�SP+{�Q�pܕ��2ۖ�ڗ�g������1V�,)�ֈkm�a3���^>n�A�Zmzd�HQ3p�G-jڀ�6ổo3����1+�Mg��_��e��M5�3	n��j�̳���:j�7̴P�Q[&�S+�"��Ԕn۵U��'!t4ɸ�&"�!e �!Qș� �0�1D
)�C�?�)��նbo1Cb�cR�9�4�c���,�����Fm��}&zD�����MfM���@>�(��$#-Sh�&C�Ը��elגmX�Ar��չ�r)=W�YH�~Ia�vЧ�2�Y�%Hԁ���#��IN�i�0�h��A�TfE��Y��# ���	Aq�^'����ř�,���+�v���0�� ����Y����U�v��%4EJ��݈J3sC�ڔR�!����1+"(�}�m�k/�ޅuk�XHS=zM�G��B�Q�J�H������D�cCh��l<1&ALӓ&������n����P�I��Q"Ի���lۂ�Ը�Aod"��Ґ'vɰbVH��c��L�'�%"k�܅��S� BlK�,%ү���{y���!�5���i�N��]1��Q�	mN����������ֶ��d~8�!Ԝ���D�n�of��ꨨ��)��F��T�3����ՐҜ��OS�W�,���/��}�%��2�2�,������֧���	;�'��9�(��fUc$�;uaP�Mj�XZ���09F]8M߆�����U��`�5��J3\�-=30s6Y�D$���y+�`�;���*Y�ț5�U��]B�'�w�������+�@c�v掙�	���;S���]�m"_�&Ə�7j�z=%D�T3�l&D����3c'Śڑ�#�:Y���N�O6 �N��,��XՔ�u	5�v���D��2�)�k(Zs5�$�L�j�N��%CV�6!��Ͳq^���Bt&�#4'{D��O�-���[��� [Y]a#*oJrTn?m��ڣE�`Xi����,�fSj� a���$�G䜦=���H[ޤ�0�6vA��Zz.pG?Jm�k�cͤaeY��I�
Fݲ^�1Y���2�1�"J[�f&!��W1Ӣ1�@ٚTl��va�%	����l8`�T�F��x�$��&LD����E{���&�1�_�	�#zݷΈX�&9M��B�&DʔY��Ԛ,�k�	��7TLr��=s7��)b�!��
���#��Ŵe"/(]C�ݾ��'<Y��l�j�͊A���-�cV������C-w�gl�$,*�5��K�������4ߌtiٲ�����F�)�˩n�F��>�A�w_e,m[�!K���r�Y�v��o����xTxZ�
��Yգ��k!�Mmn�A�Qܖ�QR� A%e�=��h��q�ܓF�ڟ(N2M�Q�����+�Nglω4�q8d�8� R�Dl��y2�fG�ڕ�K���	�{���?�k`&�m�1�����{��P@ՙ�3jcA�������'���|�lKD�����v�z�8� ��C�P��5i\Bw�ٔzj��kں�����㸽��l)��+�n�M´�cf:��jM3�k�<%��(=F��3�x��7vl����yM?�j��&�9��9Z2�e�K��'^�uz�y�D�P_�;��F��H�!5��vGT�
�]��gi�:X�nb?x�ir����D#��ۙʬKcb��hW�jz�����4x�d3s���
�b��h����I���q~P{i��,�)�n�l`�h\��ڦ�Wf)�9#�#4���9tN��;V�ſ��)�|0˅\�V��^0n��E����Ռ�166S��w��;ԩ�l�F/-ЬIB��~�z��Ŗ�fC(��fMH�ç�(C�H����-�}nti�ݞ��&Kh��\�6s�yf4~�Ӯj�JrD�gߕ���<�u\�UӴ��4�7Te���j�����9%J�fm��qb&�X@��t�B�FӐ�mf;HM�=�ѥ��y�b����7��f��v�����,�W��n/��m���as�K��Ԍ�6�HS_�v�I����6,���s�9��?bnc�h��z��,e��]�<X�Q�y*�M4a"|pH5��R�pzll�˹�L:�;�K墕X����vo�Gi)�%`n��z�<m@Zܘ`���'�\]�n�Pp{�ٙ�i��^h�������W��S[w�A�|nRB�$�|��* �Lr����vh��2���yxC�3�v�Q�_ʍ��3��A[3�uc��Bgƻf��+h��{��7>���C�0G�z���##Ȕ��'$(S� �Z���\5�DJ��,�,"�s���ۃ2T��*�2t�
�bbꎐ"�WD��!$?�TkMz���7��ǣ�3'cY�j�V��~��&��m�f�$��
)����jR6�#�&b�_�vg,��G,�vq!��V�e�����������)<]�e�f.D���HI��ƣ��k�����iA���4ɷ�9Wr6��(�~�n�Q�\�r�B�L��8�]G�da�X�Qh��4����i�Uh~JO����LI��C\� cLKU�q�ٙ�)�p'�zתf0��Ie=��;���"|hH���������fـ�ʆ�Z]�)��e%1餗�r:���ηڸI��J�3�Y�huX�<�Y?��O�8�.|�+���DL�1��t�K���HS��
�S��[f��f�dQ�����+I��ҳZ+6?�:T��?�'K�~����0!��H M���bŋ�Ҥ��u�y���6�{4&���2jKcB�Q%5�1�LXY���ŀZ��&,oM��E�
Ҏ�<Ӓ.�� m�l��O#m_t���>W���4��,8���ya;�z�L{ؤ������F�M|!,\K��Z��-[އ�ɍ{�6���L�[�l2ݦ���C R�T�@l`H�hr�5�ת"��H��#J�\�G,��JaA�f�ͲfoїZ���R�\k��H.E�F���^5�O�_dl:�AFک0:<����)CդZ;ϕq{�N��9v�h���T�L%*%M<I�&u�����٭�b��#"q�E�z���|���L���b+GzZ���3 �Z�l����S�Z�C�����?�+�q�T�03�$L�9�H�-``iI$�&����$xbf��oP�WI�*��+�I�6�:b��TDܷ[ID��s�;E}�g#'̈́Z���c[� �B���g��4^ �����++����ɨ�F6z�#�Ba����[���4�'IO�o��,M�|��F��Ѝ�m�=�F�zSUS7���jJ("���T�,ˮ���U���++�ZU�j{ďYe���b��d��m��/�^���\*�+[�Z�%�/Jk���V��r��W� ���O3�CFIyI�DZ/�<H��s'I��p��&혴�4m�O�
i��ք=��J �d�`3)+>	OV��R]3ٴIB��:ѱY IR�6�|E"�^�$�j �2M��;&��{V��4�HDGnq���3��72>MR��J���[#6XY%�� q>.k!z���Ƽ�Ī��^%44�I�H�#z���T��V�SVS��OD��&�)��+2�֭5��p/�m/I���W�J���"�	V*�⩂],��*�:�>r�S�:��p�Ңh��V�_�f2�j���
u{4�g�㘙HH=J�pH3����'��T�ʪH��IW�oUU�q��q�"�C$��@Z��b��D_O�V+�E�χ�C>�LX��q"N����h$��E��"#"��CG��bY�<KSQ��vc_���t�֎eS٨�Q�Q��#�?"����Fu!�<ႄC#R�rlH:���!S9Y�`2�������)�S9��ԁ�l�$�3ci�y��$#�N�<�XtMYEmD�)	��A)��k�|Mm��,���9b)%FD���>��aX������}�_Uc��D�D�$��Z�ȩ��_e-9i��ԩ�|�E��Pr�#w\1���j�D�ȔO����l��n���`��U�^Fϧ�� ��&B�eL�������b��O*5����������Ӫl�� �(]��b �r|��ֆ�M��x'�o�, mii��G�*AS4�e����$�^x��k"��_��_�z�ڵ������{��������D�xǽ/�t2���kkkk���q�?��'���G���}?��#G�K_��ذ�&TV��
ޫ���l����_ۘ.���"d_ۓ?��?m˘�>��G�{��8����?��o{�G�H�!����GIX��.7���N�������>�g���:�I��W��Ǟ�f\fk�5�.g�9٘��?��̵c;��.����sϱ�._��#g�q�	��U$YӰ|�_��g�4[0�b/?w�=G����?Ώ��Y�F���_g�_xa�q�~�c��YU��{��c�X�"�C$�����C�f�?p޼=q��w��'>�Y6v]�3�w	���g{��엿|`���3����H����~oe2��?����坔����󗏭W��C=t�N4>B)i�C������ߞp�߶�ʢY�*�Pj�|G�eݾ}{哟���C���,~�~kH�Z���?��O|b�� Ԯ�������{n[�v��c%����C��Z{��(~��~���_����{���/�_�"}�GN>����S�M��������-��<�K��K?%�|��}�?0��wh@�����US>��zWy�o����}b��?�ó�|��'���_��������?K9���p�����ɟ�ɿ�q�ֱ���O�o�z���7�>������GD�����y�Q��*���ī���{��>�H�o�������[wBV`F��*K�5!��;(���}�;�d�`�����w�)�Z�a����es�؅;�n�~�wVW}�Q���v�ś�nݸ�����_�jz'3j�<����/|鎶�~�_������K�~���w���g��o��o�mA�O�c9D��=    IEND�B`�PK
     $s�[Q��0�U  �U  /   images/a88da2ca-7e0d-495e-a5bf-cdc1eeca5e78.png�PNG

   IHDR   d   �   �M�m   	pHYs  �  ��+  U�IDATx��}�eE��{�ݯ�LObf`��$ad.�	Y]XWQ\1�((k��]WWpwq]�]&�5�E�I��Ȑa�c�t��U�שp���h�k����u�Su�9�j/>���k�v���xZ�N~���� �:xQJ]e(tuH ��0ٌ`�e�o�* xJ����^(W
 8�HH��"�h�B#��(-�O
�R}��Υ��_�x�/PW0����Z�6j��3��D� ���zܜp�H ��2��h&c ������Q�ejL1�Z!��� ��t�>gh�rY�Ѽ/~�D�� ��R*����{Ċ�+��� ~~�Mp����_��𶷞}��𠹽{w���������Р0�4pp��Ȍg��p�PdA���6�g��]4��!�I�;d������ 2���k�lڣd��i����j	������������{�����a�Z��o���ǏC�@���������oh�(��d��Sh�h�lG�����;�����o��}"�'�'`�-�Y�f͛�����_�^���ܓ���'��`x��BF��d�`��4S{*��.��9��/g����ߝI���T��c�e���󩧞z�Z1×~��n��g�dooߟ!�tK��X�c�U�һ(�!�(�h�8I�.IM�-�ӴAs=�$!��tJ1�e�H|f����C;�����'���|F�{,��L|���!�y��c�]oT�<��ɩUk׮=��h^����֭[��o;�Vɽ��y�s��y��ŋ�{��ժ#�A�SOb�`�N(�J�qb_���w�"�:�/eNc��/u�f��� f�� %y ΄��=�K��$9���Svh�=J(0�Nu��@����wl�r��ŋr)�Q�7� ^Vp��R�2�����3��n��!��t~^�W>���I�Vԁ��۷'�w�ɤ�ǵZ�Ҟ�������+d,�p�A`�]b����cǎ*���><�9�4���!�6#¤��8�{)K�ST�Z���dOOLL��C�{������緶o�~t":�+���I�U~�P�9���Wp��뵝s8�I M��v��;<�&�~	��%�H�#�$��1e[��v�8���<D���WRoo�Z!�z{N��H�"��sS���'I��Sk)k�?1\ĭ�'��
���J�c��5��S���%�Iw�E0�T�˜�,bD�3-/#��1/�is����b�ۣ�Uˉ$<_� �!\"bu�>�鬗����f��G=�Ԍۧ>c����WN���9
����#V��R���דkx�Oպ��*H�Z|�S����.�Ӫ 	-�e��D/��H�[��UO��N�*ޞi���2u��F4 ��Tߊ�s�s߷�r�8e��{(c�FH��5=�P�����'���z�
�����rd�]��^Yt�W����R��	�4z*4+��P�!$#G�,QHU'� �g*c��}ߚ;t���+[�9���R�]��9��*�#	MM������9F�Y�֪�����mk�&Ec.��؝o]4��#�ꩡF@��IVآ� C��nDB�	`�:z�����8Ozjʴ2K*��=����@��'D�,��t����q�}���/���-K�D2�Z�4+!�t�j\G��W����kj�#��;������|��j�I��H)*��0�>�K&��45���^�s>|�׆6?�A`d��o����/R��P��Yˎ�p=�����c�V�k7}�E�~��K� ��8���79�a2:>OM	!|!I���9%����ܼ�п%}~�?�s�ҏ��mG�\���S�+DiPFv�Yڔ�t�7�Z��4֌�q�N��38(c���	ɽ��������{�B�꟎���0%z�!!�����߲�L�3�8�T��p'�O<��j�0uC���<�]ҁ �����;�E�ViJ�+=�/�Z�d��GhP+��q4��������я���+�pTA!�8�Q0񯧧���dk�w�<k�s�	�@:ŤC�����쓤\�%*̚���O$�Mn�]	��V�bɧ��+��>Q�R$M?^@L��!)@�O�N\��Y
��|����~�O�C�����K;V�7�埛e��f���5��V�|�-�á���HQy5� ���a���N��d]�kh�
�kI%D�!IEmW]���^�פ��ܿ�W���2j�Q���~�85�@�(�[�z;L�?�<D�	����
�Z�
YD��n�z�m�ȌEX��f%6j7&+�9�@��}���W�Q�SQ�$AV5���ñ��3ڧ�xw���.���|,�Ο�j|�#�rY.ʥ�vM��"��B��^h��d������?	�I^�J=���$I��B�/_]��q|���f���y <A���b1��hY;}q�%��D ��ET@/�:����W?���\r�d$�pM*� W�q3%\�MTB�z ����a��]͸�y^����Q-_I��D�;i�)�#I��/%���pu�D`��n�#�N�%�c�F�|���7� ����()]�MjO���<x�e�\�㯭�RD� I��c�Qb8f��j��Y!�%c|KN�6:Lpd^%�p���-=>���\q�{�pҮ]'#��~)��F"�F��J��yγ�'^61U�� �����kg���`��� ϝh�S87d��MO��Z����&g;�����d�HtA�~�
��A���jx�y���f�AH>f���[�Ly�&�ZVJ&s�e5�Q5T4����b,f�79m����"��cpz��K��$��P�DK�ӂ�.\uo�
������3г3 -�i�x�=m�!�]L6�|x�D��=\�XUk�$�V�Lt+�SH�&�3�X�<h�/�q�s�KgK���|*>��-��u�eN�r�9��y�ppʝ�sH�4��5k���+�%�Q�L�L�n5����>�@�v���y�D�5�/$�bzo����R���*�S�s^A<������s�G��3)�qe1�����#���uu L�7W,����}_���ht�����޷AI��јvmn��1�U����դ����`�lRdLZ|�c�5�v)i�N#$6��p-I�#"H�=C]��E����A�	���r!����
�7 ��.+�i-���<��B���(�ӒS�!��H���&�ȼ���O���{K�љ�K��J���&<�E���߽픓[>>��"�v�����~��aӑ�eH�x����-�J�%��j��@<�,�Κ�r����B���
��Q�G�#�����Vr�:*�<�y���R������	����0/���2v&<������mDj���%5y�Wb��ⷔ� �'Ε,�l�3^�!��5��G���W��Kʁ=�<o��׳��w��1��,טA��P!D�,�9ʤY��D��gpߝ B�Ժ��L�21�1F�<�d1�E^�;,��e'/����w.����C���c!��T�H!�i�6)R���R�@R#�(�������5�"/TZ��b���u�u=���Ln��A�[��~CV��Wv����Z�Dz�r���+)�����v�#B�V����j����H5E"j�Weqj=���s��=�)�?R$.$Q��y2�d׀!��f�d� ]?9�;�#>6"�x��2U��Z�<'/���0j��Р͐��[Ԏ���������Iy
x�����c���Zp�b���$#X��]�)J����Gz��4r�3X-*�[^'*l'�a�r(s0��.<V(�5Az�sڊ�zj�K��P��v8s�1w�����h����[����I\�F"��P�q9�\cW@�G��Z�aK�3�Kӑ!+E1���zV�t�F����D�������vRB%�@�~�W���U���J��Bc�Bþ��|.��H�1/G���ዹ��z�gM���R���(�!���C�9f���6��'D�--$(�X��Z�����]�~w�#%Q@��X|������^'qr�*ђ_G�$H�$�;*�a�p&���o® a�T�-1�� ;;6by�̬:�_Y{��T�8�
���V=���bD�>�ݯ�����ሁ��+H�Uhf
���:�-e��<��AU��J�L�Y�8�w2�ƟBZ:>V������ݔ'�/#F��6�M�&&��F�cj!�����g1+iIp~ə�XR�!~�D�יD+v3��^����M;s�I7��(G![!m:q�9��@	9e4
3�wO�������Q1!)�ܔ0t:#���E�j�1o�O6P&2�#br�������4H�pf��KE�Q$%�l�9���0�b?i����y�eO�IfPv�YR�Oajr���b����1����`?k�AMt�!,��w�ϐ���q�GލRh�Ɔw�E�h�P���//�8�x$=����l��_�O��\�iXEAL��9� Kg1L�t��_t��p"~���XR����'b)O��s�=z����#�؍g���X�|�qT�Q�SG�_\�RQt�� �@3+�7��_�}�ލ}�����[���+�.(�V�~������T�	��;��� �?��<��������R"A�/�:��d��T�%y����]O!ĭ1H�h@P3p䫛�_�y�ّ }�:N��[)��#}�M�gCV9�}��>r�O飣���ȋ��,�ڦd�Uup��՝��/�n�:�1�D&/4�c�����>�"!�����}�ek��%ړ�QA�! A8:a���	���T�~uUC����}h5�Д[TD�����Ȋ��#��W$/q<d(�R��-�N�J�<�5$	y�H)rv4��#vqd�������:/�%j]�i�qZKgN�nR!���u$` A��Y��}$�,Qb�`�yY�zR����tҞ�zY{���gM��i#JlYZ�˨�YC,��9�	HU���QBJ]��R0�T�����&��� i���q	)j�Oq�>�9�M�N(I��ޕ;MM�"}v�9�h�&��b�J��׭m �Q�tH�2��S*u�GXA��L�$�p!$�(�3�U۱����{�1�E� acb����G.	��
��/�B�O�
HbiɁI�O�G�3x��ƍɕ j�J� B��e�݊B6�#��� �K�C�X���\�&�g���SY-���2o2V�.6A)XI��Iɴu!+�0zE(I��.�+�~�ժ�x)ZBi��K���Y�ۿ��~��}B���"OK���
�:)���B4���o<�3�8��V8�z��������r�+�YG��;��y��c�>Z�r�o��j�:v�:�9�%�v䛿WT��X3��lY�ax:���f�%�3������nmM��������-Z��ܬ�y��"q w��X��X݌Q�F���wOL~���&���k�)R�¡�9RH4s�4�
�����=Uy�1v��mr.�?��~I�30�Α�=GS��u֋�T��6|��M''�����X|�Ww���5m�/~���]RR����Lt�{�,w��!;tK��t�>���/���x�̓�Zt��7��I���Vtx�P%ǒrg�Gh�p���x�ݣ�{�X,����<�,SW�6.�ł��@��R��g�*q���$$�mE�D}�R��0�W�0=ݷ݉2�ܷX�#+`Tk�8�~7�,� S���i�����AY�����qp�^+v�1.O��F�����G�'P;R�\>Le��e��N�p�rHÀ������-9�E�t�7v�\�p'�i�"�^�qR:J�]yi�sn3�c��\��Z��'x�y��bZ���dF��l'����#ʠ+ d�^�Ra?�٦�k�n���	o�xJ�����_F�E��e�L)��`,!��$��(��ʄ�����2�h��Sc�b�5'��є1˔�v-i�-M\�&�Lԕ��U��@��`���lDI**���JR*UX�|L�:ӈ�C%��7���S�l������#���OD��:ΊX�]��Gq&�m�U�B0BD��,�(]�ig[�ǈ���e�A�d��f2�&''1��_��ځR�Z��$N��N����8b����?�
pu{86�a�V<�
8Fn1f:4�Ix�	��>8VVS��i�������V7pz���N�1�6E�"�����敚��@N��н����۴+a� �>!����sU��g�{0>y�t����w��{i�v�l��-�(��,%�u�\�d�A1"�a,�1��5�!��
����c�T��a�zd~��4b�c?��%�=2:��z��
�ظ"CF��Y��$y�i����
^�iy�ą�&��ϸ(�L�>�$�	 m+Y�#R�l22�W^�A!Ꙥ=|R�V��z�T4���>rya��U�1<+�a�����t~H�����s�H� ��}C�X���w��z����'�K��?YVf~%vc# ���f��1 M��
L�N�3ZT@f��}�dɫ'~�ej���s8;rr��OANF�wa8y�T7�v#+�~4�*A�������C��r�H��Lmf�3�0�Dd٨��8��;沇p`�Y��!e���&_����O��"�G��ekf�g�g�^��������^i�R��{�F9{MM�����,�2�9�2H.�Jp�*���c�N��}q^8���k��{"��3�y��T�Vo�Xެ#<Tz~�#~��?LYs_��?���!��Ӂ��|�<Dm~�d�.�4z2Q��y����	���%�"��#!��^X�.��q����(�1�22NxF��f+D���s�}Z��k��7�G���ly4�t�J*A��}�u�.&�U�c�V��cC���L�_�ߵb�{�09}>'��r�,�B��)F~���~V�9���Ko��2ڀZ�U�52j�;��d8Vxw/�W�p�M*�Ǔkߵ�v�Ow���+����m�j���/�2L.SZ��}hjXuv�MU�pVǌC����2�uA��Q�����{�ފW�(e�����}�_�Q�J���UON���7,f���]V��(n�K�C��fы�Ǉ���s��3����W@��בFT�U:���kA���\�~S�dȢ$�׊�#>�@��M����"�]=��|��}g�!��i:g�@�j�I�AO�E��� ��#�Q,�,iG�����!�Ɖ���گ��޸v\��h
����pd,,�K����e�r�v�#6�� e���%��E�D���j�I�#��-7m�A��O��p:��/�cLK�N�ӡ�_eH�={<*������#�);-i%��%;��a�:Oճ�_����c�s����H�|�3���d !(�?�yT�w��qS
�թ�9/��x˝�E��������NJ�z.���0���WH)��?���΋=����?X|�b��w�� �4!��307L=�a�d��4�rc�����C���0��K�6������ˣ5u�"��允
��\��!��3�7�4w�Ԅ�1��Qha" Q+�J,�[y�p�s���$�����,dTX�BvZ8&\�`#1��*���sz�~�����P�k�e^�>W��F�Iҁ��3����؏��I/�c��@D3�NNqu� ���	�I�N�?�����ޖ�׌�5��҈�+AM�$d:�:G2m�~���.������Ԥ?���\$+&A��zS61<�#sQ.�q���	Y�֩iM�S�����M�6�-��j�y��ҷ��&�i�ѹ�:���1]q׶�ѹ��B�)�4�mF�"�%���I�� cQkoH���	�i��>y�&P�&�H�0@�dIy�)	|�!!$�F*�NN������")�<��SJ**8�O)�0li�I����̐�Ț�:֢&���U��a���-lt���"n�R� &us�k�������t��z���F>�o�XN1#\h��=�x�^:ި�y,2.;p��<����y2.�s6�a����n���K�7R$< �i����J� �V�L��NF�(�0Je���'׏���Î�������5��	͆ޙ�(��%&M=�e��ap�����x��\�$^����'�ݯ[�.,]a�����"����KA,�����x���,l���m������ώ ��]�I�fF8Z�F��
=��fW���	�R3a:&k$�!��љ�:��'���ӔL�{�O�JN�4�LW���c�-��9dy�oP�i���
Q�#M����o����^e<&!�I'.Ca}��'�pt����}Ǎ��+e�x�>.�u�~�C��t{o�������{aj'�<a�U]vbȝ�UO�m|�k|���@T�P�]���{��� C4�2.z3�t4�Ĵ^�V��q6>Q`��tJ��{QD-����ܪSw���p����h�L�Fx@���������&��on��kl嘹C�l���['.SZ�v��f�!���c�)
S]�F����t����_���?
�a}�i�u����Y�e��������?�ڛY�8�����EFV4�-�O�ʎ�@>������	;��[PY��(���ڥEq���"���߅$WO��B�|u7�˰*Qx؎*�!2�i�dhAkPC���s��lL�Wq�0��Sc@���U~��B�%��P��3I�L���5������'Fw�����uˀ�U=6�ڽ-�diVj1ȸ]��B�.%�U��:d��m!R�:4��_p�)�]rʅq��M���܆&�2�sX_�2ֈdq#�xӿtU��}�$���W}nū>���J�0���|+ۀ�4=��s�{���=���(޴W���oX����T�Y�	K�]�ƕ�2ӌ�F�u1s��}Z���������B�5�����Y���É(G",B+��lƓt(�Q8Lh��_�9|�P,O�Ĥ�gU�B4�JT+�D&��7p݂�]2R/�����iB�;,��BR�D�5T�{��_���/]zm8�:�w�s�s[��^�r}I��E����hr��+4
��}��Z{���Į��d��G���?+��J*�����W�b`ڋ�H���$8����z��x�s9��s�!#�1�u�As*j:�D�7=K3���Jq�[y��>�a��X�(�C�d���j�8u0��INs�̟Q� D���1�n 3�&�{1Op�UVv��>><5�����jF|�MD�C��D	_�啾Cn�ؽ�:��x�h,��r��:q�cnz��#N��BΑ�Q��61�X�C�0Ъ3_J��T�E�7������j�e�$3W��0�d�ZOfR�86A�f�D{1�VQՀ��'!��b��rRTP+��ޥ�hI,�0z(��Ek?�,bt�����A+��ԲҰC*43l�3�+q5~b��і��� �v�uI��=�U$�EmtFX�FPV�QJ+���@� im�ŸML���K�(P�s�N+�j�'��LM�M�;1%9:�j3����z-�ɨ�k��B�M)�i)%�U�4@�Փ&5+��y+@�UE1���i@(u�Yc��|rL�T�mL����0j�Q�ʌ����	�ʼ��+#t���HcxD��8i24�}��Om:�4�	��B���)��~hBmIY�� �d2�,���N�M�C�m������M)�r;��xsOQ~*�·�$I���ޮ���Tذ�R�%։O   ��ŵ�
ѕ�]�f�_R�����/���b���V�O���xKA��xb/���qk,
�8xmD?N�v3P���i����@@\(N��.��dAF#C'���HM�H��I�i�Z��q�d�, [�.����4:� �������[ԋ��0���M[�M�32	�A��K�cq���j7��Tl\wh_�j�5����G��c��<ݻ��Y���<�o=�o�EC���.�ڹ$�n�D��c K>����5�)��퓪������D4o��j��~���*!m��Y{lS��7���"��M�n[%���-�W�yZy�YX����g�##U�\g.����$�TËa�����9}��N����*�ݓd�)�`��k�%:C�7h�!$��@$�����swu���C�r����&�X�ث;AOGȧ0l[�%
Q_�Wٝ�޼�v%]���YII��47�K+&.�=7yOk�jz.X�2Ŕ�P9yh!���V�3�D����:�NW�0u�J��f��������\�J�'����1E�`Ж#�v
�v�a�f
 �A;�o&%aO3�b��h��&^�(��@�<��e�T�M��z'x]/����֡7Ӑ���e���mo"Cq	�l��z��P2S�A+U���\��h|#�L�Y��ѾJ2���/�٭Q߂H���h���e�w6�]��K~K��dZ���y�gR��<��-ab
N��}~~�uD�kl}ּ�'��l*�Νؖg�Xئ,p]�Џd_e�o�Z�9x[[�Ҷ�ڢNP�����I8�N�Nl�)j��Sl���fp�!%9�w��\��̣����@�.0�d�Z8�ё��L~��^xKc�Sgr�w�$�]�����շ�a�E�1�x�s'>>^�W��:F�#���r$����Νa��X���x�v@f���mg�?m:�i&�C��*���Z�X=�@D����rc�/F�g���d��u9)N��Z�m�j2,W�5`����qϽå���/�YxnWq�g�� ��l6$�u��G�"Y,�J/ =� �]mҏ�n��7�/�N6��u�����+Z�i_!��E��w���`������،S�IG���J&�&�t�;��2�ξ7���d ��F�pbD��v���qN{��q	�Y�S�H�W)B{-?i)|�mʥs��/(���9T���c�z�jY��:'�73_L;	5��~#�4ii����pN��Z�����:�#�%��.4�)]�02���a/xuk�q!���B�~�����)͚N�5U�RX��/I�fm[wdE�X�~s9jR3g�7P��T)��{cv��]��Z�K�1��("�&�Ńȴќ����� �mU?��fT�zhG�UA���iMRj*���pB��Q�	�ޭˋ�V��J��?Y+��6
�WBQ��H�m�$�H�!�n`�d��ʽ���{��/��ojj����K��^JE<=.+8O7$K]���5�AT�xB�eR@%T�&�R��'CM.�F��(��N�Ihh��$�������+��Y
905��kQ0���I�����Lmk�����#�S��iK�T��m 1��%I���c��.���Z�o09q���xl\<ܔ�rz��L���<JKY���;��0�K7�u1a�6��Z8'Lն:务]�/���,	Vt/�0'It;"��7���I��,��$�E����S�	j�v&Ձ��\O����ܵ�FɵԙI��񭨯M�(�*}�S��S���m����DY�ɟX�fҢ�yӉ.��.z͕nA�j��(�OR�[ ��'����ø�S81׌(4稉�7:R�-�tB�7�|�W�g��� ��Ք"R����&��T*e�[� ��2�l07�\?�KǉI>�ŊyВ%����_]���hhӶ�v4�>��$i|	�3Q��Y=45�@��Ў=�p�(ǆ�wJ�]�����fB:�;R�Dv�������S��Q���?OG]�q��#�)z��fh��Y�����"���Iw6m�ޯ��R���*���	� �����H��Yҗ�#���)�ʮ�qu����\,��Zhj�5��eVoN]�~�5.)+�ml�b.P�����,c7qY,��*�	''^���N��e���"F���~�
�LW��O���ܲ�f/����I�/��{n���V�y��z�'��ٓ�=�̏^앺��c�����'�Z�,��Tt�1m��Utb��q���W��߯�Z��oB����t��Y w*���M����=���wnz�������ջjǞ?���a�uk�F*1'�S��`�A��& '�"�����-���p�k�F��o���� ���8�3Z����|���}���ho�K�8��toF��R�8��"]V,g͑m�����sS!ъvmS9�x���f4q{��2�d^��w�����S�J����c��iy^��/��Rkt��@��|u��B'm����%�[9�{����YfS0��s��!��R�$�ri�9{��k������������D�>s�S�9�C#n_( �O��*3uI�=��'e�O��0;@I��,���E:�>c#N �Zsjƴ۴b��4	?����Om�5���-����&,4u]�P$�?و��|f�uϓV����F�2c�֫�N�$�<�'��A�Q%:��H��TJ��3? �X���]%��rDK	JD�l>Z.4���B+�Eƛ��9Y�2n9+=���w�+#�N,�G-o���bXR_L��1�L6���A8�R�jԂo��;�G'Պ4%�I�鲹�����V�a�ੈ�֊Jk�����%�A�U��&��n��;6C�e3s'����
��rF&N�Hc��C^�뫻���ŋ����4/�b���~��nM�؎��~Y�z��k�ߺ��Y-(�t�9_�r�1g�B)'FN���?��>D�Cjy���q�e'V���kՋ4_0�r٧z+�X�{�PpO�u)�:@�l�u�X`�*7���=��4���+�O��{%�N���"o�tִ5($��Nn�����������k��o����ٙ�Ki�4g
vE#���?�V;C�z6GiE�.ǌ�,n��$�m�ɍ�� �.��W��D�G+��8qo�;���#�F�%-��C�L��h�
$�7p�a_޻��ת�n��\,U��>ODNH�ט]2c���+&�`Yo8���K>���[^�h��9�Gt׾׋z(/��P�ۋ0�D�`�D�9'9s���o��퇯|߭��}"��
oD����޼L�үp�0�	B��h�#3�@QӋ}��}0��#a̒dJ%�Ƅ���pj2��*���hb��#8�lj6�Y۷�$.TkEs�ϸ.��V�c���E!�]���H��"Km�,W�G�mE6"���tM^�D�V����
�z�{:�T�"���G�ޱ(
=c���=m���N�N}=��C_���N�nk��?Q�^ϒ���5q����.�K��J�iz�E�:\Gk#���F��s�Vz�����5�GGZ�q+#ۯ��	�g���$���Fi<0��B砨�w�	�|2m��vB�����H$a�b�T�;��4UB���m*�����j�A?��DD�_�l�8%G�c�WV�ξ�t�ƥ)$  ��1�*qrޢ�������B����#է�Q�C;����`i-���RL/j�nZ~#��4��f8��������M3uM����#�Bq���Q�tj0�����o5�-|o+�*�[���n���t�c��s�5H���𡹅�wF����C���P��BqQ�m��tɄɘ.t�_ߜ;���Ւ�aX/�.*�{�k�N(F�ew�ۤ�z�����F�$�hf��~˕��5ǜ��6�X�� �t�������,�h�B/3��M �m="��xb7|Ќ�S�L.M���eBc���w������8|�ڮ�;OQH2RD��H��L#��mշ�A|�D���j\���G�L�gj�pj,�9IP"d�p��I�a�*����x?0��jN��B���Ś�S���_NE�O�V�Y�gH"����j�Pܺ�H��R�ã�l\K���. �`{bxv�κ�6�8�d����i�G@+�YTH\0类�;/�<��4�KK���9��W�E���é��if9K+OI�y�x$F�5���09Zzg�xP�r5���N���9S�3#��e;���b�wO��Q
�9�����T�9�B�0k�o�'&^4��*���ܸ�'$�/0�J`��2#����b�zt��>��R<���:5��XקM���(ɭ��ҁ4T��o�m��`ޒ�4���5��n��Ҹ�V��(���y�S�95��Vg�=a�Uݻ��|j�WKD4C�*��r���&+���F<�����{&�R(�P�u��]�{DW��8�x����{B����Z��W���7x�{�&w�t�S�F_}05?C�#��՛kj�/�מG�:a#�8�}���O�#� �����8�P���z�Ю��'���I៝p��WUW�����|Ӿ���S;\���j�׋H[�i���^��;z�+��������o����)3�س�%�e��zfW��;׬��N��58��,a=m6��l�"��.��X)¦�_�� hG6S�B/w�\:�ɔ~��hE7iw���v�?�HY�<���M���}���@��_p�3^~������#�{�>x�_ޱ`�@e�P�.��֬���fQ�Ü���$�&���.��)�0���xq�5wL��6paplD�A�Ә�V+�����y�5|R?l�y���o�F��z�o\���-�q"*�<h��s��=�E�K�Tl��W)(�K@\,�C�m땱x"y�=��5���d�ʬ"��V�D����#�n����o\�%{��'�P�߾ş���4� �^.Ň��T�B���xaK\Z���i��K���q��-�8I=��2��,R?�4�C�֨(�O�-����AL��SZz m�=Wj%�^򔠩XEA����c�+���{��w�Qݟ�>� ��}b��6\d��F>#H�t�>]��e�K[=T� 6Q���y����&�H�\�;���x߁�қ n&!%ӥq��Z�M���Z0/Z�;��UC�57�����*Ѕ]�$!�9��@θ�#�ԐY4\�}�?�գ9^�H��R˯D��~V���|Փ��K�L�������Y����,���ڧ�:�a�>�C@��=]F�Es���m�%T�œ�f/���E���"�IwJ5����(\�ҋ �v�]-Y�:as��ǡ��Q�'J��!��fqI]z�օ04���>�ʚPCCf1h��X�$�Q؃�1fn�u��Ycj����|��p�8h+^��}3�9�,+o����M�h��Җ�U�ز�;\pM���f��������H�c�bXU$S��#��7��G�d��j��AM�]�����LW�5$�9��⤴��P�I��q;-�]NZ+�&�� -�Po+�a�2TJ��̣�(���ϖ���#���H��?�\�,Q�Kf�C4Bp�f��on)�/�+= ����Wn�[[�)��o&4S�}�b�#�Im���5��י�i�Zd¤�Y%2O�����@$�%�&���>8��\}��T�rmGIh����Oھ/���,���t�OK�[D�҂6��@<�܌RRf�<���!dW�k���fS�t��i��J�	Kݡ�UQ�,R�sȓ������t<�����)���X�Z�01���6$4d�Ҕ�� ��i�OD�
c����Kr��f9N(�W�4�:���y\�t)d,<��!���d�&$�ܽ�ͺ�V�.�C�v7��8��;K��N�.E���mn��Z��;�~�T�p��������2���n�T�"!��ں���7I-��]w~����~����!�e1�e"�S�Ǆ�Z�/����)��ӂ��޵wǺ�<�Vο����v���c!�L=l7��4��4����b׃7�޹��H�����<w��+*���Z?��J�17������l,9*����ޥ�,��ٶꪙ[�A�鍂'�r#��/ش�P�tߍP�frFd��K� Ҭ��	�p�I=�K�^�����%7y̛2T�la�J������y� �g��l��
�\����̹|d�����iis@R�;'�e�{Ka���щ�%�a�^�N�-u~�K��.�[pZІ4ٴ�"d�#�c,x�Fs�����8�ⶐ{�f�iwG9BA�. ,�/"82�<~�e.�y!�v-
�� �3���;��2��63��91SS�ƙ�j�P�+���w�j���V��i�)�Ԇ���d�.�whOkO�e<�F���ƐѴ�nO�VG���j��o�w�|B�qS����z�ޜX��D)��j��AA��h6_�����Z]�ik��*��G��Gy}[;%2L]����JTE,T���{�AK޹{���ͫ�~��ybܲ}ؠ��������o��^V�z��e�2Ng�'d�@s���~Ot;)b��;Ś��l�G����u��!�s9�_�{������8h�.E�ML�dN����)ɽ��,� 0w��J�G�"c�n�A���u%�� S�	L5h�n|��6�X���u���*�=�7V��k9��[B��^a,ڪ�6V�%���㹤m~��7����"��U'[��?�\�:���/�;5"���{�|��׋B���Qo�HPb4��`xx�+FF��c�Wa0�8�j�O���Gd�~ں�ObN��%�7�3�@;%g`��8����DQ�9J�^��Vt�T*�訣��1::
�wx+W,�={�0���d����TE?ج�e�벧�;�, �3��ں���0:{]������d�i3p��-�D���4yʑ���C9��믿��s�=~��_�7<2�.���fu�Bu�?+�8��ֈ+V�{Uq���Q�f�hm?LpG7�͖5fK].�,���`�^.t�!S�W��`����I�C{�[2� ����(�$���8L�^�l�-��r�E�y�k8Zk��{�n(Kp�q��֭[�\�x����s�B
n�+2rsҿ{ȓt� �'=�W��|Ԋ�{N}�a珎57|���_;��yǜ�zś6n����n{���^�쿜М5�߱�K[��:�����ڇ>?0P���α��u?���o>�䃟��_}�c{~x�]���3�{����e���M����\�ƿ�?{Ȓ���?鰷�n�u�-�=�h���F���<Ֆ1��H`q�(�)2v�򕯼��G�Bdw�q����h�<�P��a�!�`dddC��؀�i��g�s_���֍���������J�{�����G���F���b�|�׾q��u/xN$�/�ع��������a���W������ǎ��q��vͭ\y�.~�Q�լ4��ܷ��η��*[���g��s '�~�_�@���+���u�\��D�m�����y��8:�w��7exd�����k�<��C�c�8��c���/��4B���?Ж�я~֬Y�ۆdΜ9Z��8 �����vo+R�n�[��1ZD�{�9&'������W����Dpص}��/DSSD�����b}j�T���#��w֡0ը����U���8�)�+w�#��(�\2.��:��?��2�k��)�h� ��wТ%��K>�����b�RW]u�FƧ?�i�3.��Bx�ᇓkr�E�X�����U���Bt�s#�{L�ϰ0�'^hDh�I�:E���)Vk�a�y�h��LYc��FB���X{�p�I�Z�����=X?�:q�ޜR��%�p�m�mp�%�����I'���x�0����������)�T�r,ɨ=C$�y�۪����4F�M��%�Tg�u�X@/P��i	6R�6Z��\�'i]A~@��C��E7�V�5�8��P��#��(',H�SM�TfL�vG�T[�X��Q 9]�:�ٞ�{fWK"�Řy���݅ju����`���!�nxD|8S��t��lH]f�+BK�Iv�L�t��I,;��@�BkR����G�r�ǚ�R���`�ڬ!��B�'n�'k	؄�����C�,h]D:�Ecf�l��i�|��q�2v��#��M��S]s��}4VB�|��q��l�YC���:�D0��3���a�j�X2�b]K�y�,BtV�7�e.4�fbS�Y�!#L�S�?jE���\��f!hX4>�\i3gѵ��]-a��H��(����i���9��R�RPi�yI���5��ȕ�3m��4��#Y��b/ָ�1�9���$�g�N�$-A+d޼#�]��ˤg0�Y���ٕDbH�f�[:�bo�B:�ǖ��u�̲�e�P�
�uΦC�dw"��ĥ�d_�gz�:�q(Oc�5�HS@�����HS��l��#fD1cT���y���ܹBkqO6K@�6=S1Ͷ��3�L]!8���c���%0`~gv�5��䀔�"��s��>���!����>{
^�?X�UM=����.C�N�cu�2��d����/6��_C� �����Kh(q��a��<�GO���O�E�$om���/���6M�?���<�Z�;*�b9	�߿C�ɶYe�N�N6@�Z��a��btD��2���i�`+�d�"�i�-T��ɦ�M���F���2�@��!��0[m��:t���h�璳�@iiW�[gVV���l�����5J���h���y:��El9��T�q��Um iʴ�L�Jdv�v1!�@&Z-_��Ԑ��2�2֬"��Ͱ�\���6�N�bm�P�?�|ZK3ݽ"��%��#�,�,�����"X���X�6�`c�5�w��Do>�Ѩ�� ?�gv��yRd+��>��U��\G�+1s:���fQ1t5B!c��v�s'�/N��B胭�ۦ�gTrH�"d�y�=�G�	@���)e���d�Mh�V�H��2~zҾ}�9j fz���L�h�\%$����j�+ee�5��6��r%'s�$Sfٔ�qgf?���Jo��t���0[fܖv����$��io��B���e�8�Ikꌚ�>I�;��z�L	B���3��R��:�0�/SCy	�Xի��L��DQ��6�I<�m�#`f�)K�ȥ�@���%�0+�鍃u�3qm@�7����G`Ȃٶe���B7��x;������B�����Y��%cq�q�ˤ�S�]9:1{�۬!Ĕ" �!rK�Ȍ��3b,���>�T(��y�W�6�����r'*���$c����=�� ����"�Ӿ͆�h6��:�E�&���kt<SWH��gJH
�+�v!����eu��2���;�(��<����f̘CA�����lER�S�T~��6�*c��"���q�l�>���j�?�V���~YIK����FX7�H���G��f�d���LJ�۔9�������@`*3'�И+"�鋛�{lx�WI�B�Z.e��vߔg��.E��d�Nj��R�Ξ��vg�6R���	�r�� ��C���7"iR�(d��q��*�gd\������H9+�����lm �Y�+� �ƤTo�lL�fepa�i] D�O����La<.m�BYo��+d��'��V�Uk�2d-�.��2��Hx4�1eR���%���ȴhNZ�9�S���A��h�\uf���
�Z�R�1�qH��]8�j��1w���2���������5<���Ӓs��l��7.JS��5+D�t:[7�� �3��H{�{�|��NJ�h3ɵ<�{EE�&�`�z��y��)^�����fOS�@k,%��l9"\	c���W�i[�)��E�P�ᦘE@eL�,
��uc9&uDU+}�èm���b�%B�h:���H��aK*��QO����y�0��a��P0U�f����Z��̢_=<'?wyK�<�G���V-�T��CN�T����W{^�{�!ԛ�����Zp��qb�kN<�d�;P	�����*�秬z߻�s!fn1�OT'�Q�Q��̿6o��z���YAHOO7���(t���B9���nX����|b��_��o,��%r��#��]�}����H�@����q���>��E<R8��ǭ|�V�;�y+ja�׽�g���J��%`��ms���/-�������u�W�^������*�u����ɯ�>�E�����F�j���۷kN�5'լ dx�(���������0z�?~��f�cs�R�g�|蟾����e�?����{�E�4t�"%����v�H3���}�1��+�`�K_>zч��/�H~��;��/�e~#�?a��[����)���o��[Y���;��F�_˔q��ö����w1w6ڬ �6`��N?���:�~�D��񩈬���j[�tWU�y��G���W��澡��Zy�k4������$e�G��L@��H}(4�z�}�4��jm��������YAW�!x$&x�%�L�;����<��䒳�_�rYhi����ڬ9��5ƌ���g��
B�EX�����"WϬ�T
�<�Ǥ5v��@�?����2[��BH[B�I��Tk�k�B��r�Ob��6�KdV���{�+RfuP������lO�?:��D� �	��>��'sl�ڬ2u4O<�Yς�+W�5�\�+5p^�����n�M_���3�<��^شi�>�t�R8�S�}Xfۉ'��ݯ?����o�^�*صk�]�V���W��p�M7��А>�j�*8��#��k���J@�f�dI�駟�]w�F6�a�HpA��җ���ߟ d�ܹ�X���?\#�!��H{��G�`�3�8��!�/�c����L�m�$��ں:]ө�N�dIS�z�IY�"a7n�믿>G*~���0��?�)l߾=9�w�^��ꫡ�H�"����w�N~#�o��f,�C�ӏ~���1�[�+��qw觱�^�;F*�oذA�e�wܑ\�}F|w��������yL��u7�pC������>w����HI{f�������dHғmO��#щfIS� �eKr|��3P��8�(���޽֖�#"�ZE\�o�]4M�y����$��ϧA���lN�����N�ά S5��7�ٴ5��0"�d"h0)fk��H����rćXF@,�d�	]x���u�&b��c���ȌsH�O���G0Ԝ����
V�.E.�J�H�P��a5x�����e`i�a����
�Ϧ

�;���Ԛ[&�$�A���#T?��1,��V�*���Co�T_1��1�S���Ȩ>�#��(��T�U ���҅����:�.�(*���ݫVѸ�Ru�GPR��L��|Z�9"�
ju<� 9W]�cx���}����X������=u��B����y��σ�h�q��aJ�Y�-&?KG�
�c��4t�d
���t6��$����
	�@�t�yL��z�����	�ޙ��y�:�MW���꿩�Q�qOwܳ]BWPP�E��z"L��c�&��z3��>�C�YAH9(B/��uw}f�,	���˾2�#j�nW��@�c٣ �C���`B�[��Ľ�g>)+�6�WS���P��zB��/�a�+��ȥDnQ�*�##�wI�&���O�d\]Q*�{��Yپg�-X�v̷v�ZU_��SQ���6�ݯ9�ս=�^3>�f줚��j����]K~��ڨ����!'�Կ�λ��틼X�}�E/�t�z�Ԩ��|�|�wѩ����r���EjլQ_���u��v���G�8�z�=~��Z�7#���� 3�0Na��h    IEND�B`�PK
     $s�[�����  �  /   images/879f6d20-9391-47d7-8a0d-9140b0e14aa9.png�PNG

   IHDR  �  |   \ˑ�   	pHYs  .�  .����'   tEXtSoftware www.inkscape.org��<    IDATx���y�[�}'��}x������"nZm�v���'q�x��ٱg4�EQ��g�$�}�9}fڭ�e)+���OO�9�L2q����[�M�%Y�(���Q@P؁�����AJ�d.U$P ���sJ�E<�X(������R���������K�wDDDDDDDĀNDDDDDD4Љ������ :� `@'"""""" �DDDDDDD��������h 0� t""""""���NDDDDDD4 Љ������ :� `@'"""""" �DDDDDDD��������h 0� t""""""���NDDDDDD4 Љ������ :� `@'"""""" �DDDDDDD��������h 0� t""""""���NDDDDDD4 Љ������ :� `@'"""""" �DDDDDDD��������h 0� t""""""���NDDDDDD4 Љ������ :� `@'"""""" �DDDDDDD��������h ��] Ѡ8y��l�E�TUm��n��h��u�� ����������hS=��#I)��N�3�(ʘ�r�_Q����eY!�uY�
�e 礔g���^x��ܩ�Љ����h[����)�x�eYw�l�	����l��_^!�C��l6���,�B��ѥ�M�4k�a�(�Z�U)�㊢���j�賟�l���� t"""""ڲN�<io�Z?/���ݾ��r�;�Τ�iA��������	��UU_q���a�0�Z-��u�j54��ngu]_j6��B�o����>�O,�����NDDDDD[ΩS��\.�v)���n�~�˵��r�����z�B�����m�J%����R��Z�օF�q�4�oY���<�@����	t"""""�R���/ܭ(�G\.�~�ǳ���F��$���M��i4XYY���j��l���jg:��W ����߯w}@ڲЉ����hK8v�ؘ�(��lo�^o"�J!o����cii	�B�U��N7�	!��ﾳ�R =t"""""j����|.��7TU}������L��i%��d��z��:fffP�T����i~�ȑ#_��Bh�0��P:uꔚ�fߩ(ʇ=�-��@,s��i�����&������|smm��v�/
���|��ka4�Љ����h�LOO�
�cN����w0FGG�r��]�+�E��̘�r�������v�����:��~8e��>���}>�>��7��d���}=j�Ο?/���~�h4�R(�=g��Jl�.�������z>��ϻ4M{��n������zw%�I5�Ll0���Ů]�Ĺs�� ��m!�C����*�DDDDD4������j����v�x<���3��@Ӵ~׶nn��v�gϞ����4���g ��w]4X�ĝ�������������n�����L&�����nX�\�ٳg[�B�[�i��#G����5��`@'""""���/})�l6�f������x<c�T
�Xl����G6����l�X,�7Mӎ�{��~�D��K܉����h �:uJ�f�����{�޽^���D"aO$�ٶNtI�R�V��v�}{�Z�= ��&�A'""""��;~�� ����:��z��aO&�����wi=�j���3�t���?����������5Q�m��������h�?~|��������|�����@�K�)�Ӊt:��q�P(���Ivu't"""""�t����|n�����������z�;�ɤ���[b��z$�I����������� �A�k��b@'""""�Ms��)5�˽��v�r���XLK��[j��z!�J��h4��Z��}��t"""��t��)uaa!�iژ�2 "��I)=/�F�B� �!r��_��g>� �o�h�8v�؝��|��p�����A���(\.W�K�)%�z�)�r��7M��Ç?���GTDDDD]��/~1dY�]�e�&�8�r�bv��o��������B{��RJCJ�w:�F��i���6==�*�x��].׏>������z��G1��4M{���;�����L�`�ߥ���H�ju�\.� �6�t"""�u:z���B�]Q�׺��M�v�=�p8�.�.���AUU��v!��t ��ah���u�z�v�eFA�����Y�4O����X,��|��~?^����CyǇE��Ϸ��v�L�RJ2��}�RJ4�M� p8p�\=���j�駟����_K)?r����=�:���Gy��e}��pp����e�����#��QP���Z��T*�R�X��/7�󺮟�7��}��{�5��p�z��ѣJ8~��<��׻?�8��44M���I��F>����*èZ�U�,K�l6��i�p8,�DOó�>�l6�]]�?}�}�=��h(0�]��?|���q:��y��[�nw"�!w�M�i�(�X]]E�V+���3�f���>��<~��űc�(��1��y���9�����x<׿��J�fff�z�~�V��7MsNQ� ��rLU�I�ǳ����WB�PW�_XX�����R�#G�����9t"""�+����!~�f�����t���T*�h4�ӥ�RJ��e,--�Z��V*���v�ۊ�����
=��&=��q�0>b���������L&�A8��� P,q�f�\�����V��>��O����\>��7�v�ۂ���w�����]��Z���g�]+
��}���@�
:ѫLOO�Vq�������K&��T*��!CJ���U,..Z�j�l�Z}ܲ�G����A�G�uF"��	!������\�ݩTJM$PU���]W��ę3gڅB��v�?>�����b������l�F�ѷ�۷��t:�RG���O<a����h��!noٞ�~@DDD4@ĉ'~�f��Q$��d2yh����t:��3�B�b1�߿_I�R{���5M��Ǐ����H��bzz�͡P����T,{w:�����j:��p 333��j����#G����m'9|��)�4�Z���,,,t�UU�r�����t:�]�c*<f�����ɓ'��v�_9��w�|��f2g*��wY���عs'�^oH��J�⚞�N�:u�;�S�<��#S����4�n��{(D2�|>_�Kېz��j�Z���O�����{��i_���o,��{t]w�H��+q:����z�>
�BW
gЉ��h�;u�f����_��?�{���/B �Lb׮]�p8�F�������O=z���hS}�_?~�~ �B�߈��oٹsgd�޽C��\.��n�K)���O������޲��v���V�]��n�CQ�"е;���t"""��.Ϝ������P(t׮]�����wYW�k�.�ܹsw��H�Bc�w굓'O�u]�eEQ>������=�x�>LKٯ��h�0�����^��tΛ�Yn6�][�~9�kR������������5]��'����P(t��ݻ����wI���z_���Eczzz�_��.ںN�8q�eYq�ݷy�ރ�Pț�dЭ�h�$����#�ll�Z�ͦK)���DUU!�R��>��z��������Ǐ���i���p�"�׋��Iղ��WVV'N��x�}�=��hk9v�ؘ�(��lo���^o"�� �:��UU��� ��<�(��f�^�zq1���V�
:mK�<�Ȕ��P螉�	��3\V�`�T�e����b�S?��O}�S�~�E��s�����t~XU������n�{2�N+�x|��3�(��M��B����F��,�6�����)���y�DDD��:uJ�,�H(�#����p�K�!�t�Z-�n�o�T*���&^�N�R���;�n���^��۽/�i###��,� 	�p�\#�Z��'N��c�+QN�8q��n��t:#~��k�X�  ���M��'m;�\�n��n�ߟ�d2�.禌�����ޢi�;���_��zh8MOOߺ���ǚ��A4��d2y��������-��f�!�L*>��6 �}���u_�җe}���J$���
��6,�j
!�]�S*[�������
N�<B����;8>>E��
�Ӊt:��~[�X���'O>q��r�����N)��QM�����z��t&�A0����z�R	�ZRJ!�t:���7\{"�@�\�����J�����/�����߿�����;��	o��D"ѵ�\
�i6-�Z����`@'""�m��n�����B.����r�"�cuu5�l6ok4������ѣG��h��m6ۯ��n�{*�H��Tj����똝�E�\n�>�n���e��6����4-��x"ccc�nf'��Ν;!�ܥ���\.�LOOG�C˲�v i �����@ p{0�LMMu���j�4͚�(���1t"""�6}�Ѹ��ow�ݻ��t���!FGGQ��6�������?�i.��+ǎ{[$�-��}����D"Α�h���ڮ�R�����j��L�^ڲ�B<%�\�,ˣ��.)�[��m�v����w2�\�}�l6�ڵKKK���%Z���v���aԅ��fs;������b���Ѯ�s�0�j��4�Db��wNC�������N��n��3
��[�������]��W�����~�D�����{|��r���zo�L&�aXI�h4p���N�P����_UU�����U7{�ԩS����k�a|̲�7��vo$Y���btt�x\+�;j��]�!������A4��n��ĥe��Ng��|���M1�Ѷp��)MJ�v�˵#������d2(��{���;N�8����l�k��;q�DDJ��6���^�����K�ӈF��.m]�����E�Ry��n�Ց#G������/y�Z�T��������Ս�j�ÁT*խ�׭R��0� �m��40��+
�:����Ǆ���Ì�p:�H$v�׻߲��u��4�S�Niǎ����>����h����c����p �R	�J�X��/
r�p�r���'�nƷ��L>�ߌ2oZ�\F���
!�w-�?�DDD�-H)�q:��`0��Rz*�L����9��;v�M��������o��r�^��3�X�=�Tj��}�l�x����Z�֌�o|���.��z�~�X�v�Z�f�b���Ç�������$"""�G�U��𝚦�B�POǒR�R��\.��h@J	EQ�r�
����z:��fC*��f�P����/��?��G?��PCC���� >n��_����|����Ⱥ;��F��v�]B<���>����tN�u�0G���w���
t]�������������@ 0f�ۓN�����p�Z���h4�f�9o��eY!�]Ӵ���������������h4����H��<T�����l0'O�������������z'�鴈F�}l�z��4����+�T
!V-�jr@7kkkf�^�hY���]�:my���v8�^�╕�����j��Z����(���������j�B���h��h4nݱc��W��Bd2�j��f�}_������[�ѣGm�H��������{<���XLK��C���j�B��@@��ȵ�eم� H����l6祔?��)m��Z"""�kPe��n�*��J%���6���w;�Ο;���r����ٓG��K)�G�� �7�ٳ�ѫ�u>��H��j��W*���z2�ͱc���ÿ�t:o��|���ott.��ߥu����n�K)w x|��=z��D�B����a�7��ncyy�S�՞3M��]�:myRʄ�(�^,o7M����\.��4��x��ῼ�m/7�����i�R��.^����l	r&����ڮF���ǎ�ڑ#G���@��}���4?�i�}>�A�ϗ�d2ت�~?
�B��j��H�.�+���E��؋��h6��:��7x����]��`>S�����+�(�[Ӵ�����
������߻����5V,�s����F��+
]��E��!�J�~���(;z�(����z�3==��N�s����N4����������l8�X,��9a���2==�o=�<��#^!�ox<�ݑH��%ސR�����F�R9c����|�&""�� �(��}mm�fs�_����>hv:��i4��ֺ^��%�I�����3����QO=zT���~���|�������5::����J*��&p�N�Bsss8w�Ν;���y�El�Q��nG2��������}�GF�u��z�cY����z_�M���ܜ�T*?B��>��l�k���%�DDD��	 6!���e��e��hX��5M��F��t:O�^���R�,d)��L&�V�u��j��C=���~����F]w�ر�H�cN��N��s(GGG{z
�͒R"��cyyY6��a�N�S�R�f�yG��t��鴈�b��t:�Z����r�윞��s���w/?B��ѣJ(���t~����.���üaRJ\�x�j�����T(���hp0�іv��I��R��l��:����]ӧ?�����t���X���p8�@ l�Z |�������=��q�0>b���������L&�A8�s�Ҭ���籶��Z.��0M�	!�,��iS�u����j�n�V������>&!v�ލ�/��l�_��j��z�7�?~@EJ�D"S�c�������I�b��͚��G�P�W*�t:�/<���V�k����NDDD[��늢(=	5��W�Rn8�<y�.�Ppi����E�^��h4��裏~����b�ǥ�;z��3��O�@ ���r�N�Rj"�����.�8�<
������wE9q���~����_;v���b�>)�[ �w��q��B`ǎ�þ\.wO�Z��4͒��B(6�-�t:]�x�Xl ?��f���r�r��} ��Ǫѫ��G������z����<��c��x<{�DW�9+����U[��X��������sϺ����ߟ���
�v&���t5����n�t]W��r��w��Һ	!D$y��������`0��D"�ڵk�1�]�_nyy����R��w����'>�v%����{�'t]�-�u�\���t:�F���`0�	�B�X,��d2�t:��3��|aa�V,����<|�����]��DDD�1B��] ��N n�/@Qo����������� (���{�[���;�n/y�p��x��׿������̭��w��&�޾���o����u���i��8}�4~���j����.\�h��3��� �M)��b�:�Z�b����������T��s?����ĸo�IO2��e2�|��,㦘����z
?��?���o���8;׺�U�m���]�5w����7���fI)��������ǟ4���j={�܆�ļJ���$\��JfB5��o�R���M��+�P�Pֽ�DvK�(H�u�2�*�\�^-��%�DDD]&�P���h��Fv����SCB@؝���\Bqt�� �D������|W�ۤQ�,>t�P�? ��A7:h��]ߓ��O��;�s�S��ݵF���}NL�r�$��hW�M�022����x_��xs�Ӱ�͝����,ՖfV�
i]���2���FvCq��2�:����^���\N;�ܓ�-�1�K`l$�t:�h4:tAumm������v9Ƨ^y��?.�Ȏ��
�M�\+��ht�a�&.\����9�����;O7��[���[�]�Uu֞�#9��2w����f�*0�Ͻ�u������jU�p��m�:Q	!����6r�-�=����%u�4u�K�B��w)We�=+����jp�+���h���&�^oW���|I%p�5�o�Uм�ܘ�!��{$n��#�L��vw���I$Y]���6�8��������
��T�ˎ�
M�jW�^}��<S�{���y��KLKL&ݘHz�J&�J�`����z��bC`I�cr׆��K内z���z�\���,�ϯ�E|�F��~    IDAT�5̝�;��w@I����J�
�.�k���km��k���wX���]B�wI);���j�����h 	!���'���k�����Md�/������@�?�x���-�ֺV�n���Z�:���V�sk���f�)�����2��1v�F�YK�_N�L&�b��|���U�1�JWd֯�[K��p��e�ў�&��
��_�=v`�+���p����]i��0FGG�ptw��f�u��RSb�+�km�V��
���4M,,,`q)�ggVpn����µ�ס_�dǀ:��~��}�wx���z��o=
��wIW�7DDD]�8��:���.��M�i�3�x���� JM��0P��zR��f��ݻ��*B�5$C5�����	8l@�$�L&=Ȥ�����[�`0�d,��d�L���ޗ:n�� ;׮Y�{�L�	�i�=��/|���InR��tw�I�)�	"�#�� ���nB@ Pn`i��&e�	��XYY���f��pv����W��|֋�����;�:�WP������8v��mdO�W��~�s%|ADD�B�Q58�.m��B�����	�~��⹪@�f�Z��4͞,#��lسg"�U$�y�+u�Z&̎�M����H$�}�c��d�V�`������rc��bB(���5�	G��vͧ���}���nu�M�84"qKR`Gʃф#���xߟ��p8�u�v�X�l�q\.�N��n	�T*���G6��s�E������*J�+l!��5�h>���ns���=�� ���Z��������ێ�oڼn_�Y|����m������J��p8ܳz��(��(Z�Z���B����n���n��d��:�(��3]l��s�3�Ns�{e��+�s�ԗQ���������.@�f�"�]q�Ci����IR�8FFF�v�����~ăNLśx>����bW�L��]��Z���/���f��x�B�+�~��F8���.Ch[cŰP��B���u\��{u ""�as��-��;��i�dPT���w�$�/�P,{�_�t:~F0�N�X,bi���e�;Ui3�<	Ȏ���m�'	�DF�"j���p���2]�-闸s�ڰ+�C*B&��􆀛)"�c"���TO-�o�֌�HԅP�?�?//��t��f�]�afi3�
����م&:�<A���Z;51��҇���{lB�����j^�����$dDq��ϰ�F��_�mg��5ŵ2����~��lH�Ә*5�/���f�{��{`�^A���en��P`��7�����o��{�ǿ���JL%TL������dbKC�	!0::�R��R��rSb�x��<�8�Q0��bttx�b���baa��.,�pv��'g���kΚ������zX)]�p��2� ��]˫1�u���^-��k���Fk-�+J�֚X]]E*��qq�!�![�x���i�.ױk�����W`��_�/lN�F�������-\�jhcG��M�8����Ʉ�I�KǦm�`�r>���
��Ԣ���ڝW��5�`Z����[w�cr.��OU�_�V���<�W.�3��5���V+Ɔ��KRϪ�-����@�p2�u��R�=�]Q�;��h.�x<U宄g>��5�ך�]頡�4�����^�Y�Av�{d���?�F�̟Cx�p���uͦLF$n�HLĝؙ�"�bdd����R/~�尫�jؓh"W���
$�. �F�.�L�01>�X,�窯�0�K�<����%�����.���z5t"""�~�U����W��rH���.i ��~$�L��8X0�s�<G �ÏN��N#iu�u����{#��,��� ��>{t�Uo�J�9&1�c׈�X�Lf(�u[*�B @8���R庁�ށ"\A��H8�T*5�3�e!��aqq	s�
f�e<���c}�+��b@'""�m����x��Td�ht`f:[����P��aE�����ߔ=̙Lŵr�^X6Q�s P]�� ��2:�ַ�E���ꊠ��Cw��>�1(��K�pk�e�=I�ұiq��4�Q��rn��w�a�����K�h���7Н쥔X[[���rk��X���&~:������rv0B�3�DDDD���	\�w0�#^���D_�1M�����W�_k�T��nw.��!t#�bt4����N��T�k�Vl�N70��_�O���F���0�K�ޟ�h>xFߌf�Ǩ���'�w��؛88L$ܘL��J%�H$:l���nG0��D�Ѹ�ϼ��%��xr��\�{ŷ�˟w�_M�����S*C�'��P��*b�<O_�h�Z8{�..pa����6�K4ۗ�N�&�U��ʨ��A&���lz2�D�P��J��fW�F(6��4
09`=3����{��b�[�k�Oaj�!��"#��ձ`tm�a`ii	��<f�e��kxf��9}�Ǧ���DDD[��'�:���.��Q����jK�LV"�"�Ǟ={6�۶a8{�,N����*~tNG����l��|��΄�ZӀّ��l=�@��k�J��t,;0;[�-���P4/���f�C���L��{2�t*�L&�}G����R"��ay9���K癟��8��F۔��,�4V�Y=��A6ƪ-�=�.��䀆s������A�vؓ� ͋�.������㧗&#-�DˈŊ�D"].�������|O�T��g��a)��4�ljn��@ n��'uE�Q$�OTqˈ��s��>��	{h�z��*����aíS1음`�Xc�FFF�F�ձi[]�\����+��3�Y���Y���i�̅hæT6e����8��H���1�FDD��m�Iƫ
\����U�����3����5:�O��*B�E�B!(�<S�f5�M,�Wqa���k�k�z������2b�e�ر�'��t�Z���Zr��V{��<�K��y�˫0!�g<�C�����09G*�@:��>�-��lbaa��".,�1������J�7��G����M��b4g@'"""$�Wv��Dk�-/oڱk�b�B�Ɔ�v���tŵ5LXV�>P�z�H&��(�q넁�??�Ǯ]�b����Y�G2(p��&G�H"��!���1`�1�N���X��1�\�\���t�ϙ�g��p����h�H ?�H��7�صz��rMGvmc����b��Z��F���3�3���5,�x!k"_�c׮.��pہ[0�#��"��U�q�6)%
�����b���ygM����̉6�����;�oH��rR�¡��-9�0�j�7�t��[Ѝ��Ae�B�4��)�(5p���o<��RAƮ�G5��0�`4��H:�D"�}�[H�R���}�|i9����J��]A[gЉ���:y)���{��'��HG
��b��|=OQ(���l���(B�M	��D�U��k�o�|n��]�����I/v��JđN�a���]u�����0��`a��g�&�����n�@��f@'""�0����JP���3K��0.���{��4 ;x\v���F����Nۦ����*2��U�X)�[5a�J��_���ŝ�5D"���(<O�K�.�,�l��2��U��kx!������\z������!��5:Qwp}ȝY��������"��l,�χh����}C���р~���g��\8F2�x����&����q��[��J:�3D*@&3�p8���[H�P���"�+�檘Y1�l���>����+���ĝ���h��KK��*"�%�B����D��x1+c4j`~��!]�mƒ~�b�M�/�V�T�+�q!g��������h�%�a"��xҏt:�D"UU�]uI�^���<r�%\�V�Xh�̒�b]n��i4,Љ���8�w�[�L��bb$_C$��L&ӓqE����V��44u����׎+x�S#�&CH$=��j<��&�u�Z4�϶6u�����qh̎�;G�H&.ugߌ.��9øtlZ~s�U,�6q6'1_�`��4���NDD��IH9���i��Ȅ�H\>v�W{���(�F�0L6e��t��?��;�Wqۄ�]#��Ν;zv�����i�E�X��es�G�m��W��L$��ʄ����dz���6������./c1_�|��+������D�ĀNDDD�2�:�_k`)�#
bjj�'�!099	���ӎX����M�V:���*����K�1�aǎI����s=��a$��T��|�@�db�&)]���1��L�0� �N#�r��R*�.-g/T1�\�B�����k�@}�%�v����rw��d��(�Z�f=���~��+��a�����]ݐ�*t3F�����w"�ZD<^�����XB���!"΢T������M�Tn���h�drS�M[��N��4a�&Àa�t:P�;޸��l���.QiZ���r��ͥ*���F5L�|O�J&�J�z�C�6_������k�Y�b���s9`�ΘӍb@߈N�sg<��f�ՏOUof�ͮwP�~����F�������]~��U �|ÅQ�(B2��h����u�n,����៟Ǿ}�z���������04��m(�����ճ�u]G��x��l��lB�W6�z��6M���Li��X�e��H��hK��RE��ճ����p븆�;3A$����nZ�{�=�4�����\��W�8�"0[[c��@F��`p��l@��t%$��ʉhK�<1g�96�k߁͗��?�\��ۈ+���Ҙ�n�#���M�D�RA�TB�\���/����
UUa��`�٠��+~9�N���qiɻeY�X�i�0;��R��rY�ܲ��Z禗��
n��0�pbg&���}�����%����
�����R��JW-�_U��2�̷ăJ
����:o�0�9l���h����-U�t�|�=� XX(��_�#��"���v�����J%��ut:X�)�K���N�N��c�K饔0�V�V�F�z�VF�@4`a<n��qu]b���s�fW�ͮk6����=#�	 �`$�B<���-�R�\�g^�l��욅�r@����i������y���x7;�0�k�Y �>��V��ٖ2ab���L�" �%�5�V;�j/-all��U��eY(�J/�N��������������xBh�M�^�__J�f��J�r��
�m �`w�D�ea����/�Q�^��G����}�I/&���q����&te�VX^)��V+m�_U��*��Y�5��Da@�a
���7{L!�K_�1��\;l�"��yN~�O�o�H���K���T\}yD�ѾuQ_�v��\.����˺4=�����x65�
!�v��v��L&!�D�TB�XD�\F��F�gbwRE�l᧳�fMȗ�oNTܱÁ��S� ��02��@hc:���,��..�0�o��"Pm۠
�����������6Lcn�p�PN�e�]�R�t�4T�	Gx�o�4��o���
.`���;d�FZ��0M�eA�4D"�B��9�E�P(�P(�RX��r�T*�y��mx��~:k�|�ġq;�/�3 �� 
��aP���baq�.dkx>'���FȄ�o��.}
8�Ϯ-Ї)t���0�͎��5C9��ޣ&h�d�*��g^�w~%+ku<�ZC�c!-"/!nb�Wg�&��,���a\n����^����7/�V���(
��{�x�n���0ҩR��@?ژZ�vi��jg���7�y����=�n�w@e`��l@_ZZ����5o3LAw�B�����l4]�f���	m!��n�w�ߣ���[8RwAخ|,WS7��+ò$��o#,!\@ ��k�eY��rXXX�i��t:�z����C����tbbb����f����h4�
������w��n�/�3�p~���|O.\,��K�I�n`���+MFS�☽�n;�IDD����=�1�O]�6RJ�,_:k�����F�%D�9$���,�%�z.\@�VC�Ӂ��F"�����K=ݤ�*2���4VVVP,Q�T��3� �a||�M�ԋ*-..a~����:�d�g�
�N����M�nʰ�*]�y���l��3�?������n	�e�o'�X?��z������I2삲���ލ��GˮT�h/�KO�HK�/���{���XXX���:�E����+��o�� �H �!��cuu����;w�ܒ�y++�J���Gv����U��w�9��>������|t@�P�1�aӡH����BJ�X�W��H)�u�[_�w]D7EB�O�pp�UK߁����^�F��r��3�=W2q!�#+#^���D����V�����h4�,�`�T
���υV�d�`���h4x�g�J�066����k6������J	���]5���@�����0���vr�0�0�:lcn1w
!���Y�Ѫ~"��_B4xq)���K:��"{����-���R���:��2��D�Qx��UzI.����Lӄ�n���ؖXξN�SSS���XYYA6�E�\ƞ={�t:�]�ʋ��.�vq���Kg�
,�N� ��{�{f�B�v�u���P�R~bի%�GŇ�l����w����Ý���)�o�/�Po^�e�֒xn��d��``{���I�RJ\�x�|�i"o�N�B$	�|>,,,�V��駟ƞ={����]��svee�KY��8�T����E����^�{лj�B���u�i�m�WW+�WjGůM<([�.�h��·��W�,ՠ�v\�����J����|�:ұ5�bD"����n�q��YT�UX��t:�p8��1����������P�����b||�D�ߥmk�jsssȮTpn���+<>����weDW~ӆ-Tm�1���as�{�����3�4l������Z�:`[������,,��Y�\�<=�_:v-��@ е��F�=�Z�E���Ķ[�~=��`||�l�b/^����wi�N�������"^X�b&��O�ָ����k�~���a
Uۡ��2f�jU�K�
���W]~�H��*_���-k5sT��!��� x�`�;� ����+�y�i�XY�t߅���&F�eD�y��雮��h�̙3�uN��Ǌ]��t����X\\�i�����䛠�鼴�|f���|�,g�t�~WGt�M�n�F_\�) r���nP����ۆC�@� W��fH���t>Ȃ^lٿ�<{~e�҆�SJ���m�BeD�Y���jX��rm]��v�1>>�.���D�ifgg��� ����Cz�E���ca���K5<��xb^��6�4$H��[�U_qC/�/^w3�n�1�Qk?Ƽ��aL!m�,cv�3p���٢����1k,� ���ʳܥj����S�V;xa����
���n����s���p�A>����,��˘���wI[R�Zř3g�����g���3|�4���4d���9`z�Z�i�t�j�.cj�6�M`�}⿮����_qT����i�1�(�G�}��?{w�XZ�	��<w��$K��ջ]v�U��4;t:@X��$���LH&94L�=��I&�p��$Lff���IB �a�4t�+]U][��ʻ,/��ow{�?\UTwɻ�����S� ˿��m��ճAIܽ�פw�1�fNO���) ћA$A0���+���p044�G�������������"!|Mz������E,.�b*]��rg(����)�T���u�G�|D�����n}�^��ꚬC�v$��m���ū�F<������r��h�SK���k��c���2\ZP1��a~~l?������7����0��188�4�J����duK�vc�������sx�B߾P�W���9�Y�͖?��Aw�(�]j:��N����i8�q'#�ݢ��W�����z[�㸝໸[h�z�,@Y{R�6������R*Fb%�G�e2�F��>�1���IT�P�    IDAT�Ux<6޼�۝P(t3��������s�w�1�\.���V
��XµUߟ�(�+ps��A�{̚�S�SFI�Ⱦ�j:��ɭ�Z�cG�v�&�zH�#��Э�������0�)�=>�/�o�����i�2�C*��a[~=c׮]C>��yd_s�<�p===0���PU�Bj�*�
&''q��9<����Ǘ�7��Λ�C��l��3�A߉N]픚N�u��m�PaV�A$ �:f����t���͖����xBpD�~��Z�i�fW5�,W�+ �Nc```ӯ]\\���* `xx�Ը?n����P��Q�V199�cǎ��[PUKKKXX\��bS�kx��Gq9��3�֍#`9�5�;����)A�z���X�h�X�n`���4��"�/�C:�N|�v�]^��������㕚�B��o!���k9��K�D"�]+�XXX�i���(M쁻��� �^��b�������Zݒ�0ư���Tj�Ky\Mp!����*���,������HZ�.�5	�MŃ.�iE�V��b�0+Y�9�b��x�\�K ��i��xe���f�&��U$#���111��M����t]G8��������a\�v�������-��Xg���J��9\[V�̴�\ż�5B�P�>��2��s��嚌�0+Y�e�՜��%jEe��B�<����t��/L�?
�����m����혀�	�Sj:���>����jvH����w�{�l��L���r3�����d�L�,�U�Vą3:%����JQE&��?�+Pw-���,@�>��p���D�PmI��gUE�HF��^�gggQ�T I�DK�s/�(
��8VVV055�;��й� P��0??���:�,�1�T�3�RY���_�џ������?�ȃ��8���n`�
cm
�򥬺:Ycz�B�S}ά��(( � P  T�c�"�Q���8��G}B���8x@߭N	r��k'�l��C�K53�o���/��H:g�&��h��2W���d��i�1m� ϙ��0�k � ,0� d ! ^ #�������`�I=]]b�H��<B��s�ސs~r��>�^��`YQ��4��*b�9�C�8z�(!(
X^^�i��µQ$A>��LGFF�n��al�g�^��bS��_�q1�����A�B��:���P����M�n���Ԧ_5ss0��f��E O2��{5BH��_x�6���a�x�<toH��G����ħ��E�@^�^�������9סl?����3�_{4cdg�0�/���_�>cL��e �������x�2r�Q�� !�=��=Ay���ͦ|;S�� 2�r���Ї�\��MarQ�h���h��
b��]��0�D���)��DA?�]��t:���ގ:z�1�L&���"��P�䒆g�uT�]�o	2ı��̾�� ��OA�� �M�:�O��W��4�j���;��o�[�� ���]��{����5����=&����mm�t'�N��^���F��+�P a���v,����p�"��Ow�|3�������;V-����1�L���ډ`u��^V9�C#B����3�}tj�C7�i%]Pٿ������3�;UM(l��������L�2�B�dz{���\m���ͪ�w�	/AUU�j5Ȳ�x<���\c�������똚��ɓ';bW�b����9�W����ROOi�V�7�@ÇA|IT.�_x��)z�Is��L�g�֯��:��j�c喔b��3 >C/=�$t�N)'��v��J�MC�c���\'��I5i�hyŠ���꧛��ld���w	�7���`S���W��U�n��� �0,����U��|o.��GWz �V�� ����}U<:w���$�}G�N�c�Qf�
wyaί@~m����=�a~M��R}�,
�A@?i�R<G�P@�R��ʊ�?,���H�RX\Z��T�����qm�hZ�	A>�s�_��z�~	�4Fv��O��*���1k����)�{��
����;JO���{������^��&q��)�״��6ç��\������?Ԟ��q���;��/�^&O��wԑ����C�����g�O_Fi�m �Sm�U�X��@h�ۜVm�ș�9HċX4�wm���x���G$q݆q�a �N#�^��r	W�83�����p�#Ȑ�ڕ��
��ZP��f�z�j��9V+�$clֲV;�D������|w�d\��f���A���$�����\^��5�ѫ5��1���D?��&��	@��\����-�< �P�;���x�����\������/�oQ-	�z�!��~���� ��� 34K�i�$@*\������JMC]�nY�0� Q���޶��6
���z�i����n��2�Ν;������e|�l_x��s-
�7
i��г�P���B�����~bU[x���j�UV��[1����vW���x�z�+�-~�=�9`�.�2�6����9�f#7B9������{���_�C:�t���2�W�����|g�n�>�%����;G'�}�a��U�[ڗ�_�QJC�h�x���� ��		���� ?�&!H$0KKK0��M��J�\�/��s���i<v~_z���Nj����~C(��wB]=u�t{jrmg�X黟�7�+o4j��Y��K1ƖX��Jm�������k07�@�������~���v��N�я��a��C:�2����3��t=�/�SE�o���琉/�%��37ou;{T$��!l�S}�Tk[/^�`,&����s�	�z�PU+++V��g��bjj
g�]����|�L_>[�J��C� ���:���\��s-��^1KO��5����1ն��0ƘQ/��.|���e���x[^����:aݴ5���~��H;�r����D>�>���� (���&���u�q;GE����3���3��?e��Ӊ �6����s��	��	�[�n�c(�� ��醉J�}��O�(~=��X,���9,--!�LZ�ή�����%,.�1�\���"�-�87�C3,ޜ�J�����>"��8�N�_�eF����b����K�^|5c��rE����g��]/}��4��F�|��6>��q#�2��G�[W��v��s!�Y#� ���,�C�K0����ϩ~�.�����O�K��Ƈ��������W����&!�F>^(�msa0��xD�b����v����(�^�#�w�ƣ�\.\�����x���:��f����zD�0�&T������ͳ���z�Ջ�qJ8���6*��-=���[�����5Gtty��<o3|
����9�f�+_�O����N9�����K?�E��_�,9gMz�"��f �>^(�oz�xRD�'��x��Y>vDA8�i����^�Tp��e�9��8��;���~߾��T��u�G %���cV���Y͢���ϳZᵌ�����Ӵo�r��ʧ����	x@߽N�V��<6�C��D>�>G{3���;�Y���9e�gq�8�����M�C�/�?������l���6f3�r�ǋ������=�à�ַ[�F@___����M�033���]�s�Rx��
�v��>�"��`��.�C@]xf�93�[��O�٪Y-��1�����0���42W�X��H���6�-���鄠봚��)�����էa��G�9��ne�����]J�i��2�#�cx���խ�WMC�4�8R�M�Z{v�E �-�#�|���dY���i��d2V��"�1������8s�<vn	�:��?~���K�3.�D�8�&�&���N�=���R��r��p�a֊�]}���[ �����]��tz(��|�tw��߅��߾��d�k����AޘX�{��V�$
bu�?���rUm[/��$(>ŋ@ ж�������.��r9\�xg�]������}
��lO\�PӜu�]�0F~��V�]0��LK�{ި�>au/��3X���s�w�E;�ڌ#��B�5;ed3<�;霓`��x�	�=�>$�6��A/��o�ՋV��)�#�,/A�5���1���xe�����`��oUm��I#�ZW�\������I|��+��S)|���|չ�>q�Ԯ}��6lʆ��(���V���խ4clZ����32l���c�����<^��5iWP恼�vzۋ���8;0M�s���(`Z��:����o ~����z��V�� �G � (���]#�bAY��s�[g?���~T�U��yK�%��t:���fV0����k\�ʀQ/���ieə�>���)�c;����k�k�>�XZ��c�V��
f��_�����}l���SBg'���u�`'!����3��tS}�AU]y;��pT�������V�s�,����wͯ�z[���y(^���s�3�N]]](����rm�1d2�1�Zŵ�e�0��3��7f	�C$a��@����f�^�����E@�,`�_}4k�J���Va�i���f36-f�)�N�NnEM>��=S��T��m;ݝ�l�x�s�w䣯��ퟬn�!���|3��m7!K�~g�tv*�����|ۮɅB�.]�����3S����៾sO�O��%�L��(̲�7�����X�`u+��sO�ah�s�T��`�M2����-l�w�]w�l�M���P�s�O���~�#���:��+�����5�E�[�����z��n��9 ă�$R>z�0^��(B�4�J���RU3338��������k��S3X/4>ҐH
H���B�j�i���6�P��Ⱥ��gc8'r���Bg'�tz(wC�w�ޏ�O� ����սp��˫��|��6^�R
�f!����W��	�B>
Inn<�9G  c�e�0�R)�}��=7��=�Ʒ�����U�d�>Ϝ�
X=ג��I�9m�y���6��� ��6c�lu/���k�_���vO�ʹ#��u���d�2~�ܛ)J?F>���=q\�:#�US���M�{��,�`�<Hh���j�F�{^�B�D�|���s��(
��<*�Jӿ���R�W����bgg5T���Pi��*�������,�7lu7�Kԧ˘��'���9"�;)t�{����>]>'���v\���;O$vM�0�a��c�&�����O���5�$�i%R�3�U�=��{H"���mK=���^/c�V�M���J���H����|�+U��V�Zx��$$l������*�K>������/C�{�խ؃-�E0��t�1��խt:[���k{�䡼�ud�Pc�=��.�
��;nT8Ή�_������n��#��5�q@�ڴA\o�(|�ܡn|�R�T���}��iXXX��JӋyL�K87[����Ʒ��`����1C	05`��v���Q���y@���%�� ��}p6��)A�I57c�Ql;��8���^ �j�i T�����PIi�x�FЃ>
A �x�1���A L�D�V��4�y�
cKKKH/-av1��t/�T\XP��[�3l�M�'Vρ(�?�����Y^���%���S-|��>8��N	�N�و�3��q����#�y�=#V�A������K׷ހ�Y��>����^/j����z.����W�:���J���(Twx�@��-g&�'C-:>� �f� �lu'�u����Q����;%�:id�7��v����8�x�^�c˗�l�EA�r�a�'�+�|��$IB�Z��5�n�V�a~~K+k�����rgf�Hgw7s�l1�1�J0wMM|1��4��խpױZIc��[�砀�)A�I57� �:�q�2@���qAl���l�2OYDa��7>��\��qk�������:�^Z��b3�.,����`��g�l�\����1����Y]��.L0͂�mpl�;%�:�f#n
�vx-����AD[��r���h�s�7��cOIi�|
���p�ΉA clˀ�C&�AjqKyL�r����쌊����7�U@@��M��@��s���(g�(���n�����t�4�߈�������!�-��8n?( �ԬAg�d�&h�m���= �Ϳ�r�u�Õͦ�
����y\Y�bfic�y�҄e���0*jm�ul�H�Ҭ�m���9k�^a��}p\Нt�Ts3v	�n�C�����n8���G
����Vm����o� ���ěS�9gE��z�V����V�pm!���
��U1���T����~�P0-�H�9	�l�ߝS�c�#3T��y���68�*⤠봚��-�ڽ�^�H�D����8�.�Z�X���	"��H�����5��PT�h_ �V�g�;!���74�t��斋�J�qaA��
��{ns�'�.��N��n�
�Z��6��
�N�N�o��A֮u�[�o�q��	��*���@�f#��_x	N{0��1��`"�P(�T*Ji��q�G���:����T��kKu��QQ���T��{ �%�ā�{a`��H9;pD@wR�uR��8!Ⱥ���i��`��8�@��5a�����H�=U���~�e'���/�D"�@.�������a�d2X��pu>���*NO��[�3�uo&@$K{hfj u�kq"z A�Z����}/��SµCy��8���Ğ�m��q�Y��� [�L�M��R���RB�Ѩ��2���F<��� $I�^g#��m:s�k�Z��J��|E�մ��gU̬j�n}xSlw_aj���Pkj ���.�����ku�[���p�C��u�RCU�����|���A��8{���-: lz>4��{h4(��C1/&�H��@ x�׉�B��QVn4M��Hej���:t��-� �͇;�F����L��J��7�k�H
!q���68:�wB(��sqK�uc���F��֚�q�U} ���6`B �dw뽎��<'�$��b$�`�}}ID"�����s��l�a�1�R�]��ݽ35�| ��<hσvA�� `V��mp\@�p��Pޮ:nz-��q�le" � &(�&k�w;�~c����� ����LđL&o��FnLu�u�1~�Ci��1TU������L�qJ S����V��]���鶺n��W��p�Cy��ᡜ�8��0l0z �n B��UJ	J`�۽�2F����q?􇐸�����~�� ���1�4��}i��d(�-�Noq.8!���;֠��*�����	�$BH�1V���Ng��	�|��m�Y^��8���	Ĭn ��:����U����Oqר�1t�?���<�Q��*��ݡTU�n�ȕ��f[tPL�@�Lq�* r`����F��ٹW��{�t��,�z'T'�kʭ����q�nOS��Q�!��lq� ��{��"plЃ#��1�����htO�i�׋j��Z�YvI��0���0�K�ߍ�e���Z����Q���]�9[�b���³�薳m@�)'��V�G�A֞u�Z�*�y���6�WYUhh:B�d6���x�@���"щ��} �A)�����cI|��� I	'�<J0�B"C��F�}>��,j�ڮG�9멪
]ס�Ś��m3�n��<�_&l�!t���%����z���Н����Fx�uo�� �����lR;���x�&�=�n �Ʊ7|&��c@	�b���j*���� �=�=.K?��nw���)�F"ڃ��A(���|��|���^o��<go�j��P�Ll�"�5���wBE�z�F���<ɻ�n�{)*�bB�8c���t2Gt'�kʭ�����:�y!�� �[��q�\���V�qC]�ADL�Ai�Et)w��8��`�/��D�����M�DQBP�՚�=��)�0�J�k3���[��x5 fq��w���y�Ult�g�U1���A Y�K'�}@wR��S�;�����)��[��    IDAT	!�@�����`'_eu7�S���n{L���~��>��0�����X���m�ocՍ����5*���t+֟���_$l��ݱj�������	�?B*����ƶ9��k[�v����Q��� ��p>r����NW/��p�dt/���խ��*� ֳ7�7!@���@��HPA,�D,�����g�7� P�b�J~?���$�j�nb>����ۏ�3�
���F���]V��m�
����g��. ou;��#R������v�l�1v�O+��N;j���nO.p��ܭ�"c���9���3k���n�6��� ]G���1���q?z###-�7tww�R�b���:\s��u�ju���t΂t}�e�^��bO�}`0��!E�[����BD��W§ Y�����١�Av?u�Q�-u���sΉ:�X3��Eā��n�6u)
��q ��x��#�~��ؑ	>|�@{�\�B ����0�l�a"_�`�8 ��|cAB�������3�W ����m��~H��[���}#ŷX�G#��V��V�rd�[�5x(o��sΩ�^%xr����γk0�z����A(�B*���ypd��Ƈp��Q����u-x0� 7���!�ϣ��_��,��a[�����������3�O@|��mp;���0�Hq��BDBſ��ז�9�u����n�:��:��x8�Lc�^1QP��{^TΕF^au+�`��7����(N?�#�p��q��L󽢔�<���;�a(���:^HY��\�V�q����:w�Y��t�*�V��� ��9�@�z�~��^Z���S_�0my�i�Χ�ﮆ�괣�[������
眓����Үp��.y�����y�G�฀9���?���&q��	�������Aww7!(
����L6�E]�P��X-��zʹm�u� �p��ј�6��du�c�C��+"w��r��^��2O�Cމ�I�����-��>���5�V�5x(߹�R> �O��w\�3A �������4ׅ,A601<bu+PD���7p�x/?6�ǎ�u��vzzz J���� kkk���2&��t����� >{�����E�>P_��V�� ��~>F��/B��iB�L<]_�����M�9 t>���u�Q�mu����)� �O��9�p =�n|g��5w�d��炠'�ki��(�vX�����q�}tǏoə��!�2��7�#���[��]�Q(PSu\L��,�0�A'�B���8u����X��l����r�����Y�{i����ț
�A��k�}.�pd@�S��Q�5�Rǭx8���d = �����f�~SM��������;/��rH�*x��9<��'6֙��=w��F���"���k��������ȕK�W3��-vp�4h��]��Wx�� "��n��#y��G��A	��ս��|H�~�g��[g�2����~Bu�?Uoׅ�u��Z�U��h5���A6F���?^�,~|Du�O������Џ�8Ԓ�^���"ƓA�E�D(d�󠻻���xP�TP�T����n�k �ɠR�p)e��v���V"S���Ɂ����5�9y�խp��;���r-�K��5o���eu?�ED�[�`�7}w�疝7>T�#{vu>���u�Q�muZ]��pιË?"Q~�0'�pد�ɀ/�I(x+�ؑ��������WMq���8r ǎsD86vs�1�Χ��S.�C�\A�f�̬jI���N��QQz��%S�0���OX�
��{~��v'W�v������	������+�}���=l��e�Χ�;�N;j��N'��s+���6�F^���[���g�B3���JX|�@{G�(E6֙��` ���8q�8��֙�D,� ���PUk ��t:�Z]��բ��L�����B/�AC�k�L���}������;�7y�T@���+����t;b����:	�}2��_����Kl��o뀾S|��k��N;j����<t��A�9��u������P:�n�파�n������732��a��m� o���A^q(����ı���:��x<����R������nQ*���P��xzʚ��Q36�M%��H�x��'fB����BZ��lT��ޟ��'>H}�/Bl�� !D��?z��������xP{fag^��וۡ��^K��tR��R>@�x8�\j㷻�^H�@M��g?�cUw�����/�����!􌶭n���T�`�W�X�C����C+���cuu�\�X�,[�`~~պ��5ْ5�f�^��q*�a�%g,� �k_��{r�n���Z��w�!�w�M��_z��6��%����2H<�/��9����Nr�ڌ�z+���)�����^K;�����u��)���=c`�����g0VZ��:�Fx|E�z�+�*�g33�2�H8��0"�H �H�jZ��(��bX^^�������n���j��3���5�֞���֏�E�@���/��?B�!���f�6�������g���o��z�7c5��!����u������ń\Hly�qD@����p[;�z�S�?iA;�!�@�O�o��8�lu�kd�N�==�����e��k�OjW�|-w*T����B�z|�'����rޟ�^�%��ZnϽ
�h��Τ��^�}A$��p����� ���P,Q�T���rVh�H���x<S^X�Q��7�3�S�<��57>�Ʈ��Ԡ]���	x��`u7\Q/�^�P�>����x=�	��9�X[��(��xC��F�)t5��ѳ ���b���u���:nz-���1��b�ڱ�6�`�7>]�h{�q��>鏼�GȖ�i��?}��W~��K���Z�ƴﵺ�!���bx�����!��m�S�>�>��2����100�@�=����x�H$�J��J�0>>�YNR*�P.������B����ԕ��"o�m��{�P�� >ئ����E�y�u|Z{�"�������]�֟h���(+���j�k��=DR�_yྨr����_˘-߈mЛ�	���鵴��	�~��<�s֣�	]�������p��������Z��cMO��H��o��c��ѷD��D��4��H�J��1�/�D$阠��ߏ��5T*d2D�֜-��L�D*�� H^��+K8�V�Բ�ՂѶ^�Zv�ǙV	�d'#��0sW`�}ʑ�B[�g1"��{[�{��`}��O��g~W�u?jV� �)ք���^I��P_���=]ޱW�^�fm\{lyre@wS(s�kiW7�n{��?]���}p����B����z�J��>��i�_�w�j�S �f��y�iB��e�����a)y��}U��{��-wE�#���Q?Ļ�HđL&�3�^	����ŋX^^F0��㱺���N���:� ���@A2��zwfU|�\��Z��|`���.�F�l}3{aj��	���?�H|�ƾ�2"����zc�{����{�3��!cm�N}=SD����U�0�[��{p�ʾ���y+����C�<pwX�A��l����B����C��0��<�sva�V��m���P�9�~s@_��qu���������q���2�� fc՗>��0��t�˨� D��ȸG�?�#��r�f�w��DL$��G{088�ѡ4"�aii	8p���-u�R��\.Q_�� �Lbmmë%G4̬��@ts��s��VX�4�����[f�2��G�~=��}V�����3�g$ f5ׯg��B_��Ŵ*�&�2S' �B	���� �"� �+F�{�+��CB�(��`��������M��Mu��Z�U���]���9�a�跺~S� ������}}�}Fn�h�י���L� � �PQ�"��=�%�^�{{���O=
��=ƓA�Ǻ100�`�y7VN6<<�l6�j��L&�H$buK�g@)E?���^����>���X�ױ��Co�Lwf��r�9�Q́�F`��`��0f�� p���H�oᜍ*ݐ���{o��e�`�"H@�3�[�>�_/�Ȁ�CYg�q�kigW�ᜳ#ʄV�%��wb��m��p"Nq4.`4�p,���>D�юYg�� `tt���XZZ���u�&yVb�!�J�0�?�/�D��e0+�老�g[�a�Q�[lpMe?jK�A��jY��jk���)�}���΍�Ҷ`n���p[X�A֞u��Z\��sΦ(H�FН�`���d�`(�ÁD�D}}}��|�zzz�L&������y���C�$��r���
x<�������D �/b5W��b��D1��-��^��uH��?Hh;f@_|,{��~��s�]�&o�����2{�q�kiWʛ��s��LPb�)s���"���b�׳q�y$���A(�buk�744�j����u���blll����M>�G&���A�V?��@ �h/�%�������(�+�^ 36��P��e���^{���5��߄���{?���+8�m�=/ڶ�4n
en�����:���?~����mpܦH�֠�]���>���xc!���#[ݚcB0>>�s�ΡR�`qqV���r�����a���l����d�9��ʸ��a9����Feu��O7�s߁t��M��L-���8�A�/��v�u@o7�27��v�q�k�$����0��Qw��Jp4Jp,.`$�h"�d"�D"�י�(�8x� Ο?s��D�=gӻ��i�����X���FdYF2���l�r*�~�
�I�s�^��o1*O��h�k�>g��S0�/B9�N�����P'�O��Nk ̖��ne<�ڳ�q=����}p�v�{̚��t�JRG�'CH�"����k�����cbbW�\A&�!�8_�W�z���`����ccc�z�ƱkkZ-c4���rs�]3*+[>.x�Q��:���kJ��0S�g�	9q7|�~n���^���e������:��)�����^K;�t"�9Ga�+G�c~��~��&�A$"!�Ǜ����fH_]]!�X���F87M�`����B���1�/a5W���u�}��s0�x{@���^1� }�_@%/�~�Og�:��z;�)��鵴���^K���sBu�TE�ܑ�81���`4����u�|:{����`llW�^���
!�F�V���zSSS7G�<A��T�p8�D�C�2�h83��3����W� �s߁0��}��MK��'����L�Bxw�8��{sE@w[(�A֞ux(o�9G2�@\0�.R�H��x�b8��H��D�drρ�ۙh4
�������MӐL&�"ۨT*�����:���UB�����屲V��|eoǮ�����-�zL
�(��@�,�@�����������u8{����P�:nz-�s����s��(��נ3�(N%	�#
&�Aģ=��㱺��qcj������Q��144�?�D6�E*�� ��8t�PS��S�D#kܙ����=�ƌ�=�4��?��Nw؊Z�>�5���/�z��gW��ne���j���C00�߭�s*f2��e�<�ш��d�h7_gn�X,�׋��IT*LMMaxx�,[ݚm0ư��|��h4����������E:S�dZC:��c���
���s�zP� �폁�c��姡��b����Ι��#7��n���x��g7���<|��y��}p�tE�'(G�����ׇh4ʧU[,�رc�|��͐>00�?4��:fggQ�� �2���[��$IH$�8�-�T^�J�c�3ݙ^�Q]��k��k_�p�M��vf)c�_ ���އ �����	-�q��S�w��2{�q�kiW�7���*=�𳅌��pܾ8(�RL�Rܑ���0v�:sQ���AGQǏ���$��<fff
�����ԑb'���H�R  �ǃ�"��^"��~�Z	�	��<�A/-b��E�Q]����?��0f��4�N�����ߟ���ث��B����쥎Ni���ZԎ-0*['`W�N�/�c{�y����	�?��'`�ǃ�� �0�����z�n�k@E>|�t���(
�T*��ﷺ���4���(��P���-���صl��L���U5m�k�Q]��U����F�ʗ!��&v�`,=s�4�o���9nK ��u���]C�]k���^��h���W?��v8�kb��ܕ$8�0��?��� B��խq۠���㈻+W��R�`zz===��b����C6����2Lӄ�����b�Xۖa��a$���q|Hó�6ߕ�u��F��s�_���`�,-^��~��>̧�sܶ6�ُm{��׻t]���q��b7�ݒ$iO7���w�q\;��:Y N�)�����I�ЗL�5�p����p��I���#�J!��"��!�����u�>��"VVVP�V!z{{166f�fy���X[�ai��kK��F���b
�M#T�^�@y��bz��7� ߉�Uz��=9�# ��A�]��ZmGZ���B��^�F�9�s[����O�	#
Ɠ!�%b���s�����8�;c~~�l333���E"�@"�p��l�r��˨T*��BQ!m�9�Q}�8F�˸s]�#n�G5ʫ�Nm�!�����;����zz�)(c?1vb�ߏ�:�-㹍���)���b�:�9���y���>��^����c�|>�խqM�(
�� ��
�:4�@�6���eD"$	��V*�����r�J)<�����m�R2����ҙ2�,iXX��j�V�^Y����
Њ� �1e�6����@�@������̽�������xn
enz- ���q�]X?���Cp*I0�0��B_$�����a�[㚄1�L&���E,,�1�X��b�a�Đ��_E�RCzi	��n$�ItuuY����@6�E6�E�^�̓�$��-���(���rܑ�c)W�n00S�^��vGfQ����!����k���s��iP�u3
8�%,�n7b�w=r[(s�����ِezI ��)��������>��m�;Y�T���<�Vr�����rgfT�7Fr���q�_��!Ѡ�JU��Z~��P(�h4j�Y�1�J%�r9
 �y�^�b1$�IH�dq��E�Q$��NqpE�Ņ:������I�Di��o��n��%���3�:�}/�k�ǽ���1����Z�h9�q���	�HPG�'��G#�m��vOUU,,,`i9��T��e��U1����υ8?�����d7��c{5�*ud�E��K�z=���F(B0l�zuM�P(P.�Q*�`�&(���݈�b�ö�@����A�
%�fk�:���Z��9T��~�{�kpW�X5}��q��u�&���q��)��P���)��9E{�E�OpW�H��y�����B�a`yy��i�-0�.�҂�K)���սe:g�����&L$Ă���\�ILCEx<2�~?�~?�� �^�C����j7���eh�B(�������<&����^��Aģ��pbP���[}5��R�џ�yS����� ��{ ��m��[l�{�c�vE���t��5nev��v'n��V�+���C�����m̗�n��=k˅�/ܙ ���8���@4���~�����������H��q-���tggT�뻻n�4���t<?�C�񄈉��H���!�%R�Q�
Q�E�(B���,|>A !�1�]�a�&ø�u]!�E<B���?^��G����px��s����N�Q��/��v����t���8�lЧ�����68��8gh�=�H�#Q�cq���<օd���    IDAT"�d2��c���T*�י���B��U��V�R0��64���q)��^�K!����
Y$��)� %�����(X�t@�F�z��z����P�@ �@�e���0PJ۶����"�H`l(�{��'�o�*�QI=a�Ay���6��B��Og縖# L[~�eۀ�q�q�Ҫ�K���L�D�8�"�����qS���i��T*���L-0�T¹9S�Z5٫Xe�������?�DХ��	B>����#�Mz
�n�&I$I�9�.IdY��(�i���aee�l�J�a��GB0D4E0li�d��F��1ֿ��T��c�J�r�0�1��[#S�>�o`�����}-훳[fD�# ���q�qܮ�(癏�ʘ�"�Xgn�c���a�aee��E̥�Y��RJ�����eX5���1� ���w��P|��ELLLX�4pmm3��X\-bq��BYEUe ���v+�gЗ�bhh�eG�	���ޝ�y�w����{���֧O���e�`0�	c� �PS�837�ν��*[�nl�Kf��ԽUw !��-{T�6) D���!	 �lK�,k�������g{���ђ1X�Zr�>o���*I��9��Z�s����<�����Q쩪ȗXɩ��dXF-�?xŏa�����]���{��a�Vc����	���]ŵ0�m����� ^���oP��d�A���"�o��)��R�`uu�|SU\ʮ�M���~��gV��Nh� �� ����L&���p�r�-�]�QTMXWr��-cj�������t:ؽ{w�Bz,��PS�e�Q����d��?��?�˽-�v��o@vֶ�;�=����t""��ꓳ,{��H*��azh����ϙo#�VkmlZ���9�g;HW^�9�^�M��R�UDV�!˛��T�VqiqO�+��相�{���f������Fۄ �r��cǎ��ܺ:v�R�!W��RNG��7���@q��	��	��x��.�������C�=��0���hxݰ���gm�y<����-��~�0��id�y,fjXʨxv�����`;��7�3��h��X&����M��i�X^^�s���م�5���i�<ׁ�]�@��h4�H$ғ�� �C	온���3(�|?$��KgU����p��3����͞�HD/&��w�a@'""���}����F�9�k8������"ot��'B
��i��j��Z��t���h�[ �_!��b�p��,����5*�V�ȕT,�[8�����m��Rñ:����t`m�Z�\ƾ���9� [��1ѩ�X�&dw��f����.dt""�m�ƾϻ��!�2v1�add�D��̷�z��66�PÅT��6�Z�Ұ�v�W������ �#]Ŏ;6庵Z�r�r�u���ב/7Q��0M�gGE\.FFF���ƛE|��.�uu;�ix��K(����"�����Yt""��������1	w&Lz�Ιbttt�f8S���i�".�jX�5�̒���;�`��,���1+bpppS�
�Z-��.J���0L��Yh�t�Z-�Ua�X����]�4N?���w��Ə �-�E��,{�0Љ��6�P@��G$LD��=�H"���q�|�~�F�4Md�Yd�9dJ.�Tqr����]����9��u��J�H�p
������˲`��Ml<�MӲ`Y����صJ�1�7�]�HDz[�m"t""���	%�Zk �+�����CE$�v�m�T*auu�r���lX��Q�,�V���m��V��N40:XE<����K�����vJh�o���"o�$�H$��d;�ގ;�~���K�M�^��nЉ��6�5��9	nKȘN0�`dxCCC���4�R)J5�4�RU'��ڗ�xr ��\�Vh׾��\֑�T��Dz6k |>B>!�������2�^צ4��$i�a\��\��E����e��F��;ѭD`:"��a�q/v&CH&b��u��ȴ%麎T*�|��tQC���jUA��zI#���~��W�hw^yD�V�Tб�kcd��h4����]k`` ɘ;�*�e�+��o�C�ၞ�@x1�ߏ�d��6^_i�{�my̕�'��;�v%I���� ��O��FdL�\�3B2���xO�S��B ��"��b1]A6u%=�\'K���{>���X�ב/76��^�����#5$"9$���RG"$��RqǄ��;�}N�/��	7�FB�I]/gdd�R;K-��[H�l�����3���{?p��Gd��e��-_��DDD������L��3���� ��E,�9�m�R� �Ja���B���yO]��>����:��dY�xr ��˙*�7���F���$c5D#+صkWϮ511��Ak�0-��+]�܉���������t��C��i�ŜN'F���]k!W�#�,^�V��I�;	��߅�
Q_�Q�����DDD����ǝ���'�ܥ�Ў�AL'Nbxx��̷�f��T*�l���*~�d��j��G�/a|�[�~=��03��	��u+ڦ|�rj������x	�D�P�'�	عcB nW	Ñ&Υu���EB�/czȁ�I7�OE1=���dBF2�D�T�T��=C:�fm�l�V��)� F�]Ư��`�]FoIlGDD��<��#oB��p8�����;9����<O�K{E�i��lX���z���2����*2�<.g4,�Z8�*�|A��Q�@y�Ch>�%L�S�|$�+o�V��a�|X�T����VW��+cע����߳��x<���o��U��PӺ��$!�u"�adЏ�������k[�$���bW��\��Œ��ޗRȶ���^�����=��#�B�9����w�����x�V7��J�\��Fkm.��)��q"cxx^��ߥڂ�|�t��.e8��II�/�d���g�������^(��u��pێ��&2�:t���{�|F�Ρ&F+���==�
�p��mH&K�T*h6�0͵�^��P����ҵ�z"���0���8Pl���lGd\A'""�����C �WEQ�
���d2)%	[�@뺎˗/c5W�b^EQ���M����
�0]*cld����vP���Ι�k����b��/�eT�9.K$��eu��O`t������RI�0�#�"���X�^�	��Lxf��D���H�X��]�eY�����ׅ����:vmo���@��h�=�4Љ����ĉJ>��mI��U �����t���l�覛��:Ξ=��WJx>��ɬ��*`�hv���޸��*-���C�uLMM���>�t:XYYA6_��tK��Z��R��U��8������s�2B�o��w p(2&����-�(m���*�X�u��]KcbbbӮm�p��pOģ��p`���-q��d��m=ǎ�Ӳ����������������]ں\�xgWJ��R?�l�m�4�5����iՀnU���~���۝a�f�Hg�X�j��m�Tx>/�{��59<��ϭ~��cp߻�
O��n����0�bd�uT�֖�O]�`8Z�P4�x<�e^'�6<<��b��M<�
t�f���C� ��8:�5,,,�!������������]ں�E�<�n�{�Lt�3�+�
�x�@�UEȷ�h4��;�!����i��T\�jx>k�锄���+����v���;��NH��5����b�k�X�P(7`�x^W�i���6��UD�)�ٳ��%ق��E4�P���h��\E�+l��{$[&tt""�9~��O��{eY~ 8���w%�I9�L�z��E,�x&k]7�_�XX*똪h-���ڎ�VVV�)�p~U�傁�/K(i�	N�'����pf��)~÷�\���v)M���P�6�+��m&�슎�x#�e$�-uS����8�c%�wp.��j�K ��z۽!��Brڷ��v&�H�J���ka@'""Z#��ϿC��?��|w����X�366�����n�a���,Wol��bY�Z��n����v���K��V��o�锌Œ��Xʒ�߉�v���
�c��zOd��WC� ba�-Ѳ�ܮ�.p:��P��Hh���%��a��3w8�R_$A<�E"TG�-�����ĎC����~�Mtj@hW�˸%���U��w�NDD�����}B���x�_#����.��m4��m�FZK-�F[G��ζ�[�i���rH�3X�iX�5q:-p:#ð67(ɞ�}��\�4����y;�o��X��;�"cj$��.�s)�BF�ΡF5ĳY���F�E4tu�����b�F�=�$! � ��B�'��V�:�ٶ]��rp�ܼf��K���j0�o���ka@'"�[�C=�D"p8���������"����WͲ�a��yeӒ`Zb+t%����le%�t��i�sk��������F���? ��_1��������s�>�n�v��Zø�@�p�x��;Q��6.]��L6�T�D�������-#tal���DSSS�z���F �!j�B�+���h[{�m��ݬ\���Ow���gN����B�J�k�t""�%=z��X,6����
�'�IW2��6MќN'�ޛ�D'�vʶ!w=�f��9�*ί�X*�xrYB^�W�.y�](Z�O	��cx�����_WP�m�\�U�r����mt��ix��Y<�\����3Y	+	�+� ]��D���m�t��t�g�n����%`��D̿�o~m�*M��߾_�7���������~Wr˱y�N}e�j�?��Z^����KDDt���ߧ(ʿ�F�o�BC�\1��ǃ�ǉ�߁���Fw��M$���-;"K�u���"�+�RF�b���i	�2l�d���z٧��!�����Fx�^�����B�c�3�/���F�u�
�I�}%�����8u����<qIzɑ��)�BX,���f�aA�/���o�M*���ǁ�G�C�~�b+���
�&͢��}�P������IϜ2[���d�j�B��]��a@'"�[Ɖ'�l6{��r�?�=<<��]�� I"������ɥ��'w*v��HF�D�߼��/�3����˫e�^n�Ԓ��~��%��=IR\��o c�<��=?���7�7|'$�W�C��˰�� ,����_mg�H�]�`�޽��z[]]��tg�5���x��?~)Ò�Ë<�"���4&&6�|�$I�x<�{��&�چ~�m�����P��۵т�?	�r����хY<�类IhHn��J�.�U]Fe��]z�&��oY�ڇ��~��JЉ��p%������p8�橩)%������d>o��X]���_���t�8����磻#o���`p3���J���Hg2�ŋ�:�/\h���ǻ�rM��xўv!�z��- +��^W�����Y���k R+�_0���?���r��j#�͡R��Ϙ�]`=�����sN�:�'��<H$جםa(
�x�)�O|�S�7��/�Sy�����y����_Ew�\pv2�t�k]uq�ʝ#	��q^���XOoId���J�뚺��\��z� /z�tݯ%aI��_y�
 +��y}�x\�,ː AR! ����=4,! I������]Z����OK������� $ɲ����LS�I����v3�U�$ջ�O7�]ǫ#�������Bl�;�DD��8qB�d2����D"o޵k�l���X,�^���n�4M8�Nx�^D�QD"�u�@�|>���� �S�����<~��>��C�X,�����D&�����΂V��T*�j����zJ�v�����'?��wm�K���e��L�Ro�Ð�����j0cu���������s�o]�?�h4�=���tb�����п;|��?l���&����bϹ!�P{�qi�b@'"�m/��~���7��y����f��]!��,���n��;�N���ք���p�\�X�T������7<<�n���Z��������~IQ�.���(��F��������ݹs���g��@:�F�P�j�vVU��B�/W*�o9r�~m�oq�r���h�ݚ���d2c���=�f�ՂaU!�ٛx��4+�fs��,ːe���w	oQW��m�՛n-�DD��;v�=N���޴k�.ۆ�K�.�X,k��Ϻ��?9�oK�t��iZ�0��j��ۭV�v����;w:�$I���$|>_$�N�f����n�����%I�$��nw���L���7�B�P( ��M�k��i!�7�n�<X�w}tmG��y�����۲��p<W���v��,�e nf�nò,�4͍.녝)��qD�R�DD�m=��; ��D�299��������l�\��,˟����ů=�`�����j4�������;��i]���g�r�<^���[���b�����!�"�z[{�^���
�F�^���u�	EQ>s���_�wmt}�>����V�5����ǎ=���(�e�)��7S�e9(˲�c��U�$q��:mKǏwZ��၁�����x�K�&UU���[�Z�G�,�����^��_XXp��Z\\|���������F��)��6R�*�JSӴS����$�󳳳?���Pd{�㿩���r�<988��e#B����p�F�kY�~EQ½�MbY �WV���~E�;t�A����^����q��f�r9h���i��J��ń��4�d�Ѩ����=d�&VWWq��#�ɜ)
�h6��L&gfffg8�z�ﾼeY_i4�S�z��0��v'�]�<���z����0�(ʝ�'
�6�.]�a�f��G=Q0�Ѷ��c�%dY��@൓����6Ս`�&j���iڲi��\��fgg;�$�}��^�T�gO�R��ӧOciii�X,�����������������w}t�����6���z�T,{v�ÁX,�����B���z�;G���� ��x\��{G�ۅa-EQz��іŀNDDێa
��G�Q�]ϝk[�-�R��<����	!N�^n6�=�{Kh48{�,.\�P)
߫V�m�Ggff����(�6p�ȑ�$I����L&#�w;�GGG�}>�ۢ����?�ӗ�9??�$���|�����{RS�ӁeY�����\���4�A'"�m���$�7}>�n;om�F�Y�Ցe����%I�Z���E��~�u�T
�R��i�iM�NZ��������V�mfnn�G��i��ؑ�d&���{rEQ�{�n�;w,{dY�^XX�[!���� x�ᇇ�N�ݒ$�/�1
ݶg�8�c��o�i���)GD�t""�Vt]��P(�#�:z=��Ւe �e]���Bx8��u}=��d2��r��iUU=mY�W����9rd{m�!�ѣG?�����|~$�H8{�z�z�ػw������j�:�n��h�Z�����Bv�\!��;���v�B����4\.WOj�4�a���{r"��Љ�h�8~���;�^��V�T��z�t:$I�q��	׍���$i����yf��T*�R)h����j�Z��=�����f�]���������o5��ɕ���w��ճky<�ݻ�j5R,�� p8�@ �x<������ �Mm�u�$I��=�mY�DD�mt�ݻ}>�d0��g>x�9�|>�����ro��<O�$i~~��n�{�ׁ���&R���j]UՓ�n�����x�ߵ���u�������L���@/���X8F8 ��� �iM$���j��je�On�E�h�a�8""�6,�z����D"�.e��|>�> ������Gy��n��~�h+}��a`ii	gΜ�f�٧���������H$>�p~kz��˦i�h4�z=v��)���TUE�ۭ��yavv6�i&�-�+�DD�-<��C�h4�:�۝��B�K�f�zW��_YG$�����("�HD�}n�  `IDAT�7����������G���ߣ(ʡP(t��ؘt���	!����d��i�TU=c��h��_���>�}�Ӻx�ޯ�Z�w�����|>144��z�X,��n/x�ߵ�}1�Ѷ��v�����s������)�J�^�k�n7��z�%˲��tF�nw2�H(###Xox���B���@RU5>??�eEQ��С�������B���v�{``������h4ڣ�r��j5����^�����I]�$��g����]������������]�l��XL�E�~�v��T*z��X�z����z�Ⱦ�׻���8�Ψ���c�_�|>����n��8�i�s B\�$�%IR²�;E���n�Q��&v�޽�n�.�{����˗����!M���Z�գG�fdYnt:�I��7���v���9{�yn�N����T*�F��8�j���$�s���?�wmd?���?^XXx��hL����.iC�r9���%!�?����]�:m�e�q8=��b����J��]��F��/>����_{��;vlW�V�5��B�;��߿�-�N��w�F�Z
�7��uK�Y�e*��v:��h4�D";��3�L�|^o6�ϫ�z�4�^��k��]ٗ$I�VU��B�0��][���zt:
CӴs ���z���Љ�h[�ey��pz1v���bee�,��?2Ms~ff��^�p�ر��h4>�p8�Tjzrrr]ב$	�H�HB��n�P�֡X;g^,��dD��XVU�Y�4����|�A��u>|xi~~���M�R���޽�$���Wmuu�f�aߞ�����z���Љ�h��˲�����L&M��������/ί:t�P����Z�6�v�G���\�熮)I�ʌsUU���/��z����T�鹹�������/i���j�:Q*�"�x����*�Z�R�Y�ן3M���������_�����رcI��,;7zl��jUh�vYQ��Z����U!��[��R��=���..]���g϶r���
��W;��Csss���n���l]�Z����ʊ��v�]�M3MKKK���B|���p��5��1�і�j�<�,;E��-��V�n�a���C����s�?�v��F�q�o!�i"�N�ԩS�����b��w�f��J�23;;�}��ìiۙ�������k4�7u6�FZ\\��������r�gωh]�ŝ���<�áH�$�b&x�Ӂa��>W��i�M]��ф(��H�Rh6��z�~�0��X��߸:HI��c���t�\�T*54>>��n���*��b�^��D���G���]m�DD��)��H=�&�(
dY�p�΄�f�ڋ�WUU=�n�nY�g����wm��>|�4??��r��$���o�тW
��i�R�<!I�'>��wMD�u0�і�(J�4Mò6~���rA�� ���b!Ę��ؽ�+�u�t�B��i�M�N�b�T��
R/��ΞYXX8V�T<�,��k����籲��,�ˏ[������������t""����x=��wL�B�]Lw��p�\>��9v����od�X���z<��`0�a�l!r�2���i�EUU�X��5EQ��СC��P=����̷��rYB�#��$�~��Bd�Y���6+��L�|tff�������m�����n]��{�)��,����Џ-Iv˲�=�к�w;vl�����v�E����ת�*N�>�˗/g��w���_*�rxvv�3��fff����c�J��������e[5�3M�.]���J�\.�0��������."ښ��NDDۂ"c���j�bN�sC?v"�@�X�l6�����J���W�T~�ر�eY�W8~]2�tlt=��j��J�P�VUUUO�Z��������y�k�[����WʥRiN�f���������k]�F�j���Z���??|����Zmiʟ�ɟ��""�W��'���t:������ز,���J�V+��z�]�z�ȏ��sw�}���ǝ8qB��w��6!Ŀ��o��b�SSS>�m���T*����n�\>]�T7M����?��?^�w}D �7�i�?��3�VkH�u�V��E�}>ߦ��LӼ��iW�՟�����������nj!D��Hv�"DDDt�����>>99y���TO�Q��q��EKӴs���B<-�XB�,����z�{�~��X,2==EQzR�FB�X,"�NM�k��i!�7].�<X�w}D��O|"��z:��w�GFF�{~m˲P(���D��X��j�!N�\�/<xp{�S$��b@'"�m��G�!��CCC�u�w�lEM�u�R)T*���LӬK�$ �].W��������l�r^�ױ���F�Q���t]��gff.��6��x�G�"��7�絁@�@0��gJ�r�4M�4��t]RQ��r���_�Ћ�-�����I�����O���߿����>����3����nX���������7Z�ݾz���i�)M�NJ�������ҹz";:~�����G����x<��~�N��=�D�
�n:����z��J��j�j����f�y���<cY�_=��?�k��6:m�����922��rl�0�r9�r9���Ӗe�����W���n��#z5N�8��f�o�$�w�m^�w��r�\�����~?�^/\.�N'�6n�$	�i�0���V��v�MӠi���z���f���i�Oʲ����s"�t""�6���_�r�>�L&���o����t�9��r��x�0�ow:����G?Z�wmDmaaaZq7��E�v�\Q��q8AY�}��x�NI� ˲ò,]�Bt�Pè�^�t: �x��r}����|�Q�1��v"-,,����j�޽����~��W�F�T
�z�R��Ou�ݟb�9;M�-�����Vk��(��� ��rpK��B4%IR�5 YY�� ,�ųG�i��~"��p:m'B�V���l6{׭Я6�+�JmM�Nk�vҲ�/���} ���-��4��]�EDd{�DD��t:�oJ���Z��WU�@0�wI�F�|>�t:m5����z�Y!��].ח<ȕ@"""��w""�v���|K&�oطo_����J�T
�F#[��O��=˲>��d�]�WЉ�h��u�4�������B!:88��z��l"�J�Z��TU=��v���gx����]���Ѷ4??����O�D���v��r��]҆2�L�|��i��F�qR����ů9r��w}DDDt�Љ�hۚ����P�CCC�w�޽-Ʈ]��i�4��n�����}L�w}DDDt�ŝ���-������{�Ngtuuuhll��%�*�Z��9�s�?�$�sssK������^=��Ѷv����E����;v����b�.�u:����\.k�f�t����$I�;|��O�]mt""�������t:��b��ر��D�]Һ�蜹�l6�WU����n��<���>"""�X�DDtKXXX�����h4zώ;\v�B�E��ih���h4�5����|��������7Љ�薱������G�h�-###�d2i��q��"�J�^��TU=��v��333g�]�:�R��/��w�n����[��xdbbG�{�v�]�R)��喦igTU}Z���������7k""�[:�r����V�#�P��@`zrr}�Ų,�r9��i��l��4�eY���|��V_�"""��`@'"�[ҧ>��q��5��x~#
�.�zGGG�v�7��B�J%�����l������a|��t~�����oJDDDd+�DDt�:qℒ��~��B��>�ow<w$	x<��\S�r��L&Mӊ�F�t����eY����{�'%""�-����ny�=�X�0�?t8���|�<�T8v�b1�B!(���j�P*�P*��n��F��N��eY]�T���k>"""��Љ���XXX�B�O���|�i��=�r��PH��|�e�?��v�V���^���n�:��J��Z4�eY_O&��x��������1����~8,���eY�[Q��n�;�t:��#�(ʀ��].Ey���a�4Mt:aF�4�Z��-u:�|��M��$I���4"""�t""�W�g�gq��u�$I{ �B�:����J��e� BK�5�k�fK�B,K�t^������nc'""�WNDDtN�8�,//G�^�"l�� ���4UEQTI�J�j��V"""�ZЉ������l����Ѧ`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�t"""""""`@'""""""�����SiM\�    IEND�B`�PK
     $s�[�^�}    /   images/c5725ab6-c6f4-4984-98e2-b9c0e10adf5a.png�PNG

   IHDR   d   &   2r>3   	pHYs  .�  .����'   tEXtSoftware www.inkscape.org��<  �IDATx��Z	pTe����{��,$�HB$��l�"5�Q����W<�T�:��W.㎖����MtP�9��"00hÚ��N�{�e��w���f)q8ɭ{�.�r��|�W��I�@~br������;v,v��	Q��z�(
Z[[1w��.�u��C^z�%���~�7�|3���+oڴIe�����-�m����6�- y�W0h� :t&��+��0gΜ.���s�!77UUU(--Eyy���_���ݻg�����������I�܅��]j�gȊ+�l�227�x�������^���`ɒ%�>}z��
��:u*֭[j���]�v=l����rT�6��YYY�)S��?���ZW�����_�[o��ŋc���d��%��%�8������/�9`֬Ygl��������Z�---{��Y���?��M A 8��x���Ș�p8~I�t��l��+c��"Ҕ��p�u�V���(Ĭ"���d��5�߶mۈ���ƙ3gb���O�!����M����ؼy+L����;�����bq1 �k���4Mk������r͡�m��ә�'��Ӹ�_b��c�B���7AW������[��a�A��#z�&��x�F,|���Ƀ�W�Lg`�����S��9b�(dݷ����Y���c��Z��J����"t,�� ~7�?Yx�~�ĉ�%�MI���t�V_��������hU�~�>1S~����1E�Mc~���'����Ң ����>J�̜��W���C��lz�i��e����A�5+zXV�����^�+J��10�j�¯,�B��
U�L�4�s���ty��B�$0�5�4�.�R��&�@ ���i�Y���c�$EU
�q�µ��#��_;��w���Ƀ�&	GN4��׵����f�"4ͤA�t$���F���(���d����ۘ;%���Ut<�d˖-hjj���g�Jn���?RD{���h��� %��)�rt�l�Ŝ�5qcĀ|�g^v��s~]���y�Nd���W������4V�����_�ٙ�1喑�<� N��66CE�1vx���i��`���곽x��8x�����.�c�gD��E�����D`8��k\A��;v,��D�&�>5���#�WB�䙲����Rs��0�����sD`�W;�OV��![ۈ�E|����
CKr���΅�a�����+J1al	��al�S�q48�#�_�u� ���S
0Nu�6��W��aP�T�u����l��¡,Vr��6SQJ #�
�G,�1��x5�E��h�P��;��ы�����V�7Y�6��/7��t��e�m����m��|����Z�	���HvM�H	��v�1�!R���*�fb�K�]�L�u�n���W���v�sC5̞4���Q���N�Z%�GRѾ�n���=6�<�/�=GW�P)��9N0��M:�v�
�s�R'��%�d�L7�l��7�9�p��=��M�J��`
����czȻ�YL�<�*�V��˓b(��8e����2x���2�eO-�o=�k��C^7Z�[HWQ������tE�p��.D4�����h&Oj���κX��1�E�~(���A������|�qꐙ��c�:�qb���A�E&#��;�2�� *�0�-����\�~pj��Ŷ��Q�_<M���haUу�AJ	P�VX4k�� k7�:R��׆���o0��C%'R��i��)Lf	�F�N'���D� [��wx��8� �b��&Q؊te ��#����>�_
)D@B�+�Y8OX��tטH�#��PS�[�gEBz�1T�oS�#�;�oy���Jog�LpVi�#����ݶ�^���j��I�kr佦x��j
�dq��Zt��*W���-�Uy� ����cʏ-��Yb'�������o���*�6Y]
��x״��{{?X\�p��{�rF�B��XcL�0����Ά��db����G�5W �Zr<v��b4 �t�t�!9l���8	䅆�f~��0���*Zw���y���|p���v��_�+;̈́�Lh�����桪�ح�>ڀW�n������:5�b���`�V�)t��Y}�1�EA�((�}{7/��d�:�zHg HBG ؞�;rB����l�D؄�����#'V@��z���t�4�D���C�ʬ��#�ɐq��
�U��̺Cd�����4�R�����D��<ͭX��J���5Օ\E`E_4/0�x!	�v����V�W�T�M;�-$G7Xz_�3���3�6i�!�&�����x��ң~ၼ��X��Z"�H�s�$N,Q�������=	�Iƌ	%���4^G�9J�H����-��W7y��YAX8��ƅ-���x�"�`#:H�O�4�OvN��A����.�Fb�u��pD~{�sb���8��5E4$�s��FX�m.2T��F��ch�L�z�f��h���L9B<c�T���DU�S��(&���/H1�9�D�mrZ�ת���-���Zn2�I5�!v�i�M�&$Ż:�9Bߴf���Sa���3���@A����
@��:)�8)��X���}q�a����-զ��[3������gì��1nPO
[2�'dYAgD����-��Dv"A�l
�����!�&3�L:��E{�ݪ���`�7^3"'��2�'�P�J�����rH�t��,6#T`��,<$Iy�cO�{�K,XwQ��X�;�k.��K�t����ܺ!d��=Æ�c���}���*;�F�ftv���+VƠN�K��J�r��~ u��At%�U�<F���B4�vr������{�Y��7�|��R��>t.[UCK��3H8�+f��)����e�v^Ţ�!�t�F����8��m`����\�_��f�)��=7,X���L��U��"i_���1@X~�[C�/èZti��U��=�;1�������パڝ
� �\�5��H9K��(�����~sMh�����a/^HZi���^����&;���a�W�	�"��T?�9�����=q��"/���OY#(�j��c�]�]ޏ�E��3-w�2����xu�N8��g�_�t�M��
C=O9*�b��~X�ɗ�y�I&=k�E��y&�$��a�$�IB{�BI��v}�\2�H��c�����aKG��Lu����u0^�u�uǺ*?>\�9<��?f^�W+ 5�Xxj7]��!��i��uUx��*4Sm��/�x���n����>ك�>��>4�.f�<s���"�/�t��AE�89�Ho�ݜ`�q@B���9�w$ǢN����.�ێ;����o���e��n�=knż�33��-=�zUG��Ry�.�C�H���Uؾ@+7�����:���N�<��3d�~�#���1��2Ӭ|��-J������Y�twL\qI8�[�=�N�G�<����I��Lk�Q-&Y555第���?S{��aﲯ)8h��f���Z��&�,�G����<q����9�����n���_��6��V��RD�n �f��6s/	#�{�|m�t@����.)�e�=��gO�0lt�E�r'�Ȫ[�y��"���� BWi衠��p z0@U�E��F���M|J"�[�h�%��
���������Rϒ����Vk:K�[3���?���,-xwt�EY�P�1�@����yd�w/^�����'���kpJ-(�e�:l��A�����ǽcYzz��?��_oKK�e�hxIƧ��3�g�6p��3.�������Qʣ>/+tG~[g+-0����2&�[�7�l���$--�h����ÇO�����nݺ=@����\�z��E/UUU=:hР�{�݁�E�l��&4�vNR>q��h�Di��nYKL3� �QN[j~~��L��}665/�E��-�	���]	�LD�16�13�Z���*�`+bk��Zȧ�:$s��Xax�u��?���J Ijj� ������YSI	T_||�ĉ���v3�GJjcx�Z��=;l<����?���.��ݻ�?y�����̧����6����0r��5�>�(=�?I�Bln��4�����*� �+ãG�n O�.%%�y���:�}��-]`ܸq477cڴi���[�r�J�u�]gm�}�<pʔ)ؾ}�zR�%�'OΩ��v�����|�I�QݤI����<o q�\�Q3���=z<C�1��H#�%�W�^4q�D?��YYY���p�M7u�}F؛ϲ�2\��a��VS\\́`��+�`r� RYY�Q�F��TE!���7��طo���!8b���[&L8�>f̘��<���7�0e���)�c�ҥ�8�faf���cgTTT�� � LfϞ��<�?9� �w����� ?1�M����    IEND�B`�PK
     $s�[y&��:  �:  /   images/4a8a1475-7a47-485c-913d-9939fe0b1f0f.png�PNG

   IHDR   �  �   �'L   	pHYs  \F  \F�CA  :�IDATx��|U՝�WNN�&���OED�V���k��tfnי>��/���V@�u��;m��:N��i}Њ�
Z䡼!� �$�<O�s����a�${���9{�������C�{��Z�������*������C��l����s�D���!y�2p\�@FFF7��űmصr��5��gpN�}zԨQ��w�\A�a�S�N�������,?~��H�l�]A�c�{|��In����q�9'N�� �S�Y����*+**BJ0�� ���cP0'�g
l
v&�����������0''����x�w�(��B�� CQ[[�Ĺ���#S}?tðk4��h#,ʻ���#G�<�[�0l�y����3f��	�B�����(/��*��p8|r��mX�ط+�_Dؽ{wvqq�<Ծ�P�X����~ "����<�X�f%����ߟ���;"X�����������lonn~eʔ)�J� "lآ!{İ�����]VPPpɱcǶ544�4k֬%�C�q�I��p�(D����@AZ�!C�\TSS�G�Wo+!�#FUUUn0�
�K3�Ԁ0 �p�>�J�b����1cj� G���Vb���E�4��snvv�Ў���H$�j*]�b��vX�M�����̀�_�N�z~^
Qx_1P�;sss�����w�}]gggm{{�	<G�a�Y�>
qL@�Ǎצ VG��Z�V�2�3X�cs�������B�r���$����Z��q�dYY�{j�1 ��i:
�-���|
j�3999E�9 7k$2e\�ʶ��#KBs��������z<;�\�'d�((K����3�cW������DlQukk�a�\Mv�îk�V�L�B���WJ��Ջ�"\���N�g�ư@ n�آ���Ʊ���w!*��B8�J%��x	�h~a@�� ����|�&�7�o�1��� )+...��577ğmM���.�88��H/��^1Q܊����X�3hS��9�!�Ք�����v�䬝�٥������Ŕ)S�vBbZ��~jjj�̩(p~ܖ26d�\ca���
#�~.noo? ��������͛���u{��D�a�󜤁�ud~~�l�,�rP��*��B}���B�`��`pXSS�[vz�P�TL�<���O��۴F��iq�� j�Y������cRnnn,G�� hL7��׿��2hР	(��X����Ǖ���Z5X=ךk���J3�R'O���gi�磀q�)
L~Ͽ��ACp-v
��pj7�.�T��(�i�µ����u;�oy�Λ�6G��ѣ_RiD�	�bDq����bDA�K�nPhI�={vK�gnq4a{�c82����	���y�p���yW;v����l�J�J\i��'8�'��Q�'�֝��q��u~cc�]^j���B�!��<�a�*�W1�8��d�K�_X	�Jݴ����e�SZ	����F���v�C�(f�=1��9(�����BozP���½��ó�Q6��M�\+X�#��+���ҡ1�6)����vϋ�⢞�l����a�՚5�������*D� 6W� .�L�.�9*����Ѿ�
?�W>'-�QUU�HMdM6
��DD��W���Fy�p8܈6��l\C̖�vcn;2B����D;�pii�Q�c�B�쥉�+`)�q���k�
ϼ���WX �G������m1qXn����A/�[,��k݈��?ϩ�0���0��y(���$��ipU�VF���"��Q��Ōzbg�}V~~��|>.���`�=��?_Q>�� �@\o�<�х2y/(y�jhhئlN�K&G�`�빿�)X����\R�}�� H��3g��)))��x�|-��*��9�;���l�-v�2,Ǭ��Ɲ��pp2
���L=��CQ����:�ſ��uc��k��zB��
�n3����@�� j�n���B X3+���z4d�K4r��7�H{�h�[����FVV�x�v�� 
�P7��-z��팞�fպ
��։0�#����c��#�6ō�A�7��ewm�@ ֹ���zܘ1c����0P ��}��Cc�"7�y��B�b��p��p��c�G�N�}� ��v�������}�F�wap�e`Jee�������'�NhW,���xƱ�1:��=��
�|��N�A�pvO*��+ap�'.��j������!,�H���hk)�&�FMMM��Y=�ݑhpO4x�k"
�ľKȵ�o(�+aD"[�ga-�s���k#c�cK?�(!!�)�Yb���[=�m`-ƛ�~{{�^��N		���cǎ-++��{�0�>=[nt���1ն`�䶶�CJpLff�l�^P�7����fg�]�&�����i�W���O�3^P��`o?f�����|xRF�-`)v'�UЃ�Q___<d�Ow`�B����P�-E0&17��u!�:�7�R~!
q̛���B�ta�x��v\%�����:�f�W"��o�X.��U��6�i�u#�?7�0��N�";;�v����c�8H��Æ��y��ĉ\?a��n������qZ	��v���0���37
�!N��G�=�.pwGb�ِ��a�@�/r�Ӂ��rPc!a,�k*�0`-,[ X�B�y9>T�ز���a9
�	a@�JpXv[�]��/�au��N��������:h���߿?ǫ���0b��l4��/JF	IaРA��Dv9~�8���h�@��lZSBR`�F���0`)r��y�0,}��E`�z'''Ǳ�wO�>���9��j=O}:,݁uN��W����@c�VA���/�R	I�\�GI+a(灚EIó�ϳ7F9�n�f%�7"C�����T!�"A� �"A� �"A� �"A� �"!J8ttt�;�9t4ȓ��L"���˶����'���'�u\vv��믿��U�#��@].|b˖-�koo�th�d ��]�W^y���N[�F����Λ7o�[����X��[o��4�`0غ`������t���.����߶m�"����~F������СC�Ϝ9ck� ijj�(++�7bĈSn��Ν;�����X�v��g��"NIII��_�؎;����˳+��f�������="Ѱ�\W�gϞ ���=U]]]��v�t�gϞ���Q�NX9~Ȑ!u�.gaA��ʀF[[[��ӧǇ�aGA,NŁ�M�<��75� ޻w��tM�6퉱c�VZ9nd��W_��@��`�*��#F+���>|����fee�M�+4������I�~;q��V����(nkmm��مte�	5a�D{{{��Qۖ�޽{�ܹs_v��/����'i�J<7}��V��(2 ��������%���ơ������Ӡ	�r���+QC�]TT��$4�����p,�ѣG??gΜmV��˶u��aAg)!ʀ1�0�m�����ͮ���ℿ�įH���\���#F��j��x۶m����]��sa�����(�Zuڽ�(%%%o/\��9�=lo���S�N]���0��}�{�e�=eU�v�Zp�ĉ���DiB~~��E�=-�b߾}�Ѹ_�-"�4 77���%Da)�����b��<K5"��ٮ�_~���M��SUU5��V6��+"���u�x$//�������cЮ�D!���|
ܦ�K/��煅��>ts���;w������/"����6o޼G8������%;v���H$���x�������L�#F��r<�r�����d} "����ӧ�����=+������k��(<��`/"��	�);eʔ_O�0ᐕ�9	q�֭��~�l#���ĉ;u��w�_S
�F+!!D>`�ر{ƍ����<	���ڃ�`{VVV����x�W>7j�F��qJKK�Bu�E�@,-�@����۷/���(�"3lذꊊ����fF"�"n{��t�̙�W�	��ã���Ԡ�}������%A��A����M����񕕕e555�`��(((h�>}�;�����?>���z��"��yyyM3f�؍F��5�Î=*max����X�]V�T�=Qr����J�T���dee��R�8:����Pt�������=D)��bgnn��oN466�ݻw6D���aX >�i�v��6�D��A�,��#t�($�"��훕̨*^d@�!9��g�...v@�VW�9��� �`h�,���J����+�Й9��IP�d��� �߻�vgU���A���j�����9�H�HAAAU��O�2i)�NȴB~(�F	��{�B8G+??/\,#޽B�	���dX�\y�ٳg���x;��<�.�M+aPȨ!0��G%���555ͅ[�3�X=�����}�g��^W#m��Q�Fvj�{ρ8..,,�8,��
jkk���o~��[n9�<DZ�nk,�sE
a�*��X�����,uo�����6���222<ӊOad����fO�R�677_T\\���\�37nܸ?�T����@5�m��chXώ��RoU}}��~���-]����Z��������9�g����߆5�p|&�?~��Wg,Z�(��}�[a�B�Ҏ��?&$�566N@��R,,���S�N=��_V)Ɨ��w����d՚�E/�V�Ƹ�8��yꩧ~x�M7�^z"�N��hkk�4	e�8B�jZIIɟ�����v�7����a�B|W�ZZZ�$���8555M,,,�o�x��eh�_���V�"|%�&A�&�J���J�?���߱��!}??�R���Q�eW�|]*X�
X�=V��0�x饗.Z�d����z�7  :::$������Yϙ��VF����+��+�|#4��J����E�@>��j�r<����TL�KA����1�4 m���Sň���</޸q�m��K�d|!���v�J�&�8����=f�x���Dz8"����(������ya�Rdb����Y��.�ʱ8nȦM�f_w�u��/��>iq$��bi��� -�b'��	`JH;�e�b�d</�{+!�@a����������%_T�9�,�6bc]%O�J&����vp�/Xj;��".d������ȓ�i�
�Ua�l���U��0$hZ�a�ҫ���D�À̦��7�}ι�"(�g���`Z�����,���M�;�@~~~R��{Z�AM.))ad�>�s2�-77�=5���K�Hҥ��N���ia���e%�'�p���m^^^Rg�zZhca�/�H�r�fgg�0�����0aB��L�'�P(��qh����~�����s�����^plϪ0�5t�$�ia����삂�o�A{{;;V,�1rr��k�ya��'�H?���K;�*�x^%Ç��N�gϞ-�z,�!�ԅ@\�zD���u��cE��c�]�KJJ,�J�6---�i�?���_L=/r����a%������*�f��/��14A͑t�*��ԩS��W�BLI��B૫�+9rd�|*��#޹��ݩhx_�;vl��a��9
*$��L�:����*�A��~NV�A��7�`��hcX�7��x������srr,[ ��lhh�R9���;'�9sf1v�k���o��i����QPP�#++�lmmmq[[���ʬ �zNp�����aZ�!C�X�l��-8��g�xTr�=��P(tF%_	����BJ�'N���m���5j�9�Q�ϛ7/i���߄���ah��a� Adٱ#F���� �H�� �A�Ə�d4���m�*++G3����9�WZZz^;���U���\ϚE	��̙3щ��i��_VV�ua�#,Fҿ��Ka�Z�Sx�J�&������NY�����������8�O*��V�G���2F��~%x������kZ	���*�쒝��{�d|)
�A-Ù�\�o@W�����N����r
��0�&N�X���/�1f���f����S��z(�cǎ٪��5dȐަ~��R�����Ǡa�Ȕ���Uuuuԍ�
�cǎ�մ��GT
�0���ͮۖ���2�T���Pv-'	�M��q�<��:u��*x��5�.Rwkk�7ߵ����?8��}�G~~��#��󃢰Ӧ`��)S�������T��t�A����۷/���_��ﾫ�O���8Yb� K34662���s(�ɓ'w�LV���O*ExZ�5\�P�<qL�4����<�blsp�CF��C�|�ԩ�0�@1P���@�����"eA0</9mڴ�8hD(����s�B�M{�^Z�C\+s��1
��G��ݬ���Q��-ܯR�oJ6b]��YKUUUE�1a�m�Dq�Gʭ��
�V�cF��c6�)
+���G��Z�T)�7� t��>uUVVF�ġIonn�pz��Z���@�����%H-((P�}�b�������V)�W� Gyyyt��wމvBk�ΝQ����B�x<��d�"�����e%d�-g�ȑщ�V-5D�]X��.f�	#Nii)�s՟����N��6�!QSφ�n�af#��P�6뾢4�A�!x����N��ʇ��X*�m��?R��� t����h#�[
eǎ�5��-c��9ܐN{I]l�ar��F����MȤ2_h��Xd����G�0�Ӡ �z�s����z�/��g``���S w����(�@����ﳘ�h(�z�={�bKR�Nh��Y�|�T���!�\s�:x�`�z��5}cZf�u{s�HW{s&�%��jj�a'�;���l<�H�,� �둀@�9��K����6nܸ�B��>�(U"m�A��N�6-�0���ߏ�C��_��^q�����������8N� %u1�[�9��8s$�������/��b�w��h���s�ϡC-G�<��֙3g~Yy��F�^�/��	سg�9��c����)Zfh52n6� �eA������_�-�8|N��x�����+��c���t�<�y��W7ۉu�,<-��gQ��@ϴ{.kB|f��)$��-���D�$PZZu�K���8I��`zt3⛩O/;��M���ʍ��[G��%Q�K�'�3��^�>��k_n�����{�s�_�\��ia�`�n߾�d��Ƞɉ��B��(9݂� 2j�.n��2(dz�ʚ�')Rp�(�3m��݀�57��Mdt?`�b��f�1\�nr��?�g�Z�e����׾&O�̝;���z�?��MH4v!R$t�ب�9h���ԍ-��� hI�:e�)dԅ�x�"�@�-��	�w���Y�t)
d0�c��w&#�N��-���-�z��ӧ�(
�߅�:���sb!��,ōȋ}��x^��7�xc	j��!��9I��������#����]����jHn,�@(\5Hdu _�F���,�e�[|�o��<cӃ)R����!�������WUf����d<�{x��g�e{�� ���?�{��k��oFF-r�^l�xƂ299�wމ���e���vkR��3b7ܭ Gr����	�&�qM<*�0Eћk��L���2�����!��7� �f��ذa�wP���mF"�g�|�C�Ne���g�F����i�]`-��q=7/,��Lcv�R��<��������;�����g��M�
_	���v������u,\��-�L6*�!��0[O��x����Sp����B���U��nh
�s�2�)�x�|�gu���m�˗/��(��g߾}�Y�K�,�Ɩ2�@77�IX)����Y/�b��Ժ���4��QF�!/��?Z��xZ-���-��%2�¤���֝�i�(��9����50�����SOE���nf �+�{Xp)��s�P8��۠_��熚��w!�Z����I���J|/�y��<����AX3=���\G�.�䒤����i�zZ�x�P�:��߼O���V��B��񹹥r};������v}/�8�8z��Z�hQt�"�����1)Bר紒x9>`�=70�ޡ���E�br����DO�F�5�/��(�p�BW�N�p����/L5�ZBVJld�i%�8̤_���j���j�̙J�K��b�eN�׍����F�]�vE{F���b%S:{�(�t�0��� 4����Ztu�����$J�}��9}�tt!�@�XO�#k��[�F�'�Ś<yrg~~�7[�"�&�ȑ#�����#�8� ۷o�y��n{�c9j�IJ8g��]hT>z���0���FO������>\�|���hH��k��4e���}�:���d��p�OfΜ�}͚5�-����l�}��i���o߾� ��²\�k������&�6>u� L����`0�	�G�O���r��~F��B�B��O�:�5�ѯ����g ��`I�Ԝ��me��1�����I�����y��qx�3�]s���^r«�z������]��%Q=������- �	y�A���q�^e��sssW�:���u��� ����g�N`��t���1��z~$���B����*YX�H��9�X�8��S48�Q{���ꪫ,��B��b��U>�W�X�r%c"]e(�j;��.�k�c�r�7�B�B���cp�SA���vO�JŃ*�g����p�٬A�`%�){�zG�����O<�y�m��f��W�@a�v�E�� {m?VY���a�t�p�p�ҥ��~$�R¿���Ҝk��毃�:��������w+P�V(�Xz�8⻆&c��������O�0������w���<��
�j.����b[��Y��T�m�}f�����J�a�x���J��رcw�<�"F�<��i���P8g�9�]��gӔ?�nݺ{�-[��XR=�0���+;���_���Z���r��t��9(�G�&���w���[���?����ν���9p;��_U>��@M3/�Lr���Q�g+3�jf�=A��.jng�ت<������ӞU�A�NAh?�뮻�+��yap�/�Q�%��y��9F��,G���e��!�3h5��BÀu���{���:e���j �a�:���d�ya�]��+x�W�J��ǯ}�kv�~9�F�{���2 4��;�c��CȧP1=���+�|���χ���0V�^=y����=���P�T���&�py���7"�XzP�m[�|��ʣxVp�{���T�te������}�05E��������
b*,�0���?��wVYYy��{��yl�ʕ�v$�
����M3��F_���>ޯ;8w�����(�v�����9|g��l�W�QPP��؛�T1�'����z�5��qd��O�r!PC����{�=��@�g��{A�)� ---������=��>�y�.��j�1<'d�m�}ׅ�W§Md��&.�B��@2L�/���'�gV㻉T.}�
��{lŊ�)�)a�Z��J�~��h�4��]���?M�~�bWa�^s�FL\���t&�[�n²e�l����7X��������Ga9\Y(���ڵkg������6a?��%���=7خY{#33�N�@;��D>^�KZt���9���/ᕾ�a������U��.mcxBx�S �M���i�5QB��vQ֝={�-������@��O+;�8H��aK����Se�ь��nB�.�A�bR.�d��~6�!v����\�ȉ+W���}}�P��GԶ��l2��8��I�i�ٮ}�ᇳn��v�Q����\ךl��W�
�����/���;���Ra����7ㅌ7�v��_y��}��w&�󋊊�@������f����ap�,�إ����s��޳�о���a���5��9�UJ�Lܔ	��@�݌�]��C0��$z22�d�����}m2U��Ѷ0\�g!���הy&�rlF��{�II��c��գ 
֢S�H�g[ss�]Ӹ�P<`�-���+Q �gB�=�	��f쾝��MMMw^��W*�LE���W��3�P�IE���<ݥK��)����I"3&A�Fݍ�Q��X�"�Y* ���{��
�y*9Nu��3��9�H�0���(�A��W%v������n	�K&�e�nC��X��$,�'��xgnD�N�8�&�EA�����:.�1�a~�\&++�����N��#a�Ŧ�Q�tq$Ex�1|0e����cxik�I���~0�n�!��*{p�a��Fĭ���������~��_�s��=�y-�ś��'��p]I��E?gbUXgg�;]B����hB���.]���D��W�\�����ь#��!i�pU6l����E7E���qX�v��b[忔K �p�֚H+��p$��U�V},33�%e.b�DŁ�\�fW�k (�_�ڦ ��>�� ޅ�&�到2�nd��h��;�@�B���v�����	��F�����ȇV��10\�j���0b�b�ˢhB�y#
H��!
��3�����^�؄0�
��ވ�caE%�g�?��)V.���mBY�&�5��b\l�BpSx�m�M�(vN�S	!��l_ġ��a"��;e��C`��ի��<���Ԛ�����s5��M&lT����r��D-���íx�F�At������/��y�o.[�L�	�Uo�f�M�Ӵ��7������(�[��}�����q��4l������5&X�����MrM������鴏9������$��7��X�f��H���/���b!�+A��<��  ��a�֯_5*�e #�`���4_�D����/�Wn�Q��c�u�}q��L#�N_E�<{
�4�����ps����p��	jw!��K�KA�X4�����2^�*�p���KM���/�$��Դ�T��؈�=�PX����;F"4=U=�]���e��;��Q��#a�/���El5�k �{!�v+�Xl\Sc-O;�;p� �����0�����}���?�8������_���5���q+q4x��V�.��^��16�V2ݨ�iB�;Ş�U�%(�իWS�%psaa!��&�=����ߏ�r;X�7�"p��F��Ng0|Z%�ֿ�u9���gb�k� +V��1�ǋM^�����ܟ��		���x��R.�B�-���S.�\`(�L���!���e&��e��;xZ�
�h9`�LF7<���(�U(G�f�\���Q\�vt	;���0���@$�ΠIOƠ��X�	a:::8	��e`96��f�]q���x/��8Υ�vε%4������oU| <����VI�s�!7�_V}J���B���!��3�ua�5��&��v�e����;��;3%,pX�!��O���Y�V�E}G%��k��ӕ�N��$Ԍo�c��d�+ �W��9���B�BT��5�[��nI+W��Fz/�H��^X��JzoĺiO� uʬE�;e��T�~���h/�jk��>ˑ�[���'�xb��i/��QXXȖ��%p�B&�cm�p8|���Xӕ1>M�.p����4�6CZ�~�4a�U���
��+�񶪪�o�g�=U�
*�ꮯ+�X�r�J�&!�Z��T)>�v���e:�@r|7?TI�cV(syț�.]��H�u�>���(�>�G�y	���[
����4�gM��tJlR������J4��S�΄����o��<��/x���}}��Wa�]��K�;lH�(HAA�"�����p��3!����F~��%�P6�q�G�x�����r�?.L�mt��@��#���R/���˗/s��	�쳛��ڕG`�Wf��n[�3R"�2r�1�r�鴙�H�����������������d$��P��0Qv�ƮT�W���lp�v����3��D�E�Raa!�����Z�~��B�j�3�FW���b����O:��h��j�KL��gzNy��:
Υ|W&W�مm7��o���r��̓�]���/����P\�h��߸�(>��)ٽq��љ���_ \Ӭ<F�L��
Q�p��n�B8�����D(bp�ay>��#N9O���Q��tfF�S��2�p6msssBa����+p?�̶U￫�
�|�+_i�������A>�A��Գg�<a�\}��	ߴ'H�/����8��%�x�^��;���Zp�2PĖ+��r�2l�A7��s�����ن9���s ���)�@�3���3��9k���6aM�+#@o�kN�G!6*�o��>�:'X�pOUfy"���n�0�Ќڭʣ������4�������h���3��u��-�>:���+�Ue�CYYY_T��8�0�uX��7�G�3��~`ǔ�����{x��]�V�x_w��}$����ᮮ��z��}f#�^b�ٳg�*�r�wY�vm~:MyI��)a0D\�O�j�v-���LT(,���P�,4�Ny��DC�v{a~To�W�}��@Z��K���qSm� ��F���0PX�}Z�3M���]�F�s�1���}v)�@��5I$�>
3�r��QՂ�0z衂��6S� X`���� Va&�<�����c�2q~v V��9~l"=��SA��JS1EQ��777�Ak"��U�� ?�UFޙ[�7�ߪ���7�@r�����J�b�A��A�
J��t��煁g5u�n|���˵v���k*zҹ��0�=�j�G��1�~m�X%C{�DR��0ENNΣ�~֣2�u�ǹ�Hh�2�&�{����L��?<��{4>��4�K�f�N4��IA����F���|����uj�mB�PKV���#+��1!�(��p< D�FmW���0���ﴣ=��L,z��ΕA�K��q�2�q:x_�t@)�fr���NA��yMv�H�
Dp��#aĖ�r
{Hyܦ������ڄZ=7�CX����2&���fVHXM�T�g?#�"A��q��{�BK[�
Y�n}>8m�&�u�0�T����|:�g�Xx��W�4�ⲳ�����2�>��{|���U�Ã�|G�u�F8M����ӣ��S�׬Y�fb�ԏ~�#����ȷ���<�6ƪR'��c��^)A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �"A� �F�����?���:I�������o�T���f͚�����I�"oY���m�0*�U8L�����ߡ| 
	�w��d*��Nq� �Y��,��N�~K�����P��W9����O�=�%������Ց0�Δ��~�I|�` �EWW�7QX2��3��?��މ��H4�����=����L�>o����F������>���?��>�`B/�}��O+���}����y["��y���|�]w��2܋g �9��;ߙ�	,�xޗqߋ9������Jeee-����kr�dff���_ƶ�8;'A5�M�}S�V�M��H���m�e�3X&�o�g���������wTw�qG#j�k�s��9��tٲe���@-Z�v����S�;�c�j�j�3xϨE���bm�#���qn��,�(��!��3�x�>{����@ayoժU����}���1��D-�U?�84�����/��\���t�����ؾ3}J���n�c.~n���}��������s�}��wF���7Q��E����X����$����{��<������x���C ����x�x&�'�ߊ�?E�Qi@,�?�nݺ���4~�/-���x�W`��{٧Ҁ��?�
�~Tl��c^���������������?�������^�G-�>�=�ė��G���tG��
��N�    IEND�B`�PK
     $s�[�Sd�%  �%  /   images/3357ace3-f4e2-44e5-8366-d3a4568261a9.png�PNG

   IHDR   d   �   �R)   	pHYs  \F  \F�CA  %�IDATx��]	xŕ��m]��[H�����������	�#˱v�@�K�0l��AB0G��c		Y��H�N!8��M���-	K�-Y��Ö4��_S5��3�=3=R���}��t���z��{ut�p����N���>�Ox�^�w�^Q\\<ihh�����T�Ǔ��9H��Rq-	׆�y��!�����lŵ�III{�A����Evv�����I�@�o�.�t��A���-� �������G�20� �!y�݋O�z\~�ۓ���T��=�F:��:�_=��g�!8���"--M���'�# iii��X������0�`���y2{?>5 #&����@i�@�@>��\p[���L�4�ddD����bƌ���H�'�+ MMM�&�������P/sp=S���U)�@2%?8G�s>�3UUUQ�d�JKK�xѸRWWGI��7`,��"HJ��!;��	���O1Z�
�>�p,~~��j�Ki56.��ٳGJFVV%�
�>��nII�/�.ГQF�^�&�D'Iݦ�)���
06���}������) �`��������ӸN1��8059##cvzz�0�Qz}ہ��p���?
���c��Ԅ�D[[ۘZbc�hllP�7	`|���_���,R� ���Pn6��\�J�����,J��zp|��^ؿ�vH�hhhb,h� �^�~cR�:�ť��3GYD��߻�Ώ��<��W�']�ա���2Xs���ƾ��m ��Ҥ%(9x�����Q�V���Y����DӘ �Ɛ�`@z&�X(B�����W�����ALL�qy�C*�D���(�:777emFj1t�������#����M	O�@�p@��륺Z�v-=�3�ÇA�<33s�K�����r c����t�*H�Q����Cz�@Zv��uO*�8�� � ʶ��GL)���޽[��`�X��|J��I�K����&�!4���C?q�.J���`3Ƌ6 ^�2fpC=��$\�Fg��d��y�~���W"�W� a�I���zȧ�C�hi����T�7��`�F����t|���Ϣs4����BZ��e���g(# � y|�����DQ�r�T0x��d�1�4ZSZ24�޸�������`��D���}�֣�G�"(�Pt��G�bg�'ⷿ�\�Rttt���a7%~Gq{-+�)�����`�,��P`nS�����蝽�88A�ԍ`|ڈ=���Xje�u*��kAy���%��%�\�� h"(!�0zJ=0���1jܠ^��]��8C&/u>$i^OO�Z5��Ed2@F�ل|����#}�>����� �*j :�tp�$��tP�R]A%|
d(< d(��b�=F|[
G��Z��N;�dI��@}�c�*�~
�q�e:\��g0�n�Ƨ@)b�E���B:�懈J�`�7�>W=6�1$T�������-���zN��-%������V9ф~��%��bH�Ef`xa� }���`ˊ�X��t�hG�?�`�
'w8��T�K����}����Y(�`���>s7QD8��9�&�M`[s��B��_i9� ��Q����#)_��N����&�9G��x�!���N���oKƶB}Z]]MI�%B��E��L��8ж��	&v�B�����N)�-'�H�S��tT�cD@�����L$zR�T�0�ٚ��N҃{5�V���n[ƶ�E�s��d:��F��0 &O������.������H:��'O�-S� �7o�\� f���g��	������Ӊ+j8��ٕi"<��"�����ԍ��e���c���F����rߎ;�2�x�6@��
���`d@���
k�3��<NuE��/A��~�d �4��m��p L��8�#=b�%;[/M��l��̧IK插HG
*�"�K��=aht�m��3�j�:�(G.��I��s:Z�yM��#@j=��+�h���`݄cjD��Ю��#[��1��8�\@F. #��i����]s�)�ЛNMM�O̲���?#�=�n�N ����/ioo�>9�̥�,��ԩS;Y�#w@�82{�ƍKZ[[S��� �iUUU�VVV�&��#s7m��ɮ��idj�{P^Jiii͌3�)f{�O�^���9{����������̀���������hnn��n��p#�䒒���G"�JFKKKQ]]�g^F�8%���� d7�{�5$��������>%e�#�{�^\���S�^�L t���n�z�סצ��S��m۶��_F0�$����[�hѢ粲��*JKKڲeˬݻw�1���1�`��g@_s���P ����Ɠы�k6��Pz���S���=7T~j���?�����~�� �0$����M��RQ�����֔6\��a����j�(" ���{�W�A#RQ�1�B\��8`*f��h�*b�;�d���wBݭ�����*��0ƭ����q-��y�1$� \�LcY������?[\\�f c�D>L݋80��I�	%!ѐ�o޼y���˛�`��˅��ppp�������A���ٳ��������I39����f�_������2���;@L�3g�|����F��d�[��4�=]KqX���A*6y�}���+��@Mr��ڵ_��/l9l ѻc�pn�bo�7�[��X����UF� dtYYYmEE���)0<;v����Y� K�@(������v먰f~mmmU[[ۄ �4���=j~�r�EEE�ӦM��`T755U���(T�k��qB���n����2B��N�zV���ei�C�0��R.�imm-���g���a~�q�=)�MS�L��x�bub����N0*++�<�������.'�d�@:=��5�D|���иl���,q~�L�f�0L>��1�.���3X����x��s�1<��/���;/�*�	 ��h\.R�x��8��	M�w??++�����.#(���wF]]ݦ��[�&'������=�G���(�8�1�M��뛋73r�AA�B�����/����_|�x���Yg�sy	��
��g��	�$�_����A;j���z�2�����|�3k������������sΉ������K+��'$A�EI�������2u]NG��n^^�_x�@<�$��8 2M��1���+�L����b�>c�
ұN�,Z�H���[�SN���� ��qc��k8���BE���с͆��	/������a�+b��v@(�#P�H[�':%A	�D�TK��g
�~EOO�uw�}�X�xq�۽aG(}����#qxUr;����!9gVTT455u�^�Z`��*c[����uwwg����7�S�A���Wc,9�����u��Bk���=�ֈ���p�Ou�t�5�erRGG�+�M���6@o9���S��~�-��<����8�Lm����9��S�8��U��%�Ֆ�Q'�Br
��.�jժ���"�A.��Z�ݣ�v�&�ҥ�搗�8�
h�:$Y�Q��ɇ^�e����p �G[[%�	�-:@��0�rI����a���ݹ��<����^�2}���*++k@�J������6��.J@�2᧌ �� ���i��"==� ����<eʔ>ubh�ov/����
���������� Y-����,z�ف^�Ɇ1���3��bU!Q�F�
�����|_,���{0��A�	ٍ� ����xM���G��ђ�f/+��Օ@W=@T��|�j~T������I��b��l�b>T"�@8����
����\�]4�R��b�*!$X%��3Q�T�}�@��p��ې��۰i$u����꺆�Lr�V ���S򴺂a����PB���R���� �c�Sѓr����!����ǹ+7mpp�*Rd:_Y�.(�P%�f)�����������p��2�[�	����F�`�`)ra��~0�q�v@�H�H����V���O��>E�XA�e`0Z.
�J�r��T���x�H�ʬ���H�C����C���S�4ED �=��Ԕ��׫����ؾX�DM�z H_��b&�=}�pQ�E�p���l�����������B/�N��N 2Lk3ZJ�.{g�{Db��&��9���J�S�N����-<an�u#�
�i�S]MtR;������Q2� VTT�(\�F�^�v��h�V?D'V�ԃ�]���'�����Kj���flOyy�w���R:po3~�+\e|/Z���I����#S)�ZsPg4X��xB�
�H0�i_��JKK�EEE>%5|���~��8�裣.�6@�9T�s�#�v��=e,���J�-�V�K�f<��|.ծ��5T����L7�?2Z���Y�f�T��c<x��3fx���1$ӧO�Cɡ�X��X�z��<Go�#�T\\�帡�s@��_ǵ�|�����E,d��N��b���:J���� ���I�w�O@�Q�'}(|�(�^ke��N��F���Q���_�����={vLuH��E�Sl.\(_J�����QYY)�ONUFi���U�`�!��1�� _���ӓ___��޿x�x�1�o��)ԉ(�๷h��X)��V��ā�ؼy����2��WɂW>Iy�-���<��~�Y���^]�$)�����i�s�dG���P�?�dp��k;b%���a �=�X�d�|Q1u+_�WQZ ����|���4[Nk�c�o@�<h�BJ�"��|�I:;��r��D�R���Z"�!z�]ź�N q5_Bi,'V���M�6u�A�ſK��P��fΜ)A������~/D|N�� ��78�:߇0��B3c9�S����^Vi�ʷJ��2R�E������(��	q�8�hE>W@*�����x��d�cHSoŊ�_q�)�����Yi�s�Ε�jll�%�۲e#�^:�L�� N�����siX����!����R����<�_v}R���:�#�^�n]�5�����c�"�������M�{챲�M�6-n>���d�UW]E'�V��<��5d��c�L%0 ЃF$�ܹ�gWѩ���D�J5�����fs�1���6.��k���ܸ�u��hE��ʫ�p�Ag�{},GL
Н �Kxv'�СĜ9sl�m�ТZ�~�ԵTG�u���\�����a�$��1t*� X�%��I氧C��A���f��DN%C�x���NZ�����f:�3�&�������l8����2���:+x�}�鳪Rkkk�7�����н��fo�2��>MI�n�S�ܶ�������A?&J.;5��3Ƥo:�~z>��.U:���\���;)a�w{"�].˧�K]KƄ6�Ld -2C�7�^�آp=fh��c�.C��;?�T�P��k�� Yf���X�M	������b���hZR"1�����c�E1٧��ƼB�a��@p�a������L4����T7k֬[�n�����*������<l�=
"��M"AGx��%�C�����/��u����'\:��>p��9�ǳ�+��B7N�v���i�ƍs[[[�y�p�~	���!�6���� �ڵ�.��@/j�,<2~:�/�2��ׇ[V���1P���r-������[���7 a���k���ݔ�U'��f��GI9�3�����oϟ??uժU���_��������D���Ꮮ���f�gH�	��6���Z�|y��_0x���f��]/3���,[�,�E�?e�V2���_\p���z��'�`�k`�h�]��k\W����u�v�B�N��QJ� hә�+�'�q_ەW^)���k��:�X���[XZZ7�p���l�<���qh�'p�x�m�2�����_��
TI&2���i�ԛ��v�e<[��믗�y��N:I���+�祼���OeRϤ/�ꫯJ��{��R�l!�y:�������L�B6����
�:�D��/��}�T���`�jBYMk׮g�y&�g�Ò����F�������2�*���|X����T����W�����-��w���~:�^f�M`�A/PL��GYx~%� @B䅟����;�z,����������r�4�T��Ȥ�ˑ~`����Nq�w�x)n@��4�,,��c�E]$/(uT�<�V0»C-�\dM1u��oˎT�Yx��dk�����=)�¿4����Ͷ������{�K�.�P\�P糗��Щ�-�e+aO���ӝ4T�^(��#P7���_n����E2����N{��hp0�(�V̺-�>9RiR�c��rH�e�P��x���AD�@�~��_����H-|�a���µ�-<��u��!y\�)"º��|����*L҂�<���X��%h�G���j��4n���o�X(&@�y��H����/����g�֎VWjP�l��[���P?(S������SM�aY�(W�#��F�A�!]����2��4ᗳ��7��-��"������c�����,>N������z�U���bera������{,���LG]6Q�Q��!��7#�W�5>=�{Q�
=e�v�x�"�
�A�`��+Q�G�>���j�4�|�����07Zq�:~	�������.�E*���b)E���m�IDZ�t��F�x�G��Lw�hA�3&)?��W�P��eu��+g�K/���t�M�s��l!��By�P#ڪ�5;�����s�K�AA;�����_�P7��q$�|=(� y��GM*��U(��u0���k|=�1�l�#qǔ����p3������0d1#�3����@f��ƝZ���Ht�fZ�-�.�u�:���|���Bc�Z8f<&L��0P'җQ��C��س�e��l>t���_"��{�e.#B���$|>�T�$-i�s�b���ː^�OS�9�7��/II�ko�O1���y�
]��G�u0���n{,UA�E�V������6��`�o�٨�߅&�����6:�:^#0�7Ǥ� =/��B$	��,��ie3��4XSW
�(ZUS4K�AzYǋ"�A�Dyr�⠕��q��A���+�$���:Sݐ���U�����.¦�Ϲ�����QX@��(=̊|YD�x���%��jU:��y�����u� M��RZjRw�}�+�t=��X����P_�����J���>���)�7��
	�*��B|}BDa���7�9�Cو���VWK�϶�m�]��n��v�@A֡.|��Y�����p�!i%i���T��F�-�~�e�ʼB��C�̞@�TMKO���
���ڮ���*�*f+'���V�x;�Vs@NA�s�����&�����������>��5#C�2
���\� �0ue�םѭH�h�E��ba��Mw������p�U*((�*@|��&��Qu�[������0T�Eyx�>a��˧��YP�ȧ`PFb���BzZ�炈��e��4C�`@�d!�=���pi�3�<c�Bܽ��3��^���La]�N�h2:���~��ѽ��O���{}��@t�V�7�p��!���؏��]30HK�d�����GE���[e��ćy �E�O����{3��Ku@�C�Y����������q���h���ۻp)��	�4�L:#�)xv��{����ђaE#-43@�gffV�,K�J2�/cK���Y���(��h7r,���*W��рh���5�>��\�,����Z�EzG-~�ATG����+'��������DF�b���b�n@����q��Bd�A�K�[��K�@ܩ4[QS���B��=��n��I�XN,�J҇ �`�n0۔��N/^�rW�d�eP�Y��$�X]��"E�<|2�j�u��i�>�1ژ?M>��kiiY`~�x����Ew�H����`�!�`$Z��H�A�spH��ϸ�5�F�n�s��-*�ι��X�q�7��X,'������b5!��3x饗ZV��ĭ�|�h��ۧA����ʂ�QDM�_��7ס�W���-<z��>k4 ��Z�7>B����)+�Xz�d�����n��e9�'��Ҷm�$���(�ۮ�"�^��5 ���?,�8.�EY_SS f�y�������g���\����X}D��q�뮻N�BJ�s6Ǵ��z�Ϲ�X��2n&�a��U$@X'JnM,e]{�2��j��F&� ��磝?b���Z(k%������iq����;��R;���&��M�(��4$t<�%Y��lH(?�b���:���d�`��-�S����R���}���|���z�RB�Y��%��=�gX��ɮ��VY�Mn�u3N��B��8�B�oE�/
�W$�K@���?�U��4ƂL���k<��h��t���e��	��:�k���Rb����}v�ΰҗH�v��U8�F�R��b�۵���*/��&yip�" f]���fn,+��$�A��-���%4���c���hu)���B��l[g�����b;��q�c��76
�o�e*���$�4��(�v�8Uc��x��v����D2���4"����2����JV�=Y��+W��.��)+<1 ���J��c����������<G,�|yC��~0�P�ʺ	��
��XY�R��r3
�c/�{�q
c$��V.���8�\@F. #������a��0rq��8�\@F. #������a��0rq��8�\@F. #������a��0rq��8�\@F. #������a��0rq��8�\@F. #������a��0rq��8�\@F. #������a��0rq��8�\@F. #������a��0rq��8�\@F. #������a��0rq��8�\@F. #������a��0rq��8�\@F. #������a��0rq��8�\@F. #��xP��<��ʕ�x-d4,�+��|>�
d^��R��~"�@! uH�"����z��a'!��f�����fb�fm�R�(�d�NJJjſ�n�' �D�7�M�'''�a3=�tRF���c���5�\wa�����W���'��:��f+�� �y|�6�m�LA�s���!n����T$�P�I�,E�)5�=����o�d"�����%�˂~Ruz/����¯�Nq�S�"7�?W#����J�6$��.��w�|�ͶV�	��'��z\�&�|���&>�!}���%����<�L��7�s&��L8��H��Zyqd��!��S�َt>�MH_D*D�H��ԣ���K�"��@�    IEND�B`�PK
     $s�[9&��ސ ސ /   images/b01488b3-8551-4b4c-b09f-2812c4acc168.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  ��IDATx��y�m�Y��=�s����n�$�I��� �1���0(. U�D�	W���T��
�+�JR�#�B�Bʩr*�+�	6�6�hh���o���{�=��o\{�s�{��H�}��^����a���^��}���p8��N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p��h=��?���0>"�����0<�޿T�fS���bߔC�S��)�P��� ����e�C����0x`(gu��]� �(�X�_��y�����<�����:�=B�6�n���7�k���S�#�F�����S�1-0��!$�n<���!��`(���x~��'�����'�G�iX�s�q�8����:��q)v$7���GY4��1@�a�נ��?`�3��`�G1���3�����|��(��P�����ʢ⯥�(e#�]����eXq���8�W��&��n��g�^6���"t�����fq}�4��/������;�M8ٟ�瞀����O�(��p�$���yL��&�PA���-BꊠDO
����La(Z��g<�0Ȝ������I}"ţM-�I���\�C��x1D<���ؾ�,�"���U��_����>��W�7O��'��W�c7��－�y�������� R����g�H�7B$֌���fd�I���*��@�7%t2�}��|�W&��:	"!j�X�c$~���(�#l�bn:n��kuh�$���y,g~Y�����?o��oCc�F���YBY���c��pp��5�[Bo�^��|�vs'Oު7�/��>������?�R�UH�oA*|��Ȉ��;��0G��HDM��3	'}T�v:�lRO /o�g���q"�ٕ7���Zk��'�]�z�����>�=u�*Y���(��TAQ�ş�Y��+�>9����x��py�W���~z�Əݽ����!v_��Ư��T�8��:�e�����P��'mQfDr�^��L�l��0�Kll@��,�&���Mu�1$��َ'R��ь��ND[&�k_�Ch���{=m
��a�X>���D�.�-*Mź(ʋ0;x�<{aYՇЬϡ]�C}p"���w��.^䟛faqt\��_X޹���߆��N4���؟�l��)�u����	=z���S�(�a��<�ؓ	�I=�p{�|�\�b����d�X�]#y_¦_�r��
ϵCR�c�z��MQ�]�i�Ԋ�ҡ��B�d���U������>��!��������~���~i�6_��)��;��.�K��O"W�����ߌ���)��}w#v-���]�$oB!�3� �g]�0���zg�"Z�� +*�&�_
���D�7E,���dGeO>�<{�˘�b@��|�Z�->�	���2���3h��iQ�!��$��ֳ�����_����� ycI�8�u�X�7�N���g?K����N��=��au��hѾ?��si�n�^X��"7�B�L�=��T�t�2�ĉt�
�&�υ�)�moz�G�'���}�B�Y�MS��-��;G}	�8�[\�C? Q� ��hU�P��]ࢤ+ ����:̠�j<���&4q��0o�;��{����W~����?����O���_���p�Ʊ�l�B^-�����G��}ٛ�z�����}�M���[#-���S�dN2eM��@Y��q�o�U��	�D�!LB�&����׳+s*/�GCf"/���*���ҔD/(8�4�ʲck�,��>��~����
��?E�����^���������_trl/��ާ�Y��)Q�=�������8��Cw���+=� ;&Q
��ԍy��.T7�2�q͚�LD��1�<yF7�����~6�ϳw�>Ç�cH����Bo���*{�$�t}M۲�>�WpPԜ�W��y��Zz���",XC���� �1�z��_~���������o|ӗ���_ï�*@�� ���|�����c��ɧ��}�bx��x�[/����E���4ϴ�͢�܁�d>��B���OT��s�|������T{yޡ�� I=Q��š8LeQd<��s��)M��v`�<���Y��c��kfܐ�-J1�3=Z&(�Bq���1��W���Q��A�gB���a�������������z�w�m�\܆fyN�z���n	}u�.�G7`}����3T[ᤆ�����G���}�Z�5S�ؔ���i�T�2�坑�w�'#�4e��N�d�����Q���s:�l�����A��c��(���s�G�������5�����=���-|\C�⍞�u�x�u��妄��jg�c��?���4|?.�_/����o�\U�G��ߋo���!�m�bq�&8��?./ɥ8}xx���bh\��{��~�����v}�n�7�A���j������	�4x2RzT���e���8T�Q�D�/�EٱZCs8��CR��A1G%H��rb;��l�d	[ϛL�OL���А���E���/�}�(
s�� m��#��b�F$��*�j���gc,�������^J��1�Q�'/��Q?I���g f�NN��}��Ї����'��_V�_xk�^�N��}kHm�3�'�h�B��$nN�	�svy�y;2��K[�r������F�<�t��B�� l_�&��ߨ��]��ʱ�4��;�i�Z|o�E��P���z*_KhŇ�-��H�ҕP�ڢa�K���b����g��{CQ�VY��)��o�bY-u��Q8�AY�9�@�7����ڥ� 	7�>����n6'i迹o7�o��˴z[��<�6�e�������	z^)���G�60l6h��Tw��xǖ8���F?�Y�%�n�A�$�Y��s��4|���i4L�dː7b�g�C ��Kz_�qx�z�� �TbB9E5C%�������v��墨>Z��C��̓�%~�N�i뻟���m����S��$��K����@<8^\���7�����o}s�̆�eDm�Yr�h�V��G���K�ʄ5�dYm��YcM����!�v7M�8M��ɀ/�y
�&|O��k�U�Q�je��"f&U	��r�kv�G=�.UH��hS͵�TO�%��~#�E���))Ѯ/C�>���7T��+c5��b���P����Z�Z]U/���;�=��Ւ�+�����.U�5���
{���E1G���gp�[����a�~6���0���$^�+$�5��Hͮ�'�S\����f��ް�=�h��:4С�,��Sw��s�2�
K�� �x�2����4c���ו-{���L,�P�����Q~����N�1�8����$��
�����TTo��_L}�eU}b�����8T���'O\l���3Y�A؃d���_� �,��&4��A��g!��*RW�0�Q�S�Z�du)��u�gk��S�q)M����m��+�l���
$�d�v�ZP6�'V|B�.���Z���J�8U����)X����.�"zVf�R�D"�Ԅ��ǥ�0P(fhЮGB_�tX�(V]�Gl�B[?W_�ٷB��nS�ˡ]��jV}�(��P�m.���%
�ri����r8�]�..�Cc�������e��ě�Q`<>��������ƾY>74�[�YU�6�@"�e[��_Ė��+�=Z�d t��54���{�k��}�V�F���뇒������5k(�K��U�q��'Ƥ\<&��Ul"W/F�}�O^�Tc�e7K��*s���à�����!s��9�/�e��{YY*��G�}kY�~��_[����Vy��G�7�������?�g����˟�xYΟ���c�o2u�[ 6���:��Բ�(RBG�fR��g��6��h+OB�2��Ěφ�Y��^׺�ǔ�L�di��4���L�$|Mnw*���D�F���E�"'�pգG���"��H��S7������c��E�`SA[́lzS<VE㊦|�T�SE��[U�R=�J��M���P��7�v�X����r�D�s�������X8_�`9�K��-���m����OR�^?�L�>�$�o����Ϧ�����9.�%�힓l{%�8l�:O\���wQ���m��(�sȑ��{������oт/��·��K�P����#^!�%O2��v$�6�[y����^N��CN�R�~�=���
�gCk�X;�zM�KB�C�R�}a�8��q�}E,���B�+G��_��x�O���J���߇/��y�ʬ�����	QǊ�T׮~��6-���&���)W���Q�b	���q�	��p��P]�{+ήnQA�N���dr�4UR����̭��&�WRIZQ
i#Y�r=��]at�U 瘞C���v��.���E��GQ (�G��0��.�es���^��t=��~��$�7AW�	������������hj��)��Op!�A�	����⳱�s�֗\N����1G�5�hL��m/��"\\�`6;�cjGIM9�)��NZS�Ã�r*���5
D�o��G��J.iLI2x#E���H=��Fi�"SG�rhg�'b!U��"{)�K��(�|K��<���*���Z'
}	%h��%T�+��J!�!��KK�Z�75)Ih��4]`F*$��>pl�M3���1� ��nA���ֽ�3�:��v�SCGCU�ۋ{Э.��7Mz:����ͧ���w#�7����U���,���q�yG��� �w/G��m�����^�=y�^�	�������.=�A$s�)u����~J���.�%�'�P�D��c||�7$�')Yk�7��ŉ��ҵ�U�+�x�HO\�(M��>Q�ܩ�m��B���Oԭ���j�]�Q_�_�V��b�}�ŋ�?.Nn��o���]� �W�.}y���Ot��?Em�CH�i��^<�nٔAK4̪6�[<F������;1e8�~鉻
s&{&�4#}�b�*��	lY�y��j�LT��Ob�at3��9穓`\CC�*��Nϑb�%�コM#[�ȝhus�	+ 2�;�̡���Հ¹9�*q+�������f�~>���jTZ ���{|��Me��T���^@��Xӭ>����������"�#���>��~���o�!^`���?/�"h��N��-h%�o���p�f����};��ia�p�!A7����T��,J,����8���������3��JiV�+��j(b���yR�xW���*<Ӫ$������ U�D���Vt��X�&8�(�K��	L�ہ��}4eT���� E�Aˋ��S��L�'�n
�q M>���}@8�%4�X��8�ė1Ц�������!K�8�����#�@�%#�p�b��CH�Z���[�D��Et������OǛ_���m��%8΄�������
m�F)���(���X��e;	Ք�Q�����y6Yش6HK�y��vu�2hv�Ϋ�(��?��|G��Սjv����Ko��zG��[`�<�Fǭa�c��s)J���*���"�@�5$�~#�nlq��C74���$ �+�*P=���\�K�i%lG�[P�-*���ch0�([P|���l�	�4b�Qz{�;<�2OM�mgeU]�v����L�����0Ns������
c�R49B�U7<XI�2�4��������x������/7����۟��7�^ox���hKU}p��\�5��?����C�.�A\O�ՙTlEP�S&�MD^�,���gU��L��q�#���u��|�Ŵ)ô=�	b�;%i��x(��z��'V�P����WE9M�R��9��Pc	J$�|�K0�ǊZ�ThTs�[�V*L�����S��'7`�EBm���p��[�(����CYm����(6w�P�����S�� �t���(=5?8Y��@�n�$�i�:P�O.I���@{�T����gI���+��^vE������t��~��3����|3/�^�u3���F*��0�fժ�JT_�<8���}y������Ev�HA-K��Ʃ��yE�j��!�4�5��B�d��%]���i �<��YJdr	����F�sx��-I�Q �E���j}F�ވ�2����.=��.��=N)���+���ŀ����ZS�d��P}�Cw��g��l��lx�?��Ռl�A�][�����csA��k0y���{.m���E�0L-�c�ln��uwq����@B��r�Z�7qt���i�c$��YH}U��H�MV�X��!b�M�"o��K-y۰E^�0�͆Ƥ����mN�|O�z�r�<{sHq�{N��z���<���th�]���b���J��Ē���s�˱u��EӺu�-o�O�{���4d%+�B�%�E��vgҤ�|ҿU�/V����-4qP�B"7e��!?���U��74է._�$?�fx=�5K�tcW�}HV�Yt�����8C߀��,����5�g�O #tB��'V�ul掹jLf��>���.E�>��t�M�&�������QH���ļe��r�6�
�Q[>D">��9#�flٍ�;�%�v�,j��1�GKl)8��-�9����dk��Q��l������([3�W������v=J���k���`���;*!)��)2��Z%�u�h䆢���] ��~��ۣ5CjyOk�%�p��ف����ʒCd̗����"�Ч�bٔ�.6Ų�l���k˾k��l�ȁ6d�H�&Uz��"�21�j���z��I��J�t���xYx���w��x�B�4��l���ob�?�d3�?�<4����s}����(��'ǹx��5yTe��R��s.�K(.聆9#�;[^�ǁ�5ȓӓM%͐X��yE���Ef�ܴ�<=����0Q2%:j��s�A��@�'T�-B�J~��N��ZU���J�ޢ^�Rg�70�ȑ/-g�8$�\�x�^W��ѲB�'jr�5(p�0�RoFT�bI���X�{����(�ltD�W�V�W͠���kMu�%-��#B_�E���]���g�ZVG��X�ְF�=���C�A�_�Vܧ��,}���9��H�u͊� .�S�t>��}]��NaDjޠ�49�Fu2���&��4�Iq6Y��ibq���ۖ�p��gV����s�$���-��2~�䉪>�ţ�����۟�q���o��^��~�����p���?�ͱo~.��/A���Nz�v���g0�1h�7+	��;������?u�g��>:���6�uu_7k}"6���|��C��,a/���F�Q��g�`���:	�����2Ֆ�G�u�J�2d%s8U2�q�R}z��Y��G6�uZº?��>�cΔ� @��)ǥHj����\Z�P���λ/�%�$E�=�Fu����b�V�*��`=����B�r/ǛJ"v�[�Ҭ:8�����{�Xb�s\?�h�[�鉧C�FAn�U���8�7��"eU5̩�.�nG�pX6<�7�5{�c���`R��G%1O33�A����{LЎm�E�~d������Lb�8����\B����v�g�i2�3�HF$}����1e_Ǎx���	I�<���k�y�(g8��8<"��<�y�1 �I܂v.��c"�w����KRmjua�d)����L�)�6�ԇ��ј��A�I�.����������V=��q-�R��zb�ʥ�jΉ�I���y{r���GŊ��΁C�(�ig>-y���]��;e��\�:�~p�fu�2�����i�DR���
�x�2�*y�E��bY�t�87��jr@�l��"��UPi`v5���x2�M�=~%*�ܶ�G��,�8��ʃ��u��CC(���?�w�N҇/�K8��'�����k�YB?��8{����L]��C�|'��L�"(8�&%jZ�6�Z�I	r��u��f��<�B�j�$�C��]w�|턩sm�������7����ط6�2�(�L�L.qd���:�*�P��d˛�v�GV�y'���=�2%������hL��!��(#�f)� �N�0E�6�,o�&`�{�W��G�����x�D�J]&l�d[ઔM<%��� ɉ}�*���� �h�������8�'NR�y�)o�	d� �h��o襱�0��)q�
���0��f�r��Ǆ\%�����vϓv�ں��oד�u�J�L�{g>�Jҕ#Q~�6��X����y �q�BB.`J�L�ڈ�:�u�ذZP3�R"!k��p��Ť�1�2�#��<~�bmr�&��8�e;�n�+�ΪL�ۆ�*d��*�kR�C�
�������Z�c�N�?)�9��>������	b�2M���i�6�߆L�����$I�a��A����;�CCV���%,p<o�AlDAExݒ��Ĺ�"���&��h���y�D��d�o��ɍQ�]ޯ-����0����Q�C��U&�.��Iw��-dW9I��_yi�e#��0Gq��������+��#��C��?Ã?7�y���$���6\����=�u��5t���~�+����nZ��y����!7]fi����u��!+����ֻ>l�),aG�ؙ`�<oBhT.$l]�8)IB��9�}� �������vr�L���g�8	���X�d�r����Nr��Җ�k|�vu�mZ˨J���lM���}��vT� �$&�tY`�.zV���UL�)1+@�!��Uכ�|�����|)$5��0h<�h��!������Ȥ�K̙ȹl��9�n���:��,��+A�0�2�HH��P�<�u��<)��nv2a��3ӕ�9�.�_}�x�т��)�۱F��.��Iց(�EI7�7Z��
u�KTA�6�UC�=��� �y��Y�cR���2�6��7�f��%�ާ���9.u$J؜@�
�h�$>>%0����ш�5mLĥ���L�ٚv�?��37�ƍ!���5��O��}�9{?)�z�$L1���B�A�Y�Y�4�1�5)U�;0���\o�
E��>�آDc¢��������̲mQY��@e�I�^>�y��QǮ���#������&H[�����<�V��g��D�b��0=W>Q�#~��C�����-";�Θz�UF�KF�!��ή���s�O�{p����~�f��{�����=88}^�x�:�(��w�C���ط5vm�xs��\�����Iv����4G1���mR����#׶j��aO?��8Q�h�{����p�b9���W���fVi0˗��Iɐ��%���Y�|�<N��PE�s�Rd_�T���-WH�����K�����P`��	���/ �4ٶK�H�E�{�QY�1�@Vq �HQj���+��� �|�t(m��k^֯_H�v�����
�yݣ$���:�wڵq��,IXr��ĻSq}o�jr�Ib�t�d�(<gh�6�@���*H'%,��%]c�O��qlǡ	ݬ��3��ᔼ��:���f�lW��9�M��ǆ{T:��+J$�}䡠d#$�yGLJ`�~��$v�:Eb*��(�q]s~G�]��2�{$�~]�d�n��/D�`y�doX&����׷eM���"0�$m2���a�l.�4~?���]	Ƶ�Q� ��Х�T<@��`
}��<����2��Η�}��#��u���z�U�=�K$���ƷCI��0����`���q��YwR�T	�J�I�@9�����DCi:�Lw���ԟ4Z�F���`��'�w���?��(�ā����4E�����<0F�9��e�)o �9��bhP��,����N�������S�-\�{�_�h^s�~��'䗪|��=��FR���9���K�XdWyT!i�y�u���}��'�իߝL�f������P���t�B�d�T�C~�]C~~!���S���ݎ���=�ɽ{��c�x�cB�7P�%;p��ě����k�E����s<�,����I��}�ǭ���6��|-�`�VJQU��r^B)K� ��qU�`u�I�ˋP�n�D�Z0z��0�:+�]?�}� ���]l��͠��������.��;AÀ��J�`�I�pE�>�"�{{�ٮ`�lН�����;�V��Im���y�7ޜ�i�ز�NpK�n��晓�se~eRR�@���&B�F)�� �p��F��T)����LHj����x��B��ۥ*�B8�^ݓ�D�³�A�`���{$�ް`'��f|�d�R�!�.�/�Jr*f8�G|CJ�)Q.T�F�0��q�ړ�7{�tM�ˣ���[G�*#9��ǁJjTdC#��$f�\�Z���n��%��>*	��wI#oܜ�Y� jؑ��*�EI�B�����~]!7�\m�K�-����oI��кR��G!wAE���ْ���e/�$Ĩ�y|�
�K���$1EP�sZ^�Ī.t���JGCP���Vu�����`
��+�,s0�m�\��s��c��3ߏ�NGd/N���P�)����,�_�����?�6��x��5E�ͽ�x��>׵���������Nd�Tj2��%id���T1J5~���
F�hIJ�����,[J��Z�8
L����M6�r"��%��k޲��T( 'k���#Yδ�6)]+�})*�x��+=_�Z��,x]l��IL#�r�_@�c��ڈ�����ńD@��d��b&��"lT�l5�R�/���c����T��O��d4��c�(��Y36x�{R�B=	�_1��!˞c���7�&�Q>=���f�ӸQ)$�"h�����ɅD�Q]�����Ċ!9���R��f�U�T�;���z�Y��;{��Ė�iĪ�R4�%_�xL�{=G�b4�F6��*�T�T���D�;ϱA�օPeO��X ��G�b��B٢`�)y����-TցK�&L��57[@���0�D��I>��N�Y����4��n;�q��_�,k[yT$�l����MB�1�_?M�5�a:m�&:�������R�d]!+���Fj�ˊwQ;;;��2ޣS]��^�ry�M����1��������m�u�� E���7
+u�(�h���9j�<+w,K��8?�B[�Oy�<s�^ks�5>yЕ8'cc�%������a/�:���<`	���l�S�����t��i��-����q.�7���u'��2�'_{���f�nD{�e�f��zy�7�n��}Sp�����c�w�z��MsY��MH��hxbL,��X�8fB�>'G�J�c�2�V�D��1̮��v��Ӟ�q��4u��B m���^k� �[r��SsM�E�D ��z�->�	-�ܩ|"���8�nJS���,��{N�+E�%�fn9I���P�`v���s����������I������4�Z)��M���}�������tTW/)7d��TaP-s�,sj��콒$"���(�%O�E�DN�&�����%Jee�x'�|ÄP'�G�U�{����X�%K����O���)����tUm% �͓����=�<_�$9����=�2@B)��0���m��n���B�����Q�M���$e�v��4��C��^�($a�/vyvY֮ t�lO���{�	�#�&I�N	����z��k�pDi����.�CMbp�+~����I!-�8�k;RH�H�TvF�c�a�4�|R~����@�����8�/��]�?kT.���v�H��������۬��S�zY��^��&����DS���|�܃�(&.x́���)��c���C�=7@��c�8�01�tE�Q^�g�r ��is�K�Gp��������b�����^��zp�f���o���� �͇n���l�Z�nȚr��e���(���M��Td빘X��\��DI;�6�ѻ#�sc��l>=�}����������Y��.+U�j��s�09�-�(d��(�rW<�a���@��VzB!Q��~�%5����s����V1(~�wgܣ��ϵ�!7�$���4�萳�U�N�����o0m];ř�`2�\�+{O	1G���H�G��a���$@Tb��J�8���bΨMb�Df� DRP��Vt-�?ML�R#�O��j!��-�o�����t��U1�٠36k��r�10�%�`����kdKx�8�(㼘(SI�N�:�dd��#�LÐO��f���Wa�?�4��#�QY�<�()	���ce�TE��5���d������\��!�I�l��%�I~�����X�۩I��\�@�_1Fr�!Q�>�����\S~y�����*[W'&�җ���6��#�w�����j.�a1�s��r����c���]=���Է�($�Y���mzQ�Ed<���`�J�G;��4giz,;�Ȍ�呻�}<���J���HBoAs�ݖ�)1��`�n��R�F�5�h��#�!\���ǎ�^���p�����ٷ�k�:���w��\܇/������Y�x�g(�F��ҌAk�q�s�{!�s���X� �$�]�*��t���D����^����f�I�qb�G��t�Ԯ$t���&��������[=�vۇ4�,`V�udbˍ]TI[В˽�ul�Ak��]-�k)�T�f-�,�I��� ��X�n6Ht�l�*ۻ��a��X�`��Ⓡ�'j)bN��C�R;kA� �5[#�5j�^�GU��yǥ)m��
Y�I��iY8[7<NG�^tb�S���%����(�@�f+%p5mtC�XQ��`�QJX6?�߶��D��57�LR!mϡ�0h9
S���jc!�dR`'
���S~g&�a!W�tb1S,���Cz��Ф�ˬfR[]�|��<����v�N�<!�M�I�6W���Uyͅ��!_��r�ZW��b���I=�)�Y��N�y��:c�rS�t�ɱsK�k�@��g״�W6^�A\�F�D�k$݊���Y��Q{גI�Y�q�%����!�z��BR��з=,GLt]��K<�j�\ӆ.��o6|�y�dx�뮥nN�qx����ֺ�~�I�*Iv<�����!��v^7OȘ�d�J�@T�9d���C�ׂ(�A�6�{Xv^l�g��&ޫ��w�ò�T�x�p�̛ᵀW����/����E�'o���?>��o�\��ɎBd�s�$�q7�(�7qU����Z����	 �I�:�^���0�|��ڼ�xcn�|�te-\�I��+�8�K��
"tr����ރ�8�~��2Liܖ5��!M��T5W��%���h���!�����QM*w�Ӥ;w+��3N����	mbB��]����l��h�Pn��G/~G���[-]c��>���bΖ��:\P�{����4P��>�$��Bզ�1���Y������e;�>�Y���\u'�Q)נ��8��+������ܘ$5U?mNZhŬ�Qh���Y�[����?m}l��f����x*A��!���D�Ĳ�8ւx�U��L�)�1k�@)��FY��j�
Mw3�I��3�j�y�-C5*�3�&��L����`� l��0,��d/���'�S��Q�7��}O����w�LTe��S�y�͎P�#b��K"qT47���T�V��.���	�ᙧ��'��{w���y�՚�?O{�d��B��:�i�z��3���Y���.���d|�qMoW�����7���'�P��jχIb��3��d�e��њt-��dI��/5�81�?Eq�.>�o��2~�����o�O=w��[x��w���W�Щ��ʃ�o��woo���o7({�}&�ȍĥ�V]�Qj����8��,�rm�X
�\����Jj=9d�i2�¨�e�|2�R��_�l��oyH��X�K`�m�N� mX+&s\�x=U�r�<%�����%�e�_���(��L�n�8���5��%�[6j�V�D�ԝE�QR&�1�M��#��"���P�7meK���v-��ɯ�ތ�}�ݖ�7����Ę,f&_3��������"'XQ�{ ��A�=c�-I�q�2@�޷�\I�Z�=
W*]�{��-
�
')�P�6��(�Fʯ�-
ZY1�����3Q~䦎��}�rL��5�ig�yQ�[bʅ�-��5����g/j���9�e��鐅ɒLXN�
<�Dh*��v=��(�$S����[���EU`Ұ��?l��y�Dɥ�1���b�rh�s���g����QT���є�`zOG%i*���J`r���[a�MY����P�fL�D����pr�&Z�K� 97�l��ԭ[h ��Z�=����3���{���.��p�\q%G�JYŜhG����RhF�6Y��ES���>[÷c͇��c�<
���d��=��M16��{�c*��c?���`��Q��Be�$5<l>s� y�Iߧ�L
�7D����������'O��^x-�U#tv�o������m_�5_��RO;�Q�f'�M��7�NpA��<���G��jN�R35�tڈ�Z��L[�����/�V-{\C����[�����ld���Z̠;D��s\"i�����O��UD"/�he�`1H�N���UQ�1�'�&�c�A2ԣ.�a����%Bt�lQ������aɄ^R�
7��x�k�AA���Q�(���ZT7����\qY���e�"@�ՓUGJB�V5�)&������1�3��I����T�D Q-�������J��VT��������ٔ %4od�W�jz��M��,xR��ͥ�~@W�O���x�m�C���%}'=�A�������*ق��mL�]�Ģ+����2��Z)��YK�y�=-��X�h�&��������F\�4	!XPG<�O�X�k��LjB��vO��(�<`�-�9�ӝ����)A�[����\FK��4����� '�qITUq"�Q`	�A��҂��ě�|mZfv�c5���1O����w�2�]fǯi�Q���笔�=�s�5���8V䵛�`�cՓ!T8�y������§>����wh�p��!\\&h.py)�>��q�KN�f�a��=��������~�%嫝3�D9c���O�	J3����M)��@!�v0�WY1���i����@%�*��}���j�76�O�Y�_^<��Η�=�x5�Z�;/�;������b���D���v��`z%���C��'��\���8Y�r��(�f3J�#��Qdd�2Y�-�h;NH�W��f"��=�	�+���6&�lZ4�q_!�N.p�Bk�B�po렞�$q�a����$�ʽ��I��uAP"_�;IR;���%4�x9l���P���v�@��%o�BǓ$2�(H�uM��cCj�e�m��kzKpduJ�a����L���&&�F��%J���-�M���v��ڴ�EU�L&tRU�8[���H������*o()Ǩ����#nI���\$8[Gh��̯�cu��i&�:��X�ZrBT�\��m�e�F�+3FF�ºB�cP�5E�@�Y<�kŕ�'��{v�Ǚ䮔��{����9�y9Ve�=D��7|��E/)Q8��+�y��l�'�QJ�����c���L}f�!L��S���2P'@�܃�ʥ��p-��(�SE 4AQ��wjmZ������$���������td�^�8��
��^�g��R�d�/8�������{د.���I|����x3�Z�4��,�ʻe�cA��HS���:똃���7k�����k�V�֘e�H楄3��Ys��cE�$�a?U��y6Ie����ݑykk#��p��S�Ǔ�\J�Ѐ���*�G��-��O�x�/��w���pt�Yx��zsvNN�~�� N��uH}#��P��h1r}�F���8�}�s`����Q_�w	�Ɠ�'�����p�[JȵưM#4!�b�[�����F�B�R�7� j����L��6)�2y��UKB���5��� �orC?�|-�5�)�v;�C��5[�}�HW5�4�-yG�4"9�5�lr6�kK��H_	a���&�D�a�5,����B�Z��m�v��1}�Ĺ6u<�en@$��ErCJ�m��jVHz.]��I��8��cŊj�_:kᅳ _zZ���E�q�z�t�/�UO��7����2w= 0n���jb\���|DZh��-JAR��֪d��G�G��[�!}"�.���$;���95H�L$|���������k!��S偽7Ɖ�l�p��8�2 g�ш��5��nZ����$�ܒ���~����nP�=7˱n��a>/y�ɻq�8�c��ɫ� ɯ�+���a�����{�����P�A��ީ�%XR�=��R(1fz"�
]I��Gͫ��Z��>okc+7��q]O����ŭs�[�%�Pb������W0S�Q�x���~�o����'�O��77˗�o�1� �^B盱�B�9{��.�o�7c'�9��i)����Jyw���V�FBFw�#0�~�q��ݷ^)B��M�T�Oj�(��7���T �h����Y �WJ��h}�E�Y9���
s�r�`��	��� 	.I�<m�B�z��*�|��`6�Z�Գ�w>��ۈuS��{A�|�E�F7t�^uɤ�4�
&�^]-f$����ȵ'q�f�(j�M���7!��J�B���Υ�!R5�^E'�Uڝ��������iܼ��2�^z�����}�n�"'lKD�g����2���``ۮ�G����5�$����1L��
6�7���8�M����/�t��9���lߛ��R�V�J�R�/����"����(��܈֧ݮ!f��zy��B��غ��eO\�$�Uz>�M����څI�O=OI��^&�����[��N��� JIp�g=���f�
NN��`�d^�ť�w@��е�T�6dE�&��b��_��h`�l��ym��� smnM����d�sK��9�۝���������5����W@KC9	���310���"c̰�r�Ʀ%�E���J}�U�Uku�S�|��?���~�s�j�N���]��>K5̧(x�߬�<�:[���9��d�jKCޓ{�^����7QmL,�.Fbe�MҰ�x�+o`��R��8=�� ?�g�w�W VhT�膤wS�5�$K&I�iސ���9W��.b����ӽZb�e�b˴�e�#Gv'M��K�:ơ��s)��삋��Ye���Y��uÊ��p�tL��J��y���Dr��ܥ��d-��Z�K�;�d��F��j������0�OJ]8E3Yon��q׾P�yW��(\�o��O$fg
�e�@�m��v��~5��h�
�]�`�����&!A����JMi�Z,tS��Q�n[2_C�X��e�=|��4��1����⍽z6L����#Xמɸ�\����Ҵ�_S(&��C>.�<�sV� _��� �W�=�&vlK㧍@�gcYƿ�9���1�
��LZ[k$�7�+�-o
!=��㰘��Y<�ٽ�R�f15�w�`��o>�a�Y絜� ��\P�6<B>JF~�y���^Qv��;߷�I����5z*���VVԜ�2��B,�>I�d�=��Fϱ(�]�C��R?����ֿ���\��=_�M\����߮��ˢ]/x蚿�7���mX���ZXw?b�,��d�=\nA.@�`$B$׹�G�\ՌU�]gAoY1��)��?�zVi`���e����R7��w!���F�t,g�X� �	iyS9�� �z�`�B�]�TW�}�E�������Jv"���8�t���s�%�4He|��D��yC�$�,�Y�W@ز�L��b3����
d��`�2oՆ#�/fg�{�Ƌ��8�4�D����,�l�XJb��Ś�X�i k�K�vڃ��3xжp�V��&�WD���5V�5�xW��Cf���ˎ�%@�H,�ŻA���Nj5�2�˅D-K�d:Sd�e��}[����{�P��M�A�zK�"[^V�8Q�lL���9���Zq��;M��Q1�މ1�vW}�q�5u�5�M�� ��=����=9fP�6D����w�w�	���)�Ԝ�m������'�C��%~��jV��Bߺ����{3,�h �ӎm�Iߴ�����D�Ъ�]��E�:O��t,�*�Y1�fM<��d��f/%+!��^J�r"��� &���5�ZE~S�]��șh.w�o$;���M�cE9�����W��V���?;|A	����7��+a6?��]��Y>N��ҾɺI'[�)�֨bK�BIE� 6���Y�[Hٕ9�Y�	Q�R��mvZA�א����i�^���n�3)с�C����DpqM�$i�媺��ؔ��dRW�-��I�u)[��ЙЭ_�N��]R��.uqXs�$MBt���*ĬJC�w���7�'�\�㉘b ������A�D�f1+� ���Ж���bҽ�)9���&���b�Iw��)f��'*g	��W�]�pѯڄ�v�Ǽ
땐���lܵ��<rz>z�N��e��Io��22�;z�;��=��u3
g���[�׺J�����>�"(9!e.5��q���Q�*��[�f������k���My׫�Z�6'caT&s:�T����7(��|�jS�y2�('.xs[v�g/����
��bG'��#i�~�ʣtB�F<5�[3�..a���=��S\gN��ٽy'�'N��=�,8==�^�FZA���p��1�+��	����d{�\�&��^����Vr�����+%6M����ż�ܹQ����s��8��,T�q�GjPV%{�����>�۱��Aw���܊Ο=�`��>?�A��^��'C�~>D�s1u��7,�j�LV	b�V$�/)j@�.A�����`$�m-������B���y����W������B��ꦁ||�V��GGv��Y��Fi�ܩ�O��2�M��g�'�&)����ִ�]�T�ɼ��7m�J�mM�`�voE)t���D�����nd��5O}M�U��h'�<g�j"|�u��FO��_���Kq�L����ͪ���~"̙��$�
*y����8&��"��Q2� ٤fVע0tH�\Y �O5H�ڑ���6��yr�u�ǧ�E�T��0q7�5��O:)eK]U��9>��޾�z�$.֬�ۢ��k���5��%��!RzO%瘃�:W��k�֯��A�%:$�G�'�v��C��{-+U�,���q�U���my�;��߯S��ؓ�ܾ�w�J�A� "_��>�
�ɯ�s��K �1i�
��25�s�|�V���N�H/���baW|�e�{�̏P� ��/pXpY��l��U\��� �����Pq�Uڿ��R�k���ԃ�L�������mu����2�?���J[1�Za�'��Jr8�\$�p�y���H+�,TN�ᨖy*R�\�;\Փ t�,H3�����ۼ�o�-g?�V��yo~z
_(|A�k��(@������6�ݱojj#)�C�G���	���ٹC\��9�eM%�����ė�T��4�['%��Xr����c���[��M�W�9d�`�����抓�"�Zgk4e��(`P� L�)�ߣ�1��&����d�S��
� Tiꓩ�6�����k��6*�};.$�.¤5�J6��R��JB��5*=�6��v�|�Il�ܠ���}��yF�\$�g��u�㺃YAЈ�*�</Q;k=
�V��ӆ+������Q2��h�T����-슊
)�Qq9�f���D��Z
|��엲���x�"ߚ�6S��+��0��ʓ����
��Ne/}��,Gj�K%e�Pi+YY���d��[�k/��O�[�&�?��i�YҤx���AjV@���E�	�����Ī��xt�,�q��m��.�O���#v~�]��\������"ϋo� ���k=iR�y���pl�ĭ^c!q񪬳\x��Gp��-�=u�\5��ڼ\�f.}+��G��ʧ�D2�����qP'�ڔMf���Q�޿�������k�h,#��lyu����'
jV�B���f�Dm�
�*�*5x��۝;�C<HR���x���>�+*y�0/M�p+�Q&L�~���z�7�����������i�����З�_�yw���OR��t��J����	]���i�&s���?�Ŏ]����.�	�o�g4Ɍ�����N"u���ͳ�29N>^'�Ð�n�ט�	{�)�SD��,K.���hЉ�GڧE������\��r�*y�t��C�lx����zr���U��_����bw��������ըoG���j҇5�:
L�fJ�uϊ�.֔욖x�w�;+��%g�����$q�8.�`����� �^�����>�H�?u��`���h�L.�d�G�,9�}�~[� �[�+��|)�Ňg8.sn�kQ�	����c�,?�L0W�Z�Q��H�5�G���S���G�C�Tyz�enϧ�u_��re.��}-Wb�3� 6B��c��#���� ���|~]����͛�m�۩.Jj庀�>��x�e�g��g�>����Ƃ�"Q�Z��y�PE����5m�u߄�2��M��'�}u<��e�ݞ7�Q׍�f('�'a���޺?I� ��e�
�;%ҽ�R�ް�j0�@U�+jo�BwL�
k�-�&��6�\�[,� U��{�;��o�/߇/>yp6�w����S}���خރ��[�Z�݈Ƹ9g>�eHY�-�=�7�)]�l�&�.!�4ɴ�^d[�G�u!��Ab�����Ʉy���nPS��/��c-9͍����^��kRO-�:��7ߦ�,�YE-�Ӗ�X�%u��������v�c;�)1�'n^!�ȅd��wǥB�\&l���Ucۥ+c&��B�t[���fz�-�v�ޟ1S<�X��M�t�EA�čt8Ӏ,sj&�.*�!��G{r%%���RuA-�QXPc���A?���N@���޷e�?I'�2.�>+Y��w�I=deI�ħd��)E{��Wf=p�y�����1Z���s�Q����i��@7M2덟S�ݒ�)�����~���Rj)AQs�NC�Ӷux}B�u��+�r�q��W��%� 3�ާ��{1Q�g�1�l6���S8����//6��@�s"*�(��n@�@����-$����N��E���1�y���5u>��:ٟ�6	�U����z��l��0�E>�=6~!+}��NtJ�ZJ&�V4�}ˊߞ��S�>M��i�3i�6�(�v:�0�9J����l�I	�)Q,�PH;eRBe��5�3�;�凊�����c�m._�����������4H���tެ����.�J��,b+{�Ԣm1i;2iB[��5��|��F�m?X�%�+Y��D���C��n�V��qn�kH�:�ݴg��191X&1�d
ŤDm��0j��ʠ�\��;$�%���)�Ei=��-��ص�m-So� �~�~�o9k�Hb� j
���]`B�=7[�V�&�3�a�����K|�V�uu�E&W������S����cS�<�<M�A��x�s"ur�i�R�PgŪ{К�pQ���-���a�1e5sC-Q�K� ���G���X��u�3>�p�I*�Fg2=F(]���Bھ��q��9�X?�q��ǿ(�2�ę3�r���&��6��p��v^��a!����g�'W��z��y�by]��nb�+��QK�aHJX�6�)��Vб�(�3T(G5�Pt�>*_�f�!%<v���|
���H%n�wy��3��U04�,����@�P]�}��r*T��v�����{f.E9�+s�����'d�h�)~i*���!�,�Y����c�E1GB�>�A1���o�I�5v�g�G<J�;��εC�a�7e��+����'��v����z��z�\�3?�볗�v�ڿ�oV7c��d�iQ,\݀%��>���F�����Z�$<��c�nJ���Y %\�qڍ���B)�1�ʎQ�u��j���D��:(�O��>*x�#%�¦s�꒝�QM�n`�.�I�Y�gy^��(=�Ţ�ms+�$�`�#W�}ZpB�ԄG%�"9�Js�b�m�9�{ ݞvz�����l�̇[@��:�J'��}�>l_f���y0]�����g�#�j�������}�%NJm39���#�;]].�J��
Y&d�RNӒ�"�>���:�"]���u��ļ4ꉹ����&�8�����G������,`Io����QP[�#�r�r�X�R�'���%�T��)����v��Q�񑐷�aK1���n���&�]"�
��הG҈������V�����T*q���^�Q��I��QJ�+��XN���]]Wp���a����K�Z���vg�
�K�G�5`��1oDĝ���!�~���Z9I��W�"�v݅���V�{-f�|bi�c���� �����x!}�֕ +p�x���mu.�B�&[�Vѡ�
"��̶(
5Ri����V�?���_���~�fu��x��������i87�α��h���з_ie�����s��\wXz�Ķ-W�J��Q�y����}_C�y���Z��H�8Y�6�f&���˙���da�
��s���2��S�`\�I�=��$I(��B밂U���A����3�jId��6R��>hֶ�֔`{��-� �h%��Q��'� G�"\7��)5��M:�!>J L?ÉA�|n�h�.4S�̃!���p��JmH�dT�8�90� �E�V#��ą�(���yAU�7:��I�[ɂ7 ��r�Q+>��Xm�!!��,�_�� ���[�}�C~�k�:K�s�5���CĞ
Ʉ�.M��H���Z�Ie$�[P���;,��T �"�6�&��(k�Qޝ1������:���*���6},�I��c
��\s�#n�[�V����8<>��%	�����/kr��PłyX!��ap����T� �d��|t졛�+VVc'�[�S�MFXZ���m�n�n�C&W�ǳ=/,*����#q��{���D��2U� �*�p�o����HZ��N'y:�U��$�����bQ侢����q㙏w�;/�N�y�g���B��l�8�<j���f�]�݄����n��m[zP�}��2�\����s�JY!�,�HDDL�5�
�1JIb�D_�<��� �)�A0��/�!���*����9���֚�K���k����?�Z{�S�����s����/�����F��V��t��ˋ"�A#�"���鑹,��`�̈́�[���5��������B��x�_�z�Ν���|�	�l��([�"��mܒ�5g&��1�f�S&a����_RQ�<�����l5O��؟;�vW~߇�٣�n�;�)�+� F��^`��T�h�=��Z�&Ώ_M��^�����_Rз8t�G҆*�mc$����&4/����^�eD@�h����.jW����%�	�� �ѺJ"Zsƹ�o��]�4�De��V:݀�-�?Gk�"T����6y͗�`���Gl([���\��*�B����=�����~���:~�P�=��FӨ���V�W�B���ԁCa$e%�aj'XU	��U14D1���7�o�p/���#�%l��Go^��ڝ���F�H��Q���t�TP�O�F��/�"���t���h���F#�J�� ���Wo�p�Z�23ʴ�O���s_U��P,l�$Z=��}�WD�u-���Gn�Mw2��yvs>�mn�"�}���_�_=d7�]�WFțu����ϑ?�^5�d��0_�ޡ�es��)j�3ݨ�>(��K#ǳd�D�3`m>��)$�HT�V��ΒH�-��^�"��~|������������*�]�o�B������]�@�?|�����_���ﱰ4W�� jq׼(N�E�Y���̳*`���*��m1��*:T�
dw��gIQ@����ș�ur��.�"�TK�L�g�^+Y���S�Yy�r��	�!73P��q�o�[�MY�,��N�^�*�8�ŭ�v,@X�c��>�5QAU#�U���Z��ރ���š	j�Q��
�&�tcg�:Z?8j?ۚ�O���M\P���M(4�� )>X�:R�*�ܽ�F_�����c�vV�MiOh���J�v2��q̨���#�246��L&P�����6�$B��a�9�vC��4,e����=[Ӯ�B������|��{on �J����\�2�^�h:�C���Y�綞'+"�����b=9� S�^m!8�,=��� ��ת}Đ5_1�V���L����v���LD��se����^Id��^8�Љ�\��ֺ�y�M�����tu*T�iȑ뱚�x{~�PFQ������Ⱦr�e���ʔy�/
����u��{a�D�ߊ�����f����ve�޾���\<�(G �޾�<�b8==�W/��U�z�F�W���x�z�5-���ES��!��m��|,Z�{�ϛ�����&��!J]e�+y�׈�hx�]��8w��c���
%�\�c��5��]Y���P�����iz5��O_�~�W�?����{���o��SW�K�������/��ߙ/����R���3�7�ޔ 9Zz��zG�ඉ}���?��-�[�p�G�Q�w�& Q��<Y��Xt`F7��z���b (�ZS�@3��j�m�>�/4����ۧ����ůy���A��O���=R��ٵ: ������(.2h[tC���{�gI��X����R�#O���v���?:�.�7:�:��G6zv���E����X��5mg�k�>SV8f��E�=h`x�y�2�	t����vʙldΓd?�#"���z?^�6�Q�эk?&��@�E���Mݷ���;0��~�*�J�%��T���'%
�R�m䳃��d��1M�y:t����~�Zm����O.ج���ѱ�3n�B��k���	UrC}���=J�1�}[E�-���{I�Î�	E���E�V���uAWCx�b��(�o�J���ûw����������׋vYC�1z:�z������|��ƛ���z�����M��n��V����qQ��
;��#X��6��:I�y��B�-K�o1���嫿�k�����߿���@8�SU��E�b��:������r}�̝[��܅�k�}1���ҼUe�F��& �WK��׷�z�2�|�/�����;�ë�)��ټR��x���k��My�R�!6����#ú)Ѫ
~�ho�G�A(�zz�t���$��˸�!� ��Hκ�RC�4ԑ��}Ԯ^��T^�jJ��Ew�w��+(K��kZ��L��*��պ��7�$����@���?l���[��\�^�� �Δ��Z��j�g��^"6}� %��QI��45��}?0���:�1��-�y��d����q�۵�\	���Oϕ��zG��j���uI���^ڌ��Τ���e���A��OƓ�C���Y]u�S;oto*��B��ί1XJg�d���ߎ�����Ɔ�����i�G�KΝ<�11����=r����X3x��:}�x6���u���o�%����(E��(��PN{���=P3{ʾ��Fˣ����ʚF��3ӵx��� ����_��*E�5��,��g��=�*���֢%_�O�����q'��uq���ֶ�A�Q��[�I#�̅F�*̋7p6���	F�$�D&�5���0��y���X���oǽ��:e���)���տ�L�j�>�3؞�����|���eQ�y2��W�����j�ӲP� Ǣ�K�	ia �RʂF��p|�J��3��<�R��Y?_d�슥��D�e�a�bļ��{jA�\7w0���k����s� &�Q��~-�I�C/j�x�E�>�P61�i(q�ﾐ�fDn�^B���E=Kg8�|%�v,�j���^z4�'U {�+����^��N���r?v�|��~�c���"��"�n��]{�k`��!wc/ÞܱEj��[�������g�/�t_�6a'Y1�1����ӱr%ͼ|����qS�^(f/c��hG��U��y�ݼ��a�n��h7��^��n�
��
�j�f�k0"+g�5���xM�%R����y�0��>����_��b�X���k�n��m���x�9�˽��qel�M���wX5Nξ��zd1��q@eBGE�j�B�\ �
��G��OS��4�e-fI�ā������2���y^}V���<͗`,�Z�ʆC��՚^}�u�v�.ݙ�]4��V�	���Q��6��'��%�%�������Dr0�-���4R�`�"���i�?��|��v�ǿ:��/M�~ ��?�S�����~��o�ݛo��e�������4=�}{��������
|[<0�B/
	 ��V�3������;�t�,�l�╏P臷���J�{�M&0���T�%��f���z��az��ɽn�����k-�^��I��[m�m)�ħ{J���f*J��(�L+zW��(�=x����Rf�UE���Q�'Q5 ���Q�6dw��
��>�x�;�A+�cإ���i��S~3�)�~/�#�������/��]���~���gi�`�z��+:5�)���Nb)~�F��cW� j��L��W�Z�0/s*F�j�0Pj�g�yP��y�A�j��`Е���,=�hu���nê��"�� �vh��>B�6{ġ�S�3�Ҷ��e#�:e�yVj���{�V�+�^���7A�o q��v	~B��7���=��Y��s�[���o5r��������xi߱ȴ"�v�����	��ݴ�`0�e�"'�p'<z��PB��2���^�O4���^��q�R�2���Mꮽz?Rׁx�[|�0Ѯ��~o��Z��Z�k_�� F���ϕ���VV
�WC�H�ޟ��Y��,w�X���\�����g����*O����$���)�߲B�^I�w����[����z�3����M�'�Xh/j��f����K8�}1��̛��
��-���H,�76Ў�$j�w�P{�H(�I&� >A��La�ڊ NrJWq"�`�#��/lG��!�������Cs���@�4�@M��|����=��y-�i�g"V�adi8�!4�he����r�����ʹ��Q��=�VkQ�4tƇ�ܳ�uɳ[�7��B�aý�x���Xv�~��[�@���g���ES����]�Mi{��+J' ��\C;�"?�Ctk*�=v�K��f5C~���Q���� |ٓ���5̹a7�Pn@v5�Xg���nAp���:�BGs�?�?�7�ɦ���9�sW��Z6�@:�ixI�ui�yr
Xc�����f87�҇��{x)�ѯ���|��k�z�O�Vv��9[�IG�t1DNU��6�M�GMљѢz(2�un��
�<��1�9�n�F��D%4�gww�{x[��I�����E uw,��`�P��\���R#>Fm,_Zu.rۿ�&�.�w�g~{T��H�&�� _t�m�~��"�%s���v,��]xv�b�5���Z���1�xw�����O����q! �G�|??7]/��\O�X���S`]K�g�kW�jW0�Ek�/��nu���H���T��$��g�B5����T�Ҹ3��Q�	�T���������<�Ӣ��y~g�3ⓖ��v>[*���z2��������NĚ�d��$:AMyy�>����R���R<yx�0��ё�Ex�(o�����X�v(w��G�n���RPϳ���Pc3�|�I\Y�:��g�/��7��nKy��%X��^������s�G6��yR�O�d�˂9t
_�9l�:hy������G{���<�*Dd��Wu��B��(�#�����1#/��KJ��G���*�j@p�Gq=�߶���#�#`��5�[����a����s���oU�Zֆ'W�5����
��@@%�=��iP��h���j���c���/4��X�j�����`�o7"��]�d#01�یZ_OU��� W�E�2�a���rc�^�v߮��#Ǒ���Ԩ]�GN��=����C��g���쳢�Sq¦yV�6@��"��tY�S�-�E�i�(ݛuy��y�u�Y�i�.ku�;��~zA��I-��m�]N5VMRq�6�5+;L�$�x�&�^�s߃Y�����'q\�w��������X�~���:b�����y�\�����?��O������I����r:���;����#C����^��MTDs�)�	�dJ3��-d8x��=��j�pn�gXwP�×�f6Ҳ-�lԖ���#��T@�D�d�T�gm"ϜJ�'��`�	�fq�`�nf�*���)ن�Z���� e*�)�{eIT`h}KWB7���F*��~���BN���I%E�3D���d�|����x]��ˇ��	H������Ť%q���<?E�7a�	��|k������)Ȗ>YjL8w4��l�o`��톻=|�ݩ�`4��|��m5���E��"����Ma^�߆��/4��;��e��t�Eq�ky|(c��F9[s�`����]5>_>��z�^o�|0!��V#�ټ�Z�`LF�\���EԨSwpz4WN����)�1_>���hl�s���ma�c�{�{d� *n���Y8��M1��"�d�31(����JȪ�*��.���OU���;Ԩ@Ȟ&0C�*1�qI�A�
	�X���F&���솲�_�4"G��Vͨ�=���@)�� _PE�.w���Z`��*��R<GI��eY^e��N��mr�|�^I>��V��:O]e������`_�����(6��~N�?��iT܉�0�
��� h�<��z�� QE&�=�!4�����f��ʎ�q�ȏ7�b��s���c<���K��-ʗ���)|{v*<������/?���u>������
}z���;����g�z��G���o\Ϗo��(�f�o�n_k�9�hiUT6=��u���
�M��Wa?�Cnop�Ml�:H]h�V9L�ʏ����?d�S��u��z����_/f�����)s��7��s�}�5LIDds���z󰗻�^r*�bi�y'sQ;����bя� ��:��z)C?�����ߒ���2�{��N�~$�r��nA��z%�����`JX|C�}��C��2�O���>&N���ۼ��|;ߟ>��
P������15t{��RE�&,��8"�l; �]����A��J��& ���=�Z��Z��i�Li�̅�_�?u?�z���ކ�o���Wf��n�m���TC�7�^�lS�Z�f�3Y�,��x�����$���uj���4�^/�k�j��ag�[�}��-�S���%r[bթ�hN�hk>�����f��;^A�������ϋGC�`pg$�	�H��?ʬ���P�����,?S��Md��{�Ҍ���2X��>���]�~�x޻E%t����>��e�fP����nJ�fpVo�0�Cu�܈P%O�!V:�i�#,��e�L�^�-��r�4���\�J���Ff���^.���5�a�%8���5�c)�U���$��_����Z�5�x1"��?�B�ݡ�҃���?���;����r� �j�-$kɎ\�ε,�D3��ܳ���nl�G~�؀3n�s(�k�z�5�����TA���~'�~_��P�����pS̛UG����������<�I`����ьr���-
���܅;PHI�g2����/�,S���{Z~$OO�,ro������^����=�q�N��p���b	k�k�8��7�v�K�*�AC~�4k��7k�!���y��>�����><�~�.��?d��z����ƶ�])�qP�3��M����Q�e0J�P ��΢��40��B�^��؟�[�}��
�l[�7j�'�b3g�!�[�L�<�Q����sg^����W-��Fz2�ޑ5���t�Y%S�p��Y�_7&��6����S7c���Zq%�G�|��1���H��ӏZ����^q��P�5�^�s������
!��x|(:�c����6�"J���W��g�q���g�(F�8��*熕k�
7�mܶw/�6�V�����T��!�������Hw,���
��(�=�[�*�\��4�F1Dfᑣ�eV��:?	*���, F(Y*����=���m6�=�q]��7�s�+{���F�����������G�����_����)�����Nq9?�����/ͧw��KٜW�6S�vX�Y4������>�j1�:Յ���E����6��=��� Z�����ꅺ��+h*��}��·�|��m�^ͯ�3a��Ԭ��1��6
�C�Xl���CQ��������l�}��+
�5=x��\e�'�J 2������[?/_����Y�Կ
�i<�c��S�X�.wd�4:)�0ރn�$�_��M�JáG���`	U��Xނ�^�O��S�Q��>Hj��X�K�ȣ�N]���y~92u��2L4wYv X����xO��ˇ��-�ZL��mpٓU����|�$��.���YM�er;�������]�|��#kh�b4V.��0���Մv�HYt$;�C�0�R"���HY�R�Q2��o���j�U�����ߩg��ٔ��P�^���{��cp����������K������ah�`�'�����Q��=Gy�;$�eg{���9��k�*��2CM���LK����(鬕;���U���m��aE�`.<�a%�����y�-oU����wP��+%�}i���9�7�w"���R'X��*�H�~�>�ax*â\��s�5��<rR�l�)֋���*����=%d�_�9W���(u��)ʟ\b��������w��<=�H��>������|щ<�-�g�\��t~���ǯ�Z�;ԙG(oҼNT��$��y���@��h�Xzu�&��d�.���`qԉwf��
�#ʮ����X�Y�fx��͡},gۉ�vM�b��ڭ��N��=���P�*�VEUlQU�vo�8��v��+�Rm#	l���������}W޾�L��b�;��>�I{G>V|*w��vh�`���R꽭/�=5T�B��z�~
�U�] �����龻v�����dyҒ+��C�Fs��:ۅE�wr�������E��'�;$,YS�g,�R��j���|�|������V5�7��C�*�|M�#Z*�yD��Հ�T�h��: #jpr�s�AHF�*�g�v<gO�ʛ��(�\��p%V.���#'�	��l��>k�q{�.��t<�9�܍C�>o����о({�ES�~���VC�5�Η�pxQ��f �^�7<Lf=Ǯ��p�� ����1����%ˈ�'��G�����zQ��R����ƽېf�9�_�7�S�l���`�AI�X�m�0KG뫆�6�BE։�@C��x�a���gȸ�V��HAʈzP�VR ��4F��K�� ��V�l���;��7�7=�wG@�4�A�p;�FS�
^oE�;{�a�p�2�)#�o����o��O���	w��Ǐ�����&-���r�����_�>�V�� �?+9�D�����Dn���P�ތ�J�<���}���B Q�1z�C�/�v���LD���D]FCZz82y��L�%k���Ѽ��� �k��A�u��9�F�l�+�2?r0[,g����Q�~�/9\�P4j���g����O�$���坻�����x�����>�s��r?����!f��A7��;=f��թ�r����7o���<�	�m��	�7E���j!���N�UE�^0�=�]�0ʎ�xWzp Ѷ�ݩf�+Bc�.mL1Ez�#̡յ�xnU�o�Tz�ln�^��z����.u��v��Ô�y*�w3�=��5u#�͇�0��a�����	r��X�EP�7��4�S9�U;�dݧ,�,��n�WȵwOE�T�\2Дzĝ� w��_B���+bvy�/מ�����i_�V3���9�lQ�\�/n4@bM�Ziٮ(���ӎ���l錸�ދT����C���~�B^�AK�H�؁�x��P������^���A�]O͢�9T�0We��h�H&�<�8�X޳ WCJ��u�_���P�@|_�eO<�G��X�Gp��j�]�G:�����`�y�������ȝ����.���9m��8�}nʹ����z�f*/��#e#�rT�	;��_ᡫ�D�M��~���B8��?��5���p�V~��)�ӻwEYܕ�9a�~�x�n>��篧ޯ��妴-��֯�Sd
�kiU.w�PK	�]�}�]>-�p��<DW�����db�&�ڒlK�hf���D7�O��?ف<ǟ{a�B�.�*,�1��|�<�gR<��X�Dw��jݦ�=��r�E�#<�{���@A���x�&:��C��x�k���*7���{E�iX��Q��r���G������o�#�h���hlT�-U��{� �(z�\eq�H���k>f��?��j��"���c2(N�/g�3�!0�נ[���Ƶ�&wE���p����r��������{ �s^�<g0�0�*;<�1Ve&R+7N�KG��{v��`�Y�֥�^e~����������U��e��W�a���$��^Z-�9b�A���Ú��geAiL�����4Sb6�we�3���_k�;���-�$����]�:�òq�ۯ��$���o=��R�7n<6�C�>v�-O��i�{ Os80����{��Ľ����@�j`��dW���[��As��_?��.���H�w�a�^&�,*Ӯw\ټJǭ君���)w��w�am4bi^jmuٺR�g B�)�"�"���T�����i�/:	e|�����gU=aE���}n�Ý�C�Y�tb�<��JW+m�]n�՛��c�������NW�@�fݪ�oķPw�m�9���YC��Ɯ���ǿY�\R�U���M��U�yz�R!�����ݟ-��_ZO?z��w��IO��fKN�=g״�rP�"���:�ⱆ�����Oͳ��F5�-�����&ر i"�K,���w(�Sq�)p@�;/�G>yY�������Z$uY�b��R�ŰZ��޳�n#X����+��:e�/��-���� ��+�,�c�w�5� ������;I�b�.Y���o�)�2V@ǿ>|F �~X���/ ������읟�����E�5M�	(-xS(dHKk2	X���ee)HP��i��])\���e�]O��VHF	�\P<g����Y]i���n���;֍=�t
Z�X�������#�	���W>E�G�W���2GE��/�\�2v��/㶔�>�c�OlMH�J�-Azu�l�1�F����k�^��pC��4T�J�[.��c[�c�ߣ�j�@���(�в<�j6��!W�&�����|�����W��zY�F�ʚ�F/(u��G%A}��%��ٲ��T��X�W�n3fl�A��V~]��|��\�@{�ym���|��:�v�U�r@�#��6�
v��16 ��<0������y��)G�o^_g|M8���{��@�T����^�N�^�Q2��j7ID4g���I�5�e�6�>I.���0%a�:�M�Ր���~��� �	Q�M<��!x� ���h��u��Ɖ0���i�(�U��p�J�|(J�]��ׁ�]�L]6�Dyٵ�����~��]����`z�S\�=1""�bK��QvEE��%��x�����ͯ�ӣ\���oV�6~U��y�����|�{���ry�3���'�R//`S���^�{vK����ۉ�{ܿo�Ym��|r��������jZ����P&XЁ�D��}C�Z���NoF$ӟ�<��Iw
��T��c��^�]�+s���p�Y�~����s|�#k�A0��I.E8^�<w0�t(J�(��0f��JA���;�k�KV����Px ��(��;ʮ���Kf�����|b��N�/j���roZa^�-�"5���^�OE�(X����dG:K'�(��pZ����֮��Ɯ&��|�B�y_ky�%�s�j��5����H�I�}(61\\���f��24l�7��ml�T0�_��-���kϏ�U<{O���e(�����]_B�����uL
����|�`�+���t�j���G2��	 �aQ� �0�M�#��%��������k�F3��/�H�zu���^��"��ЯG���G����J��(wϻQn�ѽ�u�������)�8����׮u�5��Th,|�M���1�t���`�Q�A��}���!��8���@�3��G���U#�u��
9U�ƣC)/u洚A� e�����@6;(sz�@�f���Q�2	�@RW�h༃�;�sU�����Λr8�Jl��/�?|G�&��J��n�����t�Gv�a�l,}9�3�Ǘ�vr���_�������7���w�vΉ4x���Q�$��տ"ǻ����r�!����|_~�w��w.~����ß��>|��H!�S����	�k�CPC�#7�e5A�7�k�xc�Nw�=��Y�l�ia}Iئvj������
EA{�@]<��K��Of��~���7 �&W�F�ҶP*6��9�����@��(�����;��ϏT�;@��%ɑ)t�Y�XD=����xG3�3�b/J=�1@ɸ��(�VTeƼ(<*�1� c[��B[�d\�
�t|Ey��cic��@�b,(*�8�T�V�<u��aC��������_�9���>m���B��(%�2(�����#�zܰ��Oh�{�k��cUVַhƗP�[��i�/��}����6�'%sx�QwH��[�u����)����Yk����W��ο�_-�bD�ƙ�%�g�_����&D�D�*��9�S��g�0�������K����_���E�0ʳ�~��fS��*W���u-�Bv�o��90!�y�V�}�����'�TY𖵁e@9	0HW#z��ޒ�#Q��ma���f^�T:Aw����Av��F9 'Hڲu@�JC�Q��L�x��]��'���e��7 ���\�SJj5��jm� Wp��,�Ψ���#��b�5
#��li� ���Q��'��7�]���d��e�$��r��xqGE���t��G����FU�Jy���LGd��pE|���~��?���ez�O����cw~�������3ǻ?F�������o,O��}�ˤ?	�������������K�:��ѿ6_>��r�����,��2��B�����(��#C�z�B����.d]�>_��Fl�΅�Y{o�;(�����`ĬV��֖�6��j�Y�͆ͧr��V_7��jt��w>z�t�|�m���P`�V����0T�r�e<�1���/x�j��ɱh���:'-J��<� ژef�|����>�G���ͥ��Aٟ��6Z��A��$�X7�_S�p�V���"S4���깣.tz����<&�����N�p`e�)��z[�|���{p6���<�����Buؙ2���T�����QO>�,h���&"��'2���	ePF5����gZ	Q 8�y�T�=���k	�	����h��B����~�`+�%i����L�ԑ�Ӵ���v����a������������o%|�=	o��^Fxxz�AF8�i�ծ'{�ޒ�S�6ɪrO��&�<qk8�X5�4w��֛����;�:��:��g�M��L
r+z*`o��ͤ����7I�v�ow����Jf�s���� #��a���SLf+�|!4�R�mQ{��U��){РZ}��*�C�s���a	�N��\k�=��(�E#?��rw�A��� 5�+Y�"�(-�bmR���̓M�{�<��k包�s����z���ȍ�����W� 	�X�n����7����������o��Q��Kx���3?.�w��zz��/������E����1�zJ���^}�����b��_^�_�L�~(i�uU�����)�\�0{2�sS�J��)i�o0�S��k������^�M�3f��2��,����]��Y��j�XRi��f�<�`���E�F�Y� f�H٨�q�� w���$��@�X�z���+n(�u_'%��%B�k���|*��*��H�v �����S`�:h-��� �b�6!p�،7D�`D'�i�]���N8�����N;�&'J�"㜨�I�h�6ʺ�TA�%�".4G�ܽ�����}U'O��(�$w���RKn�S̐c.�6Y`?tr� S�y�>�^�b&�x�	��\��\A\���U//(�M�?�� ����s���&�B���f����^W�c7��-a#�
�V�x�5����=H�'�2k�hDyІ�@�Q����[�3��B��p����hshƇ�_h��o�����'?2p>n�N�j��ޠ�#Z���j��dЎ�����o��d�\���2C�l�F��|]ƭ(��q�^aZ�*�s�>C�"�F1��tb4c5cdD
o��l����rN:��#Д����0p�*���)s���aΡ�9��K�b.z���i6�mvc�@p�ph0�|
�Z���&�e�@���J6��=�]��3���1���^��P�U�yv^<R�Z���h5��q �^�kz�'ְ~+��������Ç�����c<��7��.�Yb��e��\߭���^NOO�qH��,oW,��D��JT�U�B�8W��JD�є�hyg�vӺI\��B��J�6*xcguk�d��,��J�7҉꥛'�JK���o+ָ���Nݕ�e�m�l9x&��WE�vޠ�������M��P��=��_�sQ������l �@iڒ�J7�/. ���w)��t9��z�R'q"�@��:� �̆���\b���0��m*�QK��8�k�`"ܰ�$��? ��aEe_5E�C�჆�%���1�"F*C��{܊?C���B/F�Ս��q��s�xkY�D��╧����6H�A~��4[F�?�x� d��HE����?x��y{y�yA���h��Z�����~�=�E�Z�pg�D~D	>�8�}��lmO3�(����%�:G:f�Ww���YY9�G��Ywo��.�E2�K�����@pl�a���<e��Sj���؅��O��kn��κ�9���E��^�6����zѡ���F�2(��30

JvFU�Y�~��B���ܠ���d8�S����Ho����B������T��a�g��7��N���̢eFW�!�2�.��"Vn��R#�ڼ�;M�e��˼�^��3�k;���׌��Z횃��#�H
j�qR?�K��̈]��p��;�u�#N�Aκ*jȽ�_nijX���^�Œ粀�?����,�{w|�_��W��K����o�P&�nW��8�e~?~��0�{w�æ���7��&Xsò��Ր�W�#N�-�.�Ym��o<��+��m���t��z���!��O�X��W�UB������h���ϩ���\-��_b2/]|��í-C�n,����W��w����W�v���P��sD��&4v.4�������X�����^	9��bw��?��r+���A�T����k�"(�E�� �a���F
���cK7A�\ط��G�M�;�"���t���ר��qo���I-x�\L��@���潺���^Wh��@ܫ<u��Aq�,�X��t���Y��}Piy��x����.�]�y��6'����R �W���B�\^𸫡ZݠfH޶��7I�t���<l�zC!7Ӭy�����ׄr6�Bx��i��Iz0����#a�;3������*���*=i5�Cv���bƚg��0���;2�4(�f�u��s�Tai{С�U�(��@Xwz�96�	��p��C�l�.K8�f`k��/�_�����W��ْ�)�x'/����t���8 pV�夥���;**�ʜ�0n�FUi��}4åS U�6��
�ZD���ٕWVO��1j8z�^8�/h����ɼ��O�欶�:����c$�Jb=�����!zS�t�I�l{�y�?���� �G.�a;r�����$A<�n�C3��N�ةde��:�Hw��`�����ͿYd�����ey�_N��<}�5ٽjy�1_�O% ����b�}��_�����|�����vd�P���G��X��f��h8!�����n�m�	d�w�j�I�-#nl�B	.�sd^kf�C�D#!w�aRe�,�b�b�?�!9�a��1�6���S+��.=�nl�f�TO��C��+0I�
�<�FI�h�K}��+�B8�X��R,עG�j��J�p���V��{� ����?�.��yf��$�)�;B�#����
*ǫ�㡚���k��-q����͑-Z���"wAv�9�l�Rjq�j8 �ʜ�*^ h��fDqj�ddC�M�	��?���LP�n���Z��	x�����4���TҰ�z�D�fF��e"o��!��}�E��[w#�H&���uvZ�;���u���˕D��A�{9̛r�q|�y�;�W�7�y7q�[p��1�
�P�F}��0��憊ԥ�	���TƦ(��Pq w��5]N���Za�@����'�>�8��K	�*>�*������%kŬC��
a{&70k�q���p��,-]�m]��*���G��"Ζz0#2�yp����� *P���}"�YPB�n5��3����Q)�I;�r���)΋�����2��X�h��j�RW`[�F]Ng�=�d\��Ԩ�<:\�i4��H�Ȍ�[��`qs��	�R�m����
 ��e��F���e�,C����m|e!������fBS�`|d)�j�;k�8$u�$
��R��k��7D[&Ϟ?�LsFkHD}5:�&1�3k�K 8���g��g�����H���S3��,�拲��鼻�}�l�m����U���!��_�K�]���˸N_r�W���EeMO����d���伝γ.w�hO�pe5p�{_m+�{g��C]���6�79��Mx�ˬ��[�+��5�g�{)*1��P�@ќ�#3�.e�3��Z�֬��^T���{C���vv�\=�g�K*|�N�{-��Z�
�s�k����X^/
�28.x��lp���9��a�����bq�z�j��5�I��Z(ڽ�Uw��V9�:Ҕ��\���R58"m\k^��`�	���x�a��1Rټ�D���H ��頣���'��t��{x�QK���+S�k��=�1D���ܤo�4u�0�,{;�A�s(FJ�*�3Il�{�U�^����ж�K��c�O����F�˖��"K~�~m��:=�J����X`�i�d�� ���׳�X8Y-�X#.`B�関p���	4��K�?烬��A��3dނLF��-�P�O�u�s�;���-�"-7C񩣗o�xĔY_� �{n7/^���\���/��K��R��` d%�B�G3�c7��Xj EO���Z�b@�y1,&x�Eֳ��jT�Ҝ��2'�E��4ן�>�zյk[݇Nڢ���,��f�mx���|J+2Lm�G���cr��1jU���eF�y^x�+��"����l����]��~_�5�-%%'̘��J~�٢7�����ڵ�8}�ݘ���/��B��e�v�_,��/��t<��Ӕ����G�Я7�����ӍW�勁 ��b��Y���CUw�A�
]������f�5G�7���T!�usl�)s������7���H��,�����묗����Vt��x� >v�F��v���ϴ��ȊBNū�3s�$��!�0�arS!�[6-�o*�3-t|�aa���f�żj�!0co���	I9�~�Z�fz>l�������
�-{�o���]�E���@V�VU�/��5�l�R�.���8E�ࡺ��z�NAE�ymC������i�2Ӓ>�LG[��:��M,I��iTH4� C	��\�j��<�:c!�����n'��I��GcV���TI��](�5�T�F��-W�^T�P�R\�@�X��M0xN5��k�^)l�R�"�;�S�t� ����+J����e\��I+�ɈA�]�^ۚ/E�.\�2�|Y�I<<H��R����JP�"��t���/5�����9Ϲʯ�7M������;�=�a3HhU��0T�orHr��N�rrh�W�o�ߒ�z�����e��@��vy������Ϣ��e���AT�]Ǌ�մ)��ޒ�0e� O���҃��ү���j��L����X�f�Væ�5צ]eJ�� ����ݞ0B+`����l�25<?�F1U�N!�wa��c(�2n������*�o���&g�Ôٚcjs�Ϸꊬ�<d��p���Y�_��Af�0��N������(��?���!��5��z��@��}ݓ�_.�~x%��t���H�g�s�Y"�<#n�κj�\��j��Z}Zk�y���ÿ���s_�b����b�Hj����p:�a�[����b��l�+]�|7m�Iܣϝww n�$6���Þ1�.�_{\P]P炞j�,����}�
�j�-�= ���"~HT1cf&x�˩x�g�ۓ�,� ���_�lQ�FMT�(�������4Dsa�)�f�;f�R����U)ЋAsj����٪$�Z��Pj�ˌ9_5�5���U�5Pb�^����[�LYU���;�ژ�7ڔ�-3He((��S���|\��zb��z���j,rL��H�c�e�>�fr�{�.r��|I��5�5��r�H[�Y�����f��8��FSp����;����`G��QK�`
0m2g��!ܑ0FZ�;��OD$���`|���aZ=��dB�8�����Sj��������ӕ�2U��Y��ۜiV�R4�w�F;��hF��ٔ�a%˥v�\�eK �^KKP���)��A��r��(��#�qnTc
f�	���:q\w�}U(|�S�e^�G�
�_k��t~z���|v�]Ĕ[�*4��N��Q��$w���=4�&]5���'���9+(5ƀtƃ���(mV�/j��?Z�T����DC,Z«F�쾴[�r�h=�b���2��A�����^,ؼ<i��Ų{�|�?��b ������/RH������rxuW�O��p�6X���n0o&�J9h�`4��6ܢ�;�E�T����$7�i�z�b�s��C����d�~ּY�YoQ��;���� η ��>�ռ�zn���_��$�%�Nj�lY�`���(�q����ղ���ٰ6�8]�����_ɫ�D�k<���<�u=ɮ̻#�;�6�A]����q<)S�7�q��`�W{>�<�^_]�b���F��9.�[�S���kٻW)󟗵4���j�\�,�5���ê����Sÿxл�!Q����Q��a#v#W<��<��,ݲ�0�ؙ�z�ȓ"����F8*VܰA�f,K������ �^k�PG��j�V���Z��k�~�)��G�p��h���H/d�AO��ֻ@��Þ�º&����j�!_8	j(�t(+�)_��>�$���`�,{K��^�>-����y�����)�l�@�*n<t��k�p���w��\W4�{�;jgyoW��N��bH|��f�>(�J��#E(t'a-�{��x���c�̇2�����2�߳�C�=��_�8�\.EV\�ф(�x��[h#խ�>�A�s����^gk P��#Qcx,�O�14J��I�����:C�FK}�hA2'�S�T��,JlFͨ|�]���T�����/��Y������6*:fz��y���>�(�N����r�2;�7�C���d��Ǹ��dr��d:�dBn� ��-H?4>�
ָ�k�]�݄�{в�T,d�5�ja�P����^�:k�-�TE{��u5x{V�f�J����[E�pc@����/yX���zo!KO������wEi(���c�2(����/:_���e�����<�X>��7��}���?��˗r����H��x�[k/rL-��FmF�]x+3CX\��BL6�5��C0�}�J�j�n�[�U�Ì��E��\��z��/j�2�s�2!�˓�	6���  ��(�	�rMG��쵁�iJu� 2�({������LN�'|�!�J!�0k��܋��M]�zO���-B��^,���H*Ą���hB1�wW���~�t��=n'Dhj��H��ܯ�e�~P�c��!�ދ�P /�׈�l�j����TJ(�J�{Y���ԕ��h�l0�H	���F��8YjE�EANq^ߌ�'����?���d#Ϝ��	����u���[�n��O���uͲ���酘�x�^��T��h��S��H_15�ߧ��O_�r~'+�9�1��YRԸ�M�/�{+i�[���S�mܺ�Q���a��"Ug�v��ji����1K�{��C��T�u��'�*I;?�"�CB6��+t�1�^�@�0����Π�"�:�W*T\��%�2~Wˊ���S�6E�
�F3<E��e���;a2� �f����b�9M��ray*�x�{F��#�t�-�+��_2�u��W�fZ�8�?�2W��� �]U��Ԉ	��������A=�Z��r������O��lR���Dj�X��^6�q��u%�߫�s+�ţ��f����G#���_Ex�7�y�B�zF��F���l�f��`��V���
S�e|1��ꗴ�T�M^C.�@�`M��t�K:˵x�;z�څ	`%ҷ��l�_W�k`��0�+�D��Us5��ZUw���ɐ�bv��5̮�E�tRj3_I%\9�E�!+�y�Y�A�Ϻpԇ/:�Oҁd�m�'���%m0Z���9;Qs�S9�u���	�cC����|-�P���,ic�-#|�;`Q�����͍d�Q�5���D�N�g| �}���T�\�����%�^�E�o����S�A�US�̎a-�IM�hx���=�f
 9�.RG��|���LX��yR��e��	�Zd��9�e����<��K��)��,�B���d�Ժjz �fT����x��OGvΆ|s=Ίh
m>��I*7��܊���^$�B1��ӏ�B/��I��;&�~��>X�ԓ������si��s/��m�#�{UIg���4�<�5��q�5:��W��D7R�F�S��⍲D��B44+��:_�5������ƃ;�v�xR�ol|�ը��!�ֵ�K�(���U_��)�Ք���$�������1���[�q��:f��&^�o��e\���ڴ,6��Yǔ�K86d�7h^���YrUug��EZYWP+?c�&��'�jq���6�D-:��m���s��DVj'�mj�����m"�-M�D5�j��;@�7P}�O��n�v�7��(Fs�s�4q8�p�Ѯ��9��L��;pYhZy���4/^>�T�2��M�ZԣKy�۵Eu�1R�g֍5�Bnat��l�'"r�F����K��^�ΤOP�%=D���׉��m�l��mfX�sX6�Z��zs��9\�/��Bw4�S�s��Ra�Z�3���2(P�Q��շbp��]�EC�;4	v��Rk�1�E=v������H�k�>E=�$-�Y�Y�=t�Udu�ʗ:b;�ڣ��x�Rt9�Z����cɏ�� �O�殏�-{�@yG�R� �[�rH��2%b�kxD������qB|��U��%w{_�
�4:Ae�-:j�����U����0D�QC�.�U�j6Fd�ޡ�/�+%ș�[���H(Q?�T���1ƫM�c\�%=���jy�{� o�-G���ʉ��D������x���Te*t���*V���б��l��u�>��1����K�������+]ĕK���,5luJ]��T�k��D}3��1�!-4X�{�Zme�N����Q����~�y�P�����\qЛ:���a{S[�f�����)3x�9I�b�Cgr�#�pP��8	qG �A�%��dT3I1p	�v�Qe�=���bI�GQO&���^ƽ2�h��);Z�^��� �$����e�ު��o�+sg���i9fiHy�4�'�����Ud�1r�-�;��>�	�g��9�]k�]�)6O?�S f{�+�>�_8�4� B�)*�o͚'�.B��a�'�ZiT����kFY�P"�l^�������Z�w>�{h.�]_�sQR��v��M��`����s�G�~�U>6$�2GG-��$H*�n�O��j���rϹy��[d�om�U�W��e*[�4���#䦠0�Z�_�˜����h��O4�P�^���y���e�x���T�Us���g�u:X����n��u�y"������lF���ڢ3��{&U��KD�P���F�0��j�v��,�*�I������bYҵD�\�8��W� .����x�.2�B��K�'-=Pm~�+a�c���N�8nkIjtI�8��=��"iN��yP�i�����|4�1�M�w�W^���Tʀj\+��2��!<E�W��,�>(ۜ5�5��|��ӓuTZ�L�uVC� ��'�2!Xʴ�u}9��۷��o�][��H���t�xj�J�5�orP�����~H��y����������J[�	t���9�����T螇�]֠!��Lup�"��b���`����9K#4[�@*��`Z��Z�c��1���w�t�if�&.���ھ��4���	>[��֐OX�D9ٞh^�vÈx,.����-��{�m/��K(t ������ÑN!l'����$�K�e�����_oy�f����E���u�,�r�,�|fDdUJ&��&�8�Z~�� [nz� Թ�3�c_����{�ˇ���]�-o.��4!�~P�=�U�h�og�XH3%��Q��HqF����7c��{T:���һ7�a��а:Wm.�3�T<�� �������/J�м(��uR�
Q�{4����= �g��%3�@PT\�W��8�d��F�qԖ�=p��2��j=����d��+����[��{��ކYuL�+��
G-�A;߻�.ʚ�S�P�>� %H��A�������1��ԹGid@��9��-E�C��(��o��<�/y��(���Y+]X6������TCY��q�A2V��bڿ��]�j'5
��fP�Z{��[����Z��+����j���a��.ZX�5���an���z9�8�}�5���|p�b_��A}:�Gft�5�:Q['�)��c�Ot�MQ�x(t���5��3k�n�B�^�����4��7Mf��
dd̖re��3�U��;uF���S�7 u�4���wv jߝ=��u[7Ր��Em���X��j�:���L��i7��N�3xogL�*����, Ve�̄5U+�X>1��Ͳ	ղ�&p�y�=��ج�ؽ)�d�bo¯�-;#�sM����oW�z{!:)!wO����J�S
]ﱻyq#�3���o��S���N�u�j�QsE�����Dm4��|[���TVS�k]��pV0�\X���/ ��2�ҟ�����O�G.�����ox�����ɭ��Ɖy�®�\���B�h��y��Us��B�����љҎN"�=���l2�+�vQ�1޼��@���I�hHvd��a�SK��������nH�%;����Y�:�Y�ͨm��V�����O��u��$��/:T�\'/� pѽ��@Kւ�!^�!���ѭ��� �8_����MQiL-�I5��'�,'�����F#=&rVG���޲{��>zy[�3�O�p_{o����)�*�BS��2Ou��=�Z$�ys��>sтqT�cP�~9�.�������|6�G���{y����vd&�Z�tU�;�ᄓy�����F���(5���������{�7U9^���9>�h;R�J�D�����S�!v c����GH����W[��h���-f2�uh��K��/lݔǮ�a�����t��M��%*k�����X$:�,	Z~�����������4%��A��?qD�兼!�ߴ�+���ArM�6ewd�5o� @�e�?�k����u��n�u�&��1ED�mg����ք�ǎO��)���\��V�􎓆m��Z4����»�}�>[��� H��Fp��.Ys�:��	AX��H���9'5�ZAdN��p;���\}��u2��4�:�`�*`-nV�N�kf{�ME�k��ec���.�W-d�ls��>��\H�JO*4��Ž�' �,���;t�4(���,2b$E��dB�Ě��|ءMk��!�u-��Z�?|M4�����s�o�"*D� /C=깷X;���-KW�z����ޅ��bWe�J���3�m00	[U�.��+y���~u������b(ܽ"�BXic�F��O����@��1�8t/�M�on���C��\����h����ޜں�{��ޔ��1���UDIt���ǫ(��b�u���):�_/W9O�XT�|���������P@a���[��c����ɯS�ٍ��1k`����椦�����"�	���|�n�<p:��dS�jWx�7|q|t��'�<�փ�+MK��������p�%Ǫ�=�Ө�?&���tG.�9�b��:�t�rOM��T�����b�FPY��B��e�P�;�<����5��rR��$+uj)$�7�M���ɸ�T�5?%n��{����Yn��d�mYN���o�u-��,�q���@�k��I��j���b���d��5��i�
2 �Cq��`�,e�f#Fl��� Osy�Z�n"�.�թ������7�W��7를��`t���6���NĐ��Z�ǋ��S�P!^T@w�첵�$��)�K��t�vmv���s�C�u�:�ʎu�L�X��yV�e*m4�*����U��!�O�?�yN�7�ej�Lq��&��#����x��qhy�m(>Kjv��ﯼY�7k�ז�:N��9�u�Ϫ0�s�8��(%?�¨Mfg:5&�5�����؃g�Δ	�8h�U�+K����hS
��cq͐�0ߤ*nU�ye�BW���D�f.t웧�&�z�=B�wl�	��@������.܌�.�Շq��ȸQ��\�yY�3x��c�s��B�tr���i*��|�ӗ_J.?������#�]#{+^�ݣ*Tx��v5t�����<�͑�_|�Zt�sp�$�x�7o�U+���Q�s�fD��إ�q�'=�g�q�̽dN��E'����Lu�J��5��l��|Tm~�^$�q���t�ь��YBL��1A����o��.�r}z����s���ւzk��<n���1�������&T�Z[բ�������gC
�pb�u�s���iH��s�m�N�Я�Թ;���䣇O[�yօ���BK��?zv�hc��)[��>9�cQ�.U�^�'�f�u��:@P"o~�>3DO�T���� HaR��*>���A���Q��	���z��d�P�ZZ��^��H�bV O��k��S֒W�L��>6����`
ٵU�� �X�	.�k���T����D��@Y�H��s�S�gۯYs�@�/��uT��}�o�2[<��h��^�	��c+���E�!���-g��x���Bl{D^<����3H=O�)�A��).v&-c%���S���Y�8_AJ�P��!�>�.Zb
Q):��WOO��){K�V-QL.���SJݘl�����g.��q�ѧ�i��-#K���[:��L=E�e���v'P�Kf�K/Yˠ��9o�����F[��lNZƷNgF㰗�W��1D0�2�^)��O���"��x$�/OOdSŜX��л�]s��alo�^���؅~MuQ��}�f�\����a�x�4S�����Y�7j`[�����1���`kC/'��7'��B5���P��?��C����d\V��Z6-�#T%wZ���:��Е`6�ࣩ�c�ܢʧ	:(��$�|-F%B=g9��i��~�xSɄdp�!6!Ѽ�ҾT��/�`��!�=㩛�I^�Zۘޜ�n��p�M�&�:�F�J�dl �`�V�<yp�g��6��ã��}������n*�ȸ����V0e���	9��+����}�e_��+zI�*�Es��*�Ȗ�'6���NP��8/sA�q�.Ve���'礬M�se�^��jW/�}�.�a��:˪�W_T�F���.Q���5`sXC~m�5�csB�.G�i�K��tm-?W۰�jȬ�w���0`�T�sE) b ~�ݛ�L��6��!��fy��$)BXؕ�ꛒ�j��J5Y�k�)�X݆@�OlB�a}�ƨ��F�Q݆�v��s�Bq��wķ�r/�e�O|_NE��"�V��e4�����k���@���l\�B����YEpk>1�=g/uꗈ�닥�1�C�76��e~�QŮH��F��y����vņy-��r�F,(��XΤLV$�������|jb��"�o-���ZU�'��YB9����;�o�;��9?��L�H4��e�����\�����d�Ie=���yk��2jȇ����\/�H����q������j��>W�Q��J�}��j�;cb�r3���9�UYVI5:C��U��6�^��;��Jι!��Sg�(�Zw����ӥ?a��V���^�V�H�"�a�`����R�&\�ʈ�sq_�g�Q(��	�TF(t�8��Ud�z�]TZ�ƌd��x��F��M�ӻ��EK�Ue��=�mq���t�=����{��S��C�i����5Ёoܺk�h�Xd��8���">���٨�"c�˥�+j�͆A3�(�e�,eU�d5|��mDb�D6n��	�Us��J�C�0{NT	�1c`���A��=dޕ.�X�"��3u��Ϳ��0up+���i��l@6����k2wF*
,?J"���b���F{4쌶��ߕ�q�#��7
�f7{@�v���zdqnJ�[��������r�T_˭�OoU�**����`�&�TЈET���=m��5f�J���Ns�'�aqlJ�[��f4��k�zn}4��ހ7{��ą�&B�c���W%����hBY��A����^�t�̧"S�.�r(�X�A,DB�l�>ur�NV�J��RP��|.�j��"����͞�3�g��z!qr����k�����;��? �}��]��:�w�K����}���G����B�n4��W�i��ϛG5����S`&V��й��c��&��YGH��a3�ӎM�d3��V`�<�k+(�w���b6jZ�_HC��;zd�`�F������:�9��kx��e�\߈R�9�' �4x�B�5��ቻ��=Z�=9����s�����t���s�P}�ze�^�NG���~{�\���=�ݤy���_c�p$C��m������<��,r9'|R6$ ����n��d���m��R]-̥u�qc/������|�ڂ�\�y��m̭���Bwo��G���6v/�7���Q���T�,����H��#�U����(�~@/o�%�JAp��,����J��}��C����<�~GR�f/_�O���j%Gv����L�?��-���V���=�����/|���&�������N?����6˯�6���Ssw6�*'+u3*MOC��<�>T�J�����u7�>ro�w��Y?����.g4���)���#Zs�����._���\�/ܘ_�aKm~~{M����u(�y^h� ��B��f�@�����'t�f@!R� ���q��}�B�`Z�k J���O^2���P������J���s��Moϫ�j���jx��KV���[��,f!��}_�D<��/�/g�>q]��C��i획�0l��#Z��E6",���6�QJ쵞,�JE�2�)fӬ�ͤg<��(�l�9j�=��?>���s^ܟőϣ囌|$/��P����IjzU�a�5�7�_'����Q����0|��7��	�ȿ�������]����E���K�D�د��@♋��N �q�snJeET.F���o�Z��DJ�hD�TV��w	�AS�h�{�aC|��7�\O�m!JEs�u����e�q�yގe#q�Ǻ���戊|U�R�����.֒4g C�c�qI����1�^^Gg�W{��wk���ft�<S��~b�ޚ�'
j/I��9�����^Z��k��Y���sG���܌�d�
��IN������+�w`�u]�� ���y2�l���W3��Iޘ�U��d }�=�����V`h�E�Qۛ�J�`�t���C9_��LG�f�"OW���漸�S�,����k������ X�q
�d����E��	�LO��q5,��)����s� =�����W��I�q�ˌ~�De^�q�(l��d����V���\��mc��f��jP�h�D������T�������m�}Иs��9�}����q�Ĥ	�*��"Tj�����_��T(�*�TI�6UUTR����
A!iS�$�$`'q�q|�N��{�}��{�9Y��c̵�>�~�{Ϸ_�1�c��c�>/�1t�B�q�u�=�]x�Ơ_"X�Ew�f�g-#(Icǚ(�j�B�D��c�'��Tv���O�b�9쵵!GAc�b"���u4�����%#��Q\-�B�y����4L.ׅO7��^�
�B;��w�.��+c�M��������1�tḖ��(4����h���'-wt3���F$7��I�#�-�HL�fF�N?5]ł���7[j�T�0��#� � r��q��e���ۢQ�Y3�&�33������y1K1;����Ɣ��\6#� U�[C��T��HQ�@����\w;n��趚Y�r�ɯ���ū1�{g�I��6�u���J?8�]x�}�\ô�]�馝W��YQ��>�f��YX�<�YE�dAZ�k�:��d|�+%�{O�U>������J��,~���ٽ4�a|��>.&ĵ<*�����\��X�2�-��e��51��v�����+�na'1�?]P�H������ح ��N!���Q�s�`�I{�}�X�[�Z��t��3�b��d>�q�>_[��T�[�F��?��5�����/ҭ��ug\Q׮���
NâpW���h�Z��Y6�@I�퓺�80�lq|��\p�i�
�#J�դ�g�h\+��Y���!����mĚ�N���IK s��u��}�Ќ�%�
��ڔP?HEYj-Z�Brs��%�V�n2s��e�_����Q��h ���V�]�6�%e7���� CFٓF���iY�I*�OU�	��
j_�����"`Ò�{*1�=������]�9d|�nbT���h�p�#�i�&�x�c�X����?���0���ŝ_�ĹK����<G*8un�Q��s�}�Y�/ִF�n�axO��vX�;�փ��tӻ�7J���CȠ)Ow��ΩT�5؄08�Yc�۰:��{�A�����fD_�i��2v��U��0�6ޙE~�n�Z'Ԉ�o��7�����`��( #�=��q1Â�|��<�4�[l
{Ũ+5#�}x�X����qL���}qa4Ɓ_\֕�ĭ~rGJ��&��V'.�49���r3 ��v;y�,Ϝ�Z��޵�]ځ̜a69윀7�˝F|��4B_`"n�V�9#�tC�@�[~o���z �����i�=`^G|������\QK�P�CI�*����Q�f��]8�8����j]���^+����!u������%����V�(��r�0�E�0�i�b*��[K���63j��Z�����f�q�dj���#�)ƓX�3���������:7���R6p��G�(�NC��wT��R�u'�Q]L�3Ўj�ڔ��]�^&�ɻ���{�~��ǫ�ۈ���Ns4׉��lD��q��_"��T�j�\���#�������ALk�����Ê
,��̚�!#�2ݎ�W�\ڵhz*`�U�%d���?# ��E�kc0�⸎��ÞfC1�-�H�ܥĈ��.񹷑0��-��dk����]�/��8L�v�<f�=^�\�u}`+�hȃ V����0Q��%
�f�������X^�����܉�ee�|N���z�\d��܂i������V*e��a��|���.w�P4c��ֽ��Uq���l�g�c_m��7���:�=+7[U[\.N+���`����e��V3���͵��AƁf� �@��=��f�p)�2���iܮx���"��Ê�qL=!�X+�3�ft'L�yh*̊�Ϻܝ�G�;	}�cZ�Nk��D� `$@�q��H����q������S���h/}g�W�ݥY$�	�ȿ��Ђic�J3�5 =-�c�Y,W��3L��-������	�f	1+���
XpM���G�o2$�j�|���K%/�k�3(�|�Z�emC{�t46��2���@��׋��_���Y�pQ�ެp���"h�V#`��Ͻ�5bs������(��	�T��F�.�R��@�2<-��<H����=��ʝ y�)&_�ۆ��ݢ�v�ia�YG���o�ڣz!�+wf�e�\�ئ�][ϔ��Ev�4����{�J]P����v���FVO� ~u?$��Rv�ýy��Za��+A��"� bgA�Ҁ�"��royN�ֶE�qYd��#����GAP�JŘ�B�`!2�K���[LZ�a
>����lx�k��ժ��a�~�լ�E=��f����ƥ��L����x�gQT@����n���'� B�!qP�����4�b��� ���S;H�	��him]#.0#�Z&��юu]���ȭQ-�<X����s�>�g�5�� p��fm��0�e:mIr�	�|,���ik��f8h����s	ymqP� V�R�	eM;J��Yk}D�j�a�Ә5�3�86R��3f�=Sk:�섶혠�n"�͓.�D� �����4�B����U�g9]�ok�`/a�f�=6*^i@���Z�b$�"4%H.���NӏM��g��+��P_�9��^(��&J�T�KP%2����s�Կ�����t˛YS}L�Ե;�ۈ2���e����pÐ�t�$uD��NQ���`uŀ�[w=7482���ژ!LfZO@�"�~$Iw�}�Ih����#N�-ޠ�4`���@��bܪ���Uo�f��T-��Y �;���������y�Ǜq1����kh�Y�V
@���,�&[�J�5�Xs�6�y�LȜ�%+{ttjD��>�l�v��G
G�񩠐��|>QUP�܈�(��X�,'q�; ,(]�K	)�̤� �8�.i��pz*|����!�k����œ�j.Y����N�>,����j��1q��x6A�n�r��i�wgb�a�� ��oT�U�����z$���l��8nIﵮω�n�<��}8ϊY���Mg�����q�Mx"2�wD�Ϳ;�i���,^�.pW��NR;�$���Z����I|Cާ���#R%t�@sf��%?H�<�E$������ :u�h��n)Hޯ�н�_w�,��"ť�\��{7��4 �u3����i��d��:�g���ɭ͹Y�/n���� pz���'�o�^�ƚ�BaU�sg?�����n�h���'�6�ӳ�Q���Y�+|�X�`����_Z4Ff�m�*��7�j�#r��q ����w�`k���Q!H�,v�I�aM��f�XZ!k�c~t�Wj��e��j��
��]��ʧ��`��ڄK�O?q$��*�<zw�&V�RE��],͚eh�aA�	=��O�	�#K�k���������z-F�Z�#���|k	O ϠWy��`���k0���7��o��3���y�m�c�f"�r�q斩];�7{��UQډ30RP��������x���Y�Av��2���]Z�oRZ�@�G��rof��ks\>c�K�8=ZǏ��LU�e�µ8W�v�/[.��{��`)�"����t���ުR�����c]���������y� �u�]�:<:�4z>��R`^��p:����b��ʖ�A7��I{kI7Q!D	6^�J6��``�:� ��Wj���y�v͎��>�P*�	mC�j#�<M+_ԿT�!���\sʛ<�S�fĝ�w��%�@!=�<��.T��[Hz��Ͳn{Y;Ig�G��4�M�ϒ�dk�01�R�+� 6!���tuiz��ݏzBր��t���^�'[��1��w��`9�qVeQ�Yc
�����,���,ǿϨ-n��O��2w��dؾ�̹�0u�G��%�$��|�k�
��q�����t�HFk�R"Wz�	�*k�)�bz�����-&]�*!q�m�g5+V7*�J�iׇn�c�L�k}�z�u�F�`aL�k0�.�u�	��x6�^XZ������onT�������T~���E+\��t��b��Z.�ia�Ga�w��o��a{@S�w�]�-Js� �yŗ�����9�������{C�z����.��혩K�Izbh���b}�hq�Vw��P��5c��G��a�����hI�K��K�i��yP;m��LlYT.� @�F��kD�"�P�F�f���nv0���Q¯� !�q`��I�>�a�ȑ�it���������u���&`��_ ���b����|$H#q�o�8� �`U����|����W,]j����q�	�3S:J&:�"��֧!^�!x�y�)\.�Lg��M��߁ ?D %���D51>јM�q��G�F�)����Z����L1O6��0�p�\�+��axI���'��(R	����r����{�wt<�Zh1�	���e���e���h��<�3y�����.���>-��ӻ0b{��0�!�#s{DFg�>0fʖ	��{\��yuL�(,��Θ�2h�S��Z��+�s� ����!ɞ��Ip"�7q��"f\�7P_�iq3���Gm�;K�׳�׻�9rt{o�]v#�����·�Y֒ �-|�/�~���g�^-��[3�O%���F�"�cA '�<�_W�Bꑠ�w8���S#d��vtް»b����� ɿKᙖ�>�];��&���pԤ����E`,��TJu�är�S~��
�6��ถ�ň}au�Ƒ:���hv]|lf<�VR����sN�0��u�Ř���+y�9���L�a����I�R���>"�X�G@f��ū�T7~+A���̠��~��h�04�q6kAIa�֜� ������+ENnù�
���v:gÑ��k��9�l�*.w���H��j;�uS*��^��=����J��	��Q��̆�Q�Y��xp������1u)w*f�es!��Z ���ݵ�)�W�� ���4ֿJms�"����-�k&"�C�R��� ���x�C��z�A`i-}��	�U3�u�y�J8.�u�7��7�(|'q�2u��EF� \�,��Ѫm~Y;�tn����e ��I�ﬡ��j��t��>�ܵ�R1	Z�%@��^�w����J�����f���^�a��nx�E��^��k@�*8�=M�'���}^] �Qg�g+f+�������'wV��TLY����,+�
�P��ӣ.hlV��O��'��"��F��%�yF�D�畡��Q��`\S)D0Fri)�I�=j#�Ј���x�Z���!,�v�;~���	3����Z�&zGzF��:ޖw��i�������R�ŊDHY^�0����
"��1��br?_��!,����Ee��Z�}�x�J�Ɠߒ��.�K�/6{�����A�^JK�+����su;T�����c$��w1����X��� }X�np���� ���~q��D@_}���\lN;� ���I�E��(��{�;Msbߟ�&��-F�9�j!��&��Պ%�>f 9qWᔉ�X�s���M�#bB@G�a1J�]�(����>�� ���8hό8�n��Ҕ��x�6�$;�\��
=�CҴ�b��n����1�gߏ'�ة�w�Ҝ%�� ��2��@Ү�2��i�+ h*��xD�M�NG	��gk޵���PW�q.(��x�.�U;�us�ٳ�k)�E���\4��!����4o���YBd�����2����Z�@��Ҭ�s�֖�m�s��z03
f��в<��6&�Ŵ�6���-j�Z|�u��S(6�1anҶ�I�Ō�C���������t"�됬1/u3��bE�P������ыC��L
�EϚ�k��Na��w�3�� f%!tz��5a��qJiJ�>�&?�Z����`J� ���B��q�K!�u��'�>N�,2��[o�4���L�G�9���m�g���(�16>C��0�?s�0W��ҋ��G�?*KI�uIT&S	e-�,O�7��%
��\w��-�J�`V�G7?�!
��ӄ�C��E�!�=�> �n&r��b4�}"�k����n��V@�}�XP5N���vI�*yOK����������H�ͼۓV�b��^�3x���Ü*x�H���|!O�=�M��s�Ҟ���A��k�^T���,%���d#��W�t���~wRYF���Ýu�d뇔��b>fF?��լ>5���̋E�a}�^�Ҏ���������ʨ��ʄ3>��@�8�\K�����z�|?h�X��N��H?GaJ(l48�:6d^=��s=��	��5h$����e&^sC*�
n�Q"�7K�#W���ERM#���*�g���_����;.����U�pZ�D�X���ղ��,�P�?hZ��|B���@|����	��b�Η�d�	�#���<3w*�+��DM���\Da��m���f��V@��'H�(����3�AtqN��5�~50 �13���c\��Z3h���@q3z�T	�vճD���9,7;�`�V^�1Jܴ���!���hKb����=`N����º:|-"7���[��I'Ɂ֍WA̻�C�;Tfd�M
(ml�h�w�Vl�#����FC{)�o����y�V�o<^K׎b��z,��hu抙��|�6 �[w�h���Pn�e�����Ѿz������b���颦|���O]�*Iv���JѓD�:N����srC>�>_Y�2m�� �8�y�ZA��i�u2�ܕ����$��u��w���&s�Oi��m��6���&�n�_��:�������i�KVә�T�T���~�Q����Y[T֌�ř^C!�0
K�Z��z�R�dVU�X��r'V#$�1���LXXP�X���p.iA�ϲ�;&tu����˖�5h�*IGl��b�{HH���H�ڱ�y����9�:����i;��.U¸j?�j T�Y�b� ƌ��l��7M�C�"'��	Q��ɢh>�dD�9K�f��6	��KB��B�p���+�2s�<p��O�H��!Ee	��^n�KBɈ�ù[�j$d��(R �Z4�j/@�ԗ��V�fl"f>Y�Xh��n�w� !��̓���9�l�g!rZ����tuA�~;]�k��輐k3�ti�5*�ŉ^�]�g�C���tMɓ�SP�M�ݘ����h�L�JD�7AG��t�W!iw�U�%��fL*��H�݆j����a��'F�y��g���r9�k��D]w�YQ�+��gۣ%�1gMٙ��M�rww���z��U8i-�؊a�:e�L����G�kDN� �\�B��  �V�%���t�,�^�"P��O�����:U��r1�s:SU�����[g��')v�4eB��,������k��/�����Q��2�둾�{蹊W��4 �R�"�~X�v�=df�6Բ#��X��j�f8�h��AV�<<Vƅp�����m��A� N�C6u��ꎙ#	����sc�Y�:k�ZjR�gQ���-�h�[�m.���QD�$ؤ�YM�z�d�NXL��WH����_�K�3�̀��ʚ��ֻ�t�f��C�M�mhX�Q�&�s�S�k5�"��\�0�hzE͘RX��gr�*�8J��������C�:���-��!���^'�MՀ_����<��@D�?6/�S�-�6��u�{B����#[m��ќ*�[`�3�Q�^�GlS(�!����,̼r+C�?�_��n3�f����}��8:�AV��<֌��o�9�[+��|�v���Q�+�k��ǯ�d��m&�{�E7�-�;,Iqm�j��M\C�JE�Q08�#��bKp�`(���$�ǵ�ٓ2�������\�Pa��Rm^"����,����#j͢��j�2Ƨ�e��?��6�*,p��q�* 0��~�̼j�k($:�0������:@�-�}	f~���"���P�����g�h���Z�;��"�u�E܌�����ޭ
'Lc�VJ�M��E�L�h��p1���&�`��My�h������-89e���	a�E����_T���T4���1�N)��4����&�����'�m5���+��Ȉ+�8&(C*	�J7[�{���|���K��I(�oG����!���D�v���}SF�+�8BjR����JT̏H�'\L ����[@*6���Q���}M���=��}�N(��T��QNY�`�I^�2a�D�)$��k��]�m- ͥB``�ؙ�s�"�����'?٫H�u��7�{Z6����/q\g�����>�z���n�:�d���U
�2`������l�5�k���g��f
�� �s�5��k���8���/�"%i�<�=2�{����q���p2_�Tw;�/\̭�Ћ���|�#�ό����f��n�`�)�������q��9�a/L�S3c���R���G�S�>,ِ��>?�z�_��[�kz���S��5S;�F$}[$"�%�W�;W	�ě�Q��<��ݢ�	U(}ߛ%H�W���R�J����3&���˝��5yA"z��$^0a��BUԷ<+aBp��ު�#*�vc�
�t�QzFE�,z/�ܣdkhU�|i��S�6}��&��s7��x��c���=��@LH��>�1�FT[It�q�$/	�`��;Lm����Qp~0�<Y���K��B��f�����Ho��7O���tѨ��o���	�1��QJ>t�f�N��:aF��݂3Y�ٱUj&�IX4��L��W�G�:�Uql���R��jz���㾪�D�,i]Y�F��2ФjE)�$�:r��t�u|yǥ�k5Z���\�0���m��\� �w�2"�q_�����9<$n�9�1��И���˵Ҝ2���эg�B�!���
8�&��|U�&{�����̍V�)��R"��4w�=�>��F�K:�^���ٞ�q�uf��-qK�:!e2�q/�u�9�5J���-�ס�"�C{i�
Xo(�����	��
���k����Vz�ݼ!���T����0X��h�J�|���*n�|�\Wdn�=,�U��"��ϳ��U���>�Z)>�%d�i)y�������Z��?b^FܻJ2����ɢK[�&�H�Y^$4�&�K'�W�?ؐ�z�X���\k9=]A!�\c�xZ}]�@�|D4���&o��g�ʈdU)Z
ZkE�h��إ�Xҙ���o��ʠ�Ήq�wS7�i/�R�P�N��0�|��%L.#�����MP�/5�l� 2���&b�Q׈1����@��5"*V3���C���aL�w��7�ڜ�g���]�Hf�����Q����jy��̐�- U��vg�:��P{Ȳ�eI����C%��dyٶ��^D*	� �_D�*��@P�$m��������]C�K"�9�b�u��H\td���+�}4�$б"�(�?�4�:HNO�>WÇ���I�]d���T-�c�,�������L�����T���ր��V��d����/��J��v�@X��?ܪ[w�D�Qud��$�O���"@g�Ʈ4��XL�@|K�)~?�BKf��Ǽ:,��\��C�q��@e�´2_���D&�5�I���Y��Ц������$��|*�|���*kb��/�|��8�N�"~�N�sJ�Hx��>@�l�w�  �h���M�S.��Ϻ0�̠�:�C����K�`�
ģ�c�鉑��t*�K�ț��a��Jeϲ���D�K�j�M_r�t޹��h��l0��{��ӲSŌn]����M�B���bV�I���d�rJ���/֨�ӯ�t���'�m�� M��h͌��7��0��o�ف!D×�8:0�1�٩��#���a�����w3�kXnba����}Y�b�ikSib!E5(��˒���иH�&���H:�Da�,jB�$(m�TP���2�����
h1Z��h��F�����Y1�6��t�ݙz�O���s���F� ����#�`ܢ��B(���W2�l0t����뗙 �oc�N���*�\)i�0�e��tA�ga��Hf
iM���}��X����-�rI�MG��)�-���h�b��dunrҢ){� �>���v�E^O˴)�J<�8LPsz���2����ή���b�K�{�%���t"v��$h����=�D4^��ɜ�W%d.(K��-M�g,����r���Ͼ%i/�N�2��ė�&�;�����J�Ĳ���{�-���>sn����;����vz�����/ݵ�����.���)��&�	A
����a�w�b��^���3��]����L�p�-�)����� #�iy�����*_���	�hc�}O&&dR!P=�&r���x�})�Mэ��D�[�L��Y�Z��YM8*#A
V�R�cWW�#�=ʚ����u��x��U����)�ަ�.T��`��K��	� t��Q��k�����ha����!����L���ʄ�W�QXva�!��jc誙Ë!�6�	Ü��ʺ4�ϖ���n��.� �֙��ސ�V�s�*���r��a����`)`���<���k�$+��������m�1b���N�i��N�9_�-�L��꥜"W�.��ԉ�6k�'��
|6��n0��9,��{���R�z�΢J__�K��#�3S+۬�Ě�*�R�-(��GC=aj��f阭�+c��&X���ʟ�+]wSU�n"�j��&�� �(pc�ĉ�� [��Ť�`��J�.��H!\��7���QX)|�u�Y���h����Uk����(�B��V���Kd�J,�{i3��hw��f8Sc�H��l��r�;қ��#������f������2~z���dy���´������?���|����C�_y韨������������DL�j�Sm�Y䞘�d�^Y�@I��KD6uT*s-�S�S��#���� @k���=d�5#́+�F��muO
�J"F���a1�/Cc~�ya���47��EI=��9�Fq����c�@s��UC��j�z�\> ���3(��S^�C�ZE7N�1b�ܡϢ��&�*8�,)�G�E$��ZĻr�h��T�&ΚGŖ"�BR�K�H��Ղ){;�bk��eܾ�r�L���9�^�1�e�M�6K75[�
E3��Y��*
J����� �r��}�t7.[ʭB5k�/t�]���&���׉}G���w���[����%"��Я�TmJ�y��.V a�d����T�=YM��'��BS�$x��K�kJ�b��Y^U��f�^��̈́VߓE|������}�� �Eq���'o��ƒ�]���AB�v8��Z�_W^)�d��X�i���w��}kɐ��kx��߸)��W��ˎk<����5�9���G����^�����_�ly�����߲,z�/|�SG:�>���o�����/|�7����8>~������~z�l��e��pJ�LC-��ՈnW�P|����)r�K�|F�J��QN3�&Gi7�g͡�(�h�Sr,�6 ����!��|��Y/EMWa- �� �v�ficC��L]o�,�C˯��`�IB�dV��B�o���F�(�Z�M��(6�b5���M���7F���mi3��)�Ѽ^ete��޵��yf�0�>�l|�JᑠЌd�?W��3��Z�ϊ��w���`r�kJ���++"����8����׎5#�����=�z��@d�4�&�w�L��@@�Y/2��g`��,���2��1���Ю��l,G��ަ��\��dX�FBk�pt�+t���c�u5wnZiOc��1�����X����o}~�V��T\�������`�������F��Z�� �.�::
5Ñ�jJ�+��� \�rc���]�]���E�Y�,�b�WǮ���Z����P��f���|w����m-� ,��g�(r�܉}Y�����s�Z�����^��=���u��|������ }����;��a,��ȯГ����ϧ�������ku����������O~O�,�i6K��e<�G=c9��SMkU����I�TS���:yw�D-o�Qt�k�P!#�x}_�O"���,�^&Q�o4� �����'�@�=.
�=$D0v�3L���)-�+p�(#G�v�pDc�9ԯ�F$���1	�I�9��c�c�}����>[(��Օ��&�p��%��!I=kf荎3�	w֮5fuꦝXl�ᰴ\�`�J�|���g�'2�NG���|���Í.���#k}< ��K�^��+]E�mfkG�'f.\5���8Rb')|��pL\��vݹR"��2'L���V����nF�c�}صG`,#��m���k��+���x�� ��8�L�����b�cƠ�������;�����x�ީ�F~<�S{r���XV���Y�9:5b/�����|�`
|��F��5}�v��K���)��w�a�=JzM`���$�o�����4醦k�#_�:��{���\�S�b�m�n�e��7�G/�n���ۻG����O~����������>�iǝ����������K�ŗ��w��{~�/����ѿs��{>>��O��ߋTί� �`'��
z()aM)f�S�lf_  �IDAT��g5�Iw�"����.����~B�����n:Of,NhJD�n�ɣ���y��m ��Q�QW~���VL��]�&� Ƴ���OV����X
����ؤ�ƈ@�hJ�q7X�ð{�`�1�>;�D���[�_|��HCp(	�ڒY����i.��ťЊ�&�-�\<��|���GP�������?��-WU��zT�Kn�5!�f�Yg�0{ ��ī��Xc�4s#'.�J�hoO��u��UgzN+1^ujfAW�iǶ\��U7G�tG8��=�K��3�5C��ٖ�p��|4{�O�Uva�];�����:s�Z�m�:��������ߏ�t~�x�f~������vh�8��ą0�n�h};:Ȩ����
���~��]J��kCBĕ�| m��vzp}ש#��:9Cww�Bj�h���5s6�/R7�f�N�{U+z5Y��y��Go��������������G?���;�&�e�_W��<z����w��^����������O�W~�<����/��G�_)��Tc�d�������v��J�~�Z�������,�O͂!� ���ݸ$.lZ{`H}��k����M�7~��S�p5]E$~�R��q^$>lTj�4t��},&�M/���cg�� ��Γd�y�MC3��:�[E���ta	X\�'�׸n}Ctd�-��	�1o��d��lo��0'%��2�tJB�cq&$���:Y�.��g�w�=�R�\��+!q�.Dmb�y?z��P�����$�(���T�O��}�$�l�1x�~2��rP�����V�-d�1��KORT�4��9R0T��s��-k��#�&)�Y	���kF�2�ofNb��<��Z�V8,V�K|f�H;�ȳ�Z��v�T���۬�<�\�?��~@݉��hF���B�{8	5�1V$���d���z�ƴ����x!̇tm��I-����$�Y,����S�0t���z8#������KQ�Eh�����s�pw�܏������/���Gw��k������6���_��w����g��G�^����Ͽ�ߛizy��Ov�ףE�.��� K*&�����:�y,:�W�ڣ9����k����ڡs �a^s+��n;�"�)ļtiM3��q.&R.��*l���l:k��C4����~�JP�Y�L�lC%AgRdҪ\E��j���;5'��-�ᬱ�m�u�k�(]�H{%sN���W��X�������r��u����z�Q�g���.D5E6���d��VO�W��e���s<�vN������F��v��;��1�� ��,L�̂��*u���ي�4�;L�\ϟ�>�XA+]�~~M3�e�]�JL��#��A��G��I�f~~J�t/=�%���'��{�}��$fQ�M1�OE�7	���!Q�����"-p�Si�Ji��\Z�i��.���6�� ȣ��;�]���#pB1h�U�Bݬ��*H�i�R��@%W&�s���Ȓ�uGf.L@��HV���R�f.M	,��Q�?BQ��|/����	��ۡ��^�YJ��U&""0))5�vW>����m�}��1��d�X3�u������
���*t��7��<S�4M�,%R9P���Vn�L�^�Ӈ��?��w������"��]�NO9��p����_(����z��s��>|x�~���n�����ҝj�&Nt�sa���"���Q7T4�X#- C�'��{����с�\�8�!R۱����5�^F�f��:@��IkMSǇ�RH����?xM��I|�IC3Sd1IQk�G�#��� j�.&eڒ"J�dݐR-%��k���ՋWA܈Q�����2��klנEj����:�b�b.k��Q#�81u]ߢ��o�ϵ���U3?��%Bh�ᒶ0_qk����u� A���5�ɖ��=闿�4[[Q��Fi����S� �	e���
|�<N�1@�C͊�.p�!� ~G�V0#~Քͱe|��q��5�$�q6�\1�㌏�Z�@�F�?�nF�g��@�K)xZbipuh3�֭5%���ZӘ��9��-_yjxl�� !H`��?�րhE�f����ᭉPJ���1�6�С�5&5ܪv�����VN{Rf4X,I�0�i�0	=6��iz��I�)ڡ�����	!�@����x���Zlr�/��a�Ь�_>	]%�+�����&z[D
E��R���l�H�W71<T'LVYꈣ������+�ԥ-���i���Q43F��X���=���OM�y��:�g>�~���O��k�鹷��:d�8��>�������~��5���O�1=m�y~\����ߞ�ﺩߐ	��w��,��� �p��$,5�2@׊^\f֢e����g}�������J�h�*�m�}ۯf��6j\+���`�������@=6�1�QZ�)o@����J���gG餡�1i3QHڄe�� x�!�����e }��^��;��H�Ecl-��w���D,J���FkM*[a4ʝ��{/r�N��H�2H��O�T������k0(onIa� #1�Q��o��a�;������CѾ���y�̤��ᴚ�UH���E�F�iRw��� +
d- B��t-䦾ah�b�# �Ǘb��R�`�Ó�Ǝ�\���X�X�fB�Č{��/�ܩ��*f����q���|Uw�y>/�dc̋y:6m���T(n�ڒ Fi��Y����]�зaC��[×L�#��b����XX���Xp����0�W��Fs�?��x�b������%��'kv�BQBê�@-jYU3��F7���g���^����C�����ߩ���7җ:^C���oz}���ɀ�������ٟ��O�/�щ��H�R���=�������"�nT-i�IT�匉���V̵����+��4f�Nk9�+9��>�i�d�#/4 �h�C�ޑ� ��mL���;(X��77fiOp�}��E�V�
���I��T�Ĥ1��,n�vf�@�B����2UY��'ن�I\Q�z59�7�5���T�l�#��0.3���b<���ML�,�8�U�9��E�@Y��ςQ��^���\0���p����=^C�~6�{q!�}�E�we\�;7�IE!Ŧ�J��s�2؉f3Uc��kK�����cMW4����s|u>�W���]���9hQN���ؕ~����i�Nu�I���`6٣v����,Z$��F`�lX�S|�M��s�ék~t�����V�`����@�]s�X��8.�R:�]	0�Ep�(�Q���횬�ӊ��ȍ�!Q��DN�Oy�N"�Ռ>�^�ʟ$�د�o\lf�;����<�>��˳?�v�oz������:�[g�>��?~��k��2л��}>���i-�f1��TC�z�F��Pr�~SSx��Q'�_�xH0����7,�M��%�/�x���e8Gir�IA��\gу�/�<l��5�Y`���fj	��W1̩��,37I��A�Z���cs�S�V�ӱ'7��6@�Da�S�����
���Ip(��-a��,�:fs7��P�I�'����i>_�n�Z�L硦I�g�+�,&!�#�%����D���,*>rBк�׀Y���d���@(�N�q������dt�
�}�n���P����z�I�'�ps��ijB�z㳭���IM��OZ�L��zeܰ�oY�΁o[���täj���CCW�>�WL�M��<� �{@�a��%��!��0�4�\�FPW`�'�f���Y���݅���?`JҽѮ���)�?�o�U��l�v��-[���
��nM!��@���4"+N�Ч1IM�L��f���;�\�OЭ|/G�=���n���=�=�C���g��7�����_6C�C����I���?�������֟_&����ā2��e�`>LA�c��:pJ�%��޴i@�8Q����&�-d�i����9u�C'����m�C��(�o�.��R��8��c6���U��{�,����TB�NV���"r�t[��O0td����Է��o�2���<L�SM�8J�@*����m��a���!
��1l�f�~:�ܕ�ZE-k˫���7����"<3WL��\K!2֪�q�*�P�>������,2���MƑ�#������`¶���j���4JKYq&�;ES���v�Zz1f%��
@���&"�;?w��`Cv��``��6'�vu��Cp8����o^�^�ԇ1��Y7˷�׮9Z���C8h"�O��B�ե��MJ�	ꬁ�]�i���X��d�v���ԍ��{Pm����?��xu
�`>���'���[Ҟ&M�U7��a��ٝW�ػk�!u�Q����bj�IT{�b2e����VUek2��9�O�~u����������������=�A_��1t��L�����������G�y�"]/W���il�1��räѱ�-_�,
�{���j�U���Q3$\1���Ř�^��h�� 08|>p�6"u&!\2t%�-��͂�ҹn�p���DCԠ�b�E2ӽ0r[t5B1������D�+C`�L�&P��0�*��60A�������10�����h�n��y��LxXKb��Q�g���D��mg��ee��jD��n^76��6Ĉ1@M�]5Jd;���f�ւ j��o�1�J����t�c
�'��/�|��{�#�@��f�p�n�-�F��z'ʹ\��]Ts��ߌ�Iz���&�Ɔ0bxk>�f�o1�/q��;��ۥС�6���P��oԎA�v�����|Q�K�A��Q�z��s��+Vt�3����oi5���m��K1���K�Ef��qF�Gky6���P3����ڄ��j�mX" �r��Y��	�Xm#���;oy-�tH#�Hb���k>�NR����3��^x��V�[���1}��W��_��o��~�7���������ߟ��N���6k�/J���mJ���MӰ �K�D7r��Wgէ�J��ɺ6f��ߊ���p�s>J�w��-��"��<�a�q�2I�H+#/�����̌��hT`�v%2�XȋuSmb&"��l̤�6�k�(I���+��L?�a��&cj���͎��V�
ps��������p4����[)&��)���=������Ka��*��l�V��No��VB%4��"�=�����C�}ݛ��U��a[~?꠩�F6���v�g�B�
Ke0'�ܲIX��Y*��խ�\�F]��^;pM��M���m2ʎ`Ä¼2�����^�������;�ay�!�3q�KL�Y��� Df
�2��|G|�>!�Ä��}S{7��q�a5C(1q��	h,;�oґ˃2܆���"l)�`I*ˑ1�*Q�2�Ɉ`�6�X_��h;�$(/F�{�)��U!��4���YXҒP�ߓ��_��~!4��h����[Bk7���%hV��$���>�^������Sf��,�
#7�����x���o�����=����ߚ���羚���:o\���?�K���_�7���~�����>�C�\�ʽ\��iX�{�\R�J�#m8 ��@tf�B��`� �Vw�bC,�%�m�����6�(��Tb�3V�}��A:/�.k)w�
Y���jK��<Ka'<�jlk���]b��k)Iz��w�7n�`�_�ّ���ݘ:L�	��6���Q(�*��Ã1� ٭!A�y]�y<݈��~_�z��}��r�''��6�G4[`u��fF�0W��veR�l0h�>�����9T��1$s�H���mV<�HB ��f�S#B��`f�IV�5�
x((���� k��V%w*�����Z�ō����JW5#����_,E�TP1��1<k��.�by]z��]�x���g�}dV�i��{�!)��3�'�V׀h�f�h���;�.������{�l��*X��[:O&�j��J!Dv�N��MZ[�|��i�'��M�G�8U+��!*5Ł39����=�6U�90ԒR0��S��Ҧ}&8%��
y<��L�"(�`�Y���U�
�M�?4�u�⸞�	Ӹ�&r�y@��(z�Vt��x��έ����H�;��ŏ:���ED96L�nZ���w����������5o������5�����_C�����z��O�'?�y�腿���]���G���܎sq�KL�yqgʦ�)�}U�wVBքZe"�.`b�ǖ_l������}�#��ĭ����3�0.-ia.����@��'���(��*�B`�Ʋ?/����H�5k����K�t�K�)^��v2f��Q�`�Ed}(�i�6�kƗX����9>��^e�nY<�8��Y��M�x��)SŰ�#j5`�I����h��c\v�m����ʅt������p-(�^3tנ$�:>y'01�ca�����\(�7��/�Z��y��b9SS�\��jvlpE���.�>�	����/�X���t��������!0[�c>>U�K�4�Ӡ,�;���Ǒa��ʐb�S�s	����7�^E��o��c'q�Χ#u�~��[4�t�e�����g��3"��qpl�)�-h ,��t{3�^��w4�بiaӅ���5C�
wF^�/�C�>F�_��%>a']��X�ئ�ۻ)��n~����_�����"����M�����_5CǄ?��.s|��ͣg���6��ϧ�_��!<�)� ��ԏ���R��TȂ�	ȩCW�cD�w�,J��60^��͕���\j3����B����A��#u3V�A\g�cH��ƶ�t&�e�Y�0�cR5� �u���cU)����ѻ܆�������S�J��:��!��]�O07b< D�M�[�Q�fŵ="�R�$w��~��̟��:4+�Z5�Rc	!I��vhx�
M�,�Y�w�.��J �0��)��B�pu����3��iU%(�W&��Uh"+��1Ɋ�_+n�"�ۙ[�.�4�IN5�Ά03�q��H f�k��
<�1	6��s���-=	������ɴ�&U��QH�)�����v� ]�����J� ��kB~�:��O��.����"�h�)M�L�0�A�����݂˧e��'�������H���Ee�is�=�t'R �僀���lЙ1�9;�1?T��C����T/�Ǻ\��99~-$�Sq+���_+<;K��b.��j謼�ɓ�c�l�s������?�����ߥ��7�����:���������2��������M��{��������H�'���f��,_��^"��s�	�(�֦Qded�@��ȍ8ۙF�bѲ��D�m���AW��m�m;'"���#i��@��PQ+���6NaV��b�(��m�֛����΁7��L�	�/$\̳��:%�6��.];hB_���'��}����T�x>��k���C?r�5#�n�%/L���I���Oi3a��A��I��T�;�VZ������f~J�	�ȵV�閒��	m�Y*2�5�f{J��Z����z�����9�Y<�;���i-v���8��R���(Ym�|�ҸV]/eǈ��G�@�3�����k�,�W�>u�̓�lM<�u����
M\�jc��9Z����1���ʭ[#aM�X]9Z�%aZV����<����Z�t�óM_q���"��#N8�����Y����'����4[@"��Ѹǻ�Ňj��� 5k���A�����2�c-d\3ů�E e���{C��of~#���'<M��q\�^��u�dw��ov��S����
�������1t>�������L��l�(��"�}S�@D̈� Dbt9�t׵��g)g>�ɧ��D����?��f��g����>Pd���+���F��pO��5nb;ɾBP� ��Kmq��L�a���b=0^����k���}���ǤxEW�>��H�3�Ey��`͑�tiMd]֓��¶��6�гb�P�<��qٜ�g�{z�����ip� ��a~_��Z���.\'��%|�� !�U����Y�2�Ԅ!�\�"�j�L��@dR���B�+��"��#{j�v�&����R�=N;��D�b��G���GS��0g�a�}�����SR錉�B��]��UK�S�S�紕i��c'½D]��I��nF�+x����I6C����\1��[�E��2�XO�A8u����Si�hV�ЧJ�����V^Եҥ��N�m�O��|�zsG����r�|�s�f!��ZD�!�S��,|f����.��b6K~?���|)��n�Y���|X���[�â��q�kDγ�<��Ks���A���s�ɝ(.ӧÂއ�����{;�r��oz}���)C����>-ƾ����8�;���TΏ4��[k�F0pt 1�����Q�ś-W������8��f�&M�j�(�����ơL��f�	���2	�~͐2qE|��DZ6Q�t�Q��%�EY{00�����inBk�o����0+�� ��1mŉ��W����6�J�q'��䫣d�YC}|���N�'Ҟ�0�v0�Ƒ�������K��2t-�%�a*$g�U�J�-��X�و��{H�pa�L�O�s�u#TEK�� -_�������5a��j����S�9��M+V�����p'V��D��|gBC��T�Uf��:Y�o�&�U0�V#��:N��s*lI�!ÿJ�ݰO3�L@�@`�"�S2�,:}�}���(��([C�a��1���0�mY���Ь@�f;0��c8o��>�f�^��*��.�}���Oď���t���p�Q���+�8&��
du��1
ݛ���	�C��G|�y�=�9մV���3Y�x�k+怏k���A��g13��i����m�BE[�rN:��-L�c���ͧ���=��.�}}|���}����?�n���v�?Q{��K9�!�3�Y4@m�v�ཆ��{�Qw[��Q�U�-��w�`<H��8�(�"R"��R��������e��d6%x�>C�
�o����f�V[�ig.��k}����^}i��x�7R�T��D�:�r� ;2eQ��T�m���4�I���v{���檀I0(���*�����XCkp��nH���i�
Y%�CXh�5Ba��Q�0�G[�3��w�CۣRCohn�RI�<I�O&���H�p��	PY���	�ac�L�`�HeC%:���P	8��M�#zc��N�p�'�q��`�VŃ��3��q�b��pd�EYΘf�{0�UaN4=��������If�]�Me����@`][���f=�S��H����w��%��%ѭ=�JZ�@�%~�n7E��?
0i��u�%lK���gV����)֏�٘��d'��
�0�ݣg��V�==y�%:��[�ᶉ5�YbEK�J���\�
��!�A����%�3��y�����9bs�L��Εv��z����[�9�i��i�)���3���Ci3wQc�p[��R�k��s�Wf��/N��?t��}���\��ks|�:�}�{���W�m�;_�Ŀ�����w,0�6��=�I�ڮRK桐�.q����t#O�r��T�j�#u#��:��I��%��,��&���m =f���0\#@��^C�2�3n��K����kE� ��tO�*V�cWn����R;�?�ӱ�,fR6�I��pMflf�-���+o�Ό��m3��0�4>�{:������r�tKu���l���TV��:��U9Y�C0q.}7�RNU|�'6AΓ�z'��_�8�g��*�˳�
d�S��'*�)�l$��������S�#H�Qr�F|%N�g�
 '֬8#_i�|ޝ�)��	a���5�n���k��
8�΍=8��,=���Ls!d�R);��rLիL�p4ۺϊ��!P��=�2������q��v��CA-DbL��#�{�GE�o�_��.����uy3W�=f��Y�UF^�Q�0��*=\���~6�U�R��|RZ����0ef ��TA0f�x�v�qz9��nXC\��x�1~A���,��%ca������ځfX�-+��|�`�#��d?8#݄�ȯ��͚�?�x�����P.K]��+���iv*�V�OlO���R�2AT�a)g�����5��.�S��p�C��sLVN��v�s�wg��_�}�����6��-��ua�||�'~����t���������~�·g�� _�j`@�fJ��ZE*�4m6 >�3���&��oVŝ��~Bp��^��]@4��/fu��� ����m������m:Q�r6Q�"��?⮠��Y���gL��F���Y�0�Q��I�Ed����H��[�WG 3��0� ��i��/����FR�%D�<V�Of�QF��n������y5�����pAȨ3sumn:����d�n�>����||�Z�M��)�, Z�����E!Pj��)e����j(�,G�PX3:/�5�{�b:H�Ct0t(m=�'�����T-�\��F�Z[b�0_g���Ws|5G��P�	f�Kn�����,�Y=��$�3�G\�~-�u^5O�7y��\��=�A^�I}��0�P��=�Wr�f���๾��4G�x�px ^���+���$Ѡ\�,��X��v��J�����Z=�MȪ�0�\�}��R1g�@3�7����"@����E[��G��?�����{/}=��C����P}�S�8�����X��?N���ʵ�HL�����b�J��˻���$9��Y]�ޡ]���/�	�R�ȓ�Z��k]�Nc͓u�Z ��M\�Gjc�ƈ� ͚�G�	�`�\þ�s����̆ȳG��eW��-����d�r�t\�3�fib?��0���%y.�Z�j钺�5�y���6���*���Q*�b�B�y˒�
b~Nu��eGb�֔���*���<\�}���2�����9
#����}�%��|�<m\��Si�e��oi�hD\3f�p	Z:=pd�G��%����A���T�ӓ�z��&���"�Y��n��#�Q�fe�K�:��[D�2z3�'���Xm)�]�G�Q�"����֝2Xg`����ڱ��f-]_�kꭅ@�`7��>h�aɪF3�b
c��`������Hy[q˙/voע��J?�������o���3�d&��!����W��0��v߸�g[�֣]��D35R�4ձ\��]@��!/}>2S^j������Z���]��ښ ��/��b��[�����eg&�I�y�y\��4�o~�q��~�;�z_7�����E^{�����ӟ|�����g�N�������X�}���v̱v�<�V@�f����"9��];.��f�`�=cK1G`���c����_�z'��[I�d�.��4�ۂ�-�(�gT`�t{�;r6%��h4�B�OR�+n݊)O
�q��YL��y4�F��3CKU��'G�;hu���Cw�;�]���5�D%m4א,������M����س�|^���Y[��.��*~x^㳚yĬ6�J�V�ִg�'8�v8k���U��1�;_�Å@�a��$GF�K�{�w�4\�6�93��L"���)���M�i�s���2�Oiw<��]:$�`c����nX�҆E�>W�f�K�W�X�D�yM �$�$��-.8f�{u�|�̔��	-\!&�Z�jw�x64ʊ)��SZ1��"p�E�Ͼ `����87F�,"|5�:��,{�M�z�h�����(��̻X�͒k��0
O(T�4ǣtZ���JWi��f%�3�kʶ���
r��.J�y`�9�Iig��l���F8p����O��}.���ϫ2re��7'�s����8M����Ox_��}_]񘇎�C������::<��/�O|��,���/0y�DS�E󛔉��=�c�EtJ*�1����̻#4��Gf�L�LIׂy㛮G%�&Q4����iP.�i��3Af.K���׌�ivS1%D�	I�H���,�Nz!릉b#͢��_��!�Z�����"��Ԛ��k/�L��][��v7�4B�Eb�=�w��/w��)��ر�&�[��=�o�ŧ}y�c�&!�g���|߽N���Fʭ(%9@l�bG��F�Y��c.Zꘉ��@�o���5G*C��`d��B�^J䑩)�
`(д
�,�)��՗Xw�f��"k3oO�.r�I;���j!�����%B�n�\<�a����v�ϼ���_�9m}�͵%�'�B�3_=3�:�U&�P�T�G׽�﹒P�q�_�ԃD��^ph�M�5����pĻ2k)�k�iU<��������N,��}��$�a.<s�Jr|kf斁$�M�1�K�}V�h.��n�..]�b{�\];ZB[�52z-��5�"]�!v�D=����ۚ�#xSt|/��$o�q���}е"���w���[��_�}��g���������3�R��>����t��}�//J�?�H��R�6�3i�M+�RA��Q�����s�F��fk�SB��؄>�G)]��`� vg�N��!���\Ւ4�˝��s���o@���cD��,&�&���>Z\��L>�S�N�����izM���%Z��N��E���~9!�
�D9k�V�����bN:��&K%�5���y�:�����8C�p�NF؏`h%�L�5i���qa�e�ιj�^��5�Zj�Ko��_34�/��n���ay���[xҠ$>9Yh'n�"��E3R*�<��!�s�.0�R��dx�H�L�"f�L�ʑ	�:��O�[E5��{*˟��L0�*��L�j�T_g��Qj�]C�u�9�k�m!�^|���-���|�}LAM8�0������&v���I>��*��}��ձ��5@��OӀ˩@���\I�2k�糬A� (-�Z �)�"]�drT�'�vՒp�]q��5 C�V�����
N���"\#:6�)Z�~3����I�j��H��\4t,U��,�gv�pB�dM��#��@�jQ����V���1H�-���N�/.~��ܻ�����}|4t��������ş{qz���D���$��-�XU.� GD�FeMY4SmɝSM�J��ҧ��C���������MߏRY�D��s:5�_CWd��&6Yw%��tj�5T�`��BFLͤ�L�DÔF#]��{��'VN�d�U��$�4���H1I��G"��W�)Ҍ��_K��:�=�o黑�g�/����ߙ/ lMza����r�+�N_�h�Yk�kᜪp,��Hk�kmr��n&z�k���Z�������))?w�㒯���_���:h���'ZI�Mx�hc����7v�:`����nfo��	ڟa�Yk��\[*x*^�d��3��K׸��߰劥B�࡙vW��/[��p�I&B���f��%r��j�����Aq�!�zt嬸`Z ����w��$�Dd"��A+��O��#������-V�C -b=��鄈�"��8'����}�-��S��K�d��R"������22��� H��pݰ���/.�qf��ƥA�a����O��M+�V����1;������gir�z�X.�����H�����u`�nu���d
*ǁд��e#��/�އ���g�������7�����}��׿�)��*��o,���K;�-��0Aʓz�E����),i��Q�U[*�O{������� ��9�y��2�g�G�jM�0�5jRDF!F=�$8�g�5�,��u�!;I��c;�=K�b{�!i�2�RLL���;2��Y��$�$T�V#vB�w��Y>8p�� �SW��ޡ�[�Xl���<X�����a��U�p� x���g!/%*_������ŭ �U�[̘�ҹ�~��+mO/�G���'^N�-4��h��nγfV����wt{7��e� z�	��y��L��L7�I
�D�8��d3�a�B������T��ا��}�@D��N�ST��.m��%H�8��H{�K����r����'Rⶋ�{'- ���t��]?�᧍K�!����@�
��ʙ#�#荿�&8�>�8$m���_�yˉ�մ�N.0�P^,�ք
��kB_��4b#T�fݭX�#��'��1Ip��N��c}�R=��l�d�"���3gr!����e,su!D��X���Ҡ�.A�Uc-��BK��-VDr���p��8W2�Z�L"R^�ޭ%\w�B�e��5�\Cg`t��[
�eAA!P!sf�������<Оb�#1#��ig�G�'�������4E�8}�n�u����������}��7����7����o����/3�N��ۿ���=�����0	2GB�?�(��E" �����������]�V���t���F:�(��V�{W6���U�Q���5k�y��M���r��|����>N�G	�	]h����NBT�@¡^�E'���^�}�������*��q�C�M�B����&�}��@v]�u��'^$S��s�W�@B�+
�d�t'1\N� ����<=��i!
;�/���O�C?�u�_g@I	�Bjs�� [���c�UP�&������ih��Z��* ��@:�z����K��X`B�^���F�k��ɛ�(���V Ø�"���ڔ룖^���S��C�)����������Z���~/׼U��4�5?{��1��'�́������*�t�+�؃��1�$9���.Y�d��X.gv�
�LښS`׺��Z/<b\��ي�0=�ׂP���r �K�,2#�fP9�ߔ�����0�{%���Y�nD1Edx>Y��B��y�
�Z�����iO�u�D!�s�mvߦ���Z�)]p#I5��h�<W�[�w����ǥ���ݳo�������K�:�a��o���/�������O�6�w!i�נ��Y|�-Ȍ=��b�^���AcQ��ms��I���ދRw�����Tb3wՒ:�lML*�eb����M�JLE��lr?qj�4�>��礔_%jKC��jJ\�gl��{��/����)�Q��l׶��[�����ݴJ9jh�q���}��oK�}��z�dF��ˁ�!̳ᓦ��F~����j�F'��!���7R��1ccT|镧�7ӳ��1͂˞jP�k����,n�Yq�~�� �~v�^)��'X�6���s���^"^K�B��E�;׺ꤘÂ�q�̟<a�F�ŒYe�ZDLr��2a�#z�](�&���|����M��YK�1
�B��;k͌�%���ZDB�X;�
:�w��}T��k�ɘ���'�I�U��?[$H-�p���l�?��Q�~�<��$�q�<Dk4�D�Jv�-B��p��� �{+�{М���͸�T=��-{�,{j�Bռ�Lڮjt`�5פGk&�=UXơN��w,)n�Z���bL�:��8U��T_oj�f��A��&�ql��N7���~wf�������u|C:ǧO�4�~��{�������L*��*�`�~�چn�j@���_��i}��FV�k;%dv�L)�M1���-`fi�7H��Y��\I)�j(I`DQTD�I��J�fM�$�eA���⤂�"�l�p�L��$3�j�j1�r)p��km�#��!$�c�5q?i6QTS9�E��1c�n�K�%u�;��[:;�BO8��o��bm����yY�����NZ�hR)R��J م�"���H����/}�C
��>81P��c-ڠ(�N'H��I[I�ڮʖDR2EʒxI�rxn{���c���9�>�v�P�����������6p���{䁅*�%v*-K-�8]/����i��yj}a��8��|o]�S
�H����oJGٺ.�
�̊���@����8Ѿ�F:	�?�?��fQ�$��⮒�EU�7��U.u�$��\���
��[���bN�������>{7�tyy��q&׬�r��2�I[�g�}$ga�I�5��X�ܽ��z���z�e･+�I{#���lU+�L���I��N�dn1�ų�	t�䦊�x
nM��}O�N���@����r����V�͓b�,2��d�9�H���t�7)/���m�ˈn�n�]�D�F�A��)!���Px������h��"��+�~�?�4� �'��y����������n�O�A~,&s[��w��dBD+���4�Wn&�MB�}6�-�{�h��]���C�L5C�u��z���Z�ZNb�Y��X�z��+O�ɜnЄ0����4Z�����U�@��H�ĭ����._Q�	@�y�:��O�����d'($Fb����u�

H�J"X���&&v�21K��>Z��%,i��h�4deG�5��"��X��j����U����8^w!;i�u� ��Sb�Wtʲ�\精JHaz?�'��(��,V�Q8j8��u�\/�e��B���}�FoA�{/)M���uy|i"e[G�vV���1�:�˾�7Eb�<���)E)�����v#��_���ngF�SI�i�{w�%���c�9�3���8ȥ������ᾍYdB�> V����F�S�dI�%i�z��}(�^��ۼt\�Nי5��Uw�<�{�MV�F���Q���LY�<��k6�����)M����\�8^���Q+rg���B��F�$#��JkΣ(��P�B��wx���.V_�����ӊ�?pB'�'��7^�*�ůB��O��?�~�N:�ѠxH��LN���d�0�۠��Sk�֛��	фɁ_�m��[�w\�a
�/�5�sL	��U]�l��?|ә�y�=5�� =tlY}y������U��8Ȫd���7����RӜ'ʲb�m����� ���N[J���3N�q��e{\(�
�����-��.�� ��I��J��A�}�)���Q���[�Î��1QԣA-dxn	)A5��IEI3W�t�)M�+
����-kz�:�ߧ��TASr�͕9�9ۃA��%��S�K�����\Z<nO*�Q���qF�VS�q<K;h����'���0.!�>�s%��� �D������a� 푄�a
yk�"H:@�*d?�"��9Y�B���lѰ��>"���z�N�ٜ��JsOeM4o>���9g��8�@c:�%�n��_S�̔
j(�ݍ�N{�ŵ�?X�w_�L�����}ʫh���?��Q	�9�I��4'ɔ1��ߧv��Gg`Xf�D$�ͳ
lO��{��a����lK��(Qc��$5)_��n ��kxS�e��5���!t�=�~������o)�X��?�J�>Є�*k7*s�)���%i���YJ���þ}:�>J�B�Ek�czH���Ff)���cL泿��!�q+wV!�	���ロq1q��q3f�؅b`��$�`��K�,����Q�T��تC�Iq��T� M�&�ȣ����,�AW��W���e���1g�`ݷT9PT�c�O�)�4
�A�7oѲ��ER�+q��v��o��e��Ls�q��������Ш�ԉ�@ٳ�F=)6x�wܪXr,F�~�0��g6.���I�A	ko]�>��kLi�YQ0���Sᚵ$J�u�@����2��N�D��(��Q�%��8��t�����v��<���1������|�5{<k�C)c��Dnc�#�ȱ4�Ŕ�[�Ρܿ��i�HѫM��`-`����W(���u�"7H\�ŷ�7ރpR�K�\*�g}�S&����	ux[4H�wm`��]���םt/�̙�����X<02.��4�V_�Mv�c6�/����b�n�>���$��ae��b�P��U���^'�%�P�Q���<�`
k1� FS~4�F]Z��MAcE�ǟ��=r��4M
��܀f��������P�a���:'|`�~��	�q!�'�v_�+�[��<Aٳ)QRW�]�@kա���/�u�}����&�A���Xx�A+\&����ݪЊ���$�4`������ؠ*�#���s�=�O)���4!Y�H�If�/���8$�5Ťdnnv!�D��aP���:�>���2@��\S��4� ��,���0�Ʃ��3i���X	u��+���2�J�/�qԬ�՚����6lx�\"�J�4��u��{�D=>u��D�
[}�<��b�(;�^'��$�\�]�Xi�ѩ�P�>�����\l2O'c5iς�z�t���Z�I� O҃Q�X]�U��'�)
Z)#���R�i��|j@҉�d~y!(C:��.�j��Z�J���4�k��g����^"#á$4�^�2$��M}[#��"��Z�����T1���!�+٧�{'N?�Q�$J��ΥRB�����/�_ϼ��M����%���� 7'j�C����.M�Y.����d��d釪!��	���9Ú:�I�Pi=�`���n���z����r��PԖəȼ��M�|jSP����5-.�\�r^��FOTQpJ�zZA�����`�H��h�(fc�Sԁi��/7m�]�7q՛BcW7��P>��	�.b%��y�7�uiHC$O#S��]�z��[��?��6��p>(|`�~��'��?xN�����������/������%��k4��4;�R��u���ZtP�w�ԥ9�V�HW�m��-�؉Uez�޳�
T�2�%����B�Xד�K�Πپ ��]�6��"�k�l�$_T�G,/��`u�r��j��B�+�N��_"�Mq��e��k$�1�:j��
�zu�3]%:B�q?�@E��i��hh��R��,����C9�z�ht��w���,�ɿ��������ٚ�T�#!M�&b�k��GF#�?��y��zL��V�j�\_>+5�(n>�m��b���5��<zk&�s������j��zZ�8Ϙ�o�o�G`e1��wPWi��K��a}MQ*��Qq.��}KeX�m?*@�Xt���\��F�^�7�C�_�ە�\qF/�;9S���g{�ɮ�R�D%>kώ�[�|��Ǟ��'/*�{���L�V�Q��i(H]-�\��p	&y���:$�n'�+)�-Z�4G=������=y�
_�2s��G����ۓ��X���:��B�1��:�q��"<�7f�O=�0��<vz��&���ͮ���π�4��1.}��j/m_�p������k��%�L�>0B'<��S��+�.][�]S�]�����OQ:T}��]cMa����Y�(Y�Z��-y1�����"��ķ�<#��L��L�I���I��_�t���?�U~���X�t��˛�}�1W���u�l�V�е)��I�8&9e0�I�JcYY��4�����[�θNa,	+Bu�Շ�n-C-��� ��Ne�Z| ��B�6IR�n�� �}��5��8��	�C�~�n���>W�]��7�_A?�(Z�`��O�^��FnLS&ƾ�c�q�%Y\�j=��յ4��:����~�[(��V��H|��%��8���N�^�pe$ZM�0�� {
ְC���cix"�iw��̪_�{
�<e�:N��e�d+O��x&��a�TT�P� ���YH=���|-���SZ�Nd�(�V�9QԸ�疆I2��n#��	�.ԥ2�n����h`��9ю�� ���h��dD*]�Z�T:Fqx�����ܰ���u�Öd�'�/�C�S"���d� X��B?�0��U�I��yN�a�ӊ�d�T&��;�%kIn�!������ڻj�9�8�i'7;��?�����o���k�>�C�(G��J�߽ ���l�� ,��nH����D�Ik�w�ĸy�T ��-ɤ��tr-����Wj��q�2��r7��D>jז�P�B��L�畿퐗����f�J6��mD�k����)�
����&=�눦�Q�g:���K,�T�;W��Zƒu�*y"����(j�Y�d���;l��al�i���3+;�X�b��SB���fT렄��+D�[\�MGd�-c��zM�)4DN=�:�µkW����^�訞�]���BCB�
={�����2٫\��J�C���
�btn�Vl�5��k&d2Z���R��t��Iv�F�dL�Y�$o6uA�61W����qtM���K`&}>.��z�4�����$�Irc�׮�#7����o�K	VerkĲ�B�EY,���k�\��O�"�k*k������?v����:��+��8i���p�>�d�B�N��"�i��PO	e�kG6.{�D�+X,� �`�9�A.t�v��kR:j9������6Eɱ���魨���s�s�'�������],͵8�d�q�i�&���5���(��7��=.n�^�Z_��N1u"r�2����_=��~�������'�4|���	�ޏ^����B�^���m�����z�C!e A�8C�Aݕ*�6S�+����%n��'i�g�v�o�)Li���4� 
Q���=����UL�n���O(�>	O��R�M!(.�L�$�I6y�E�f�m`m�e�V��A]��]�J cR{����ikI��$ܭ�`��o$�\˙�� T�ݲe��V`�FژG%�j*�ز>o��EA���%t!Z�⑩$<n�Zq�ry]��%{�����{޹���1���1^�c����Z��b
�2OJ�(D��k�L����I,2�u#-����nl5=�P��"_�z��
��F��M��#���-N��սU��w��n�Jf1��K��[J�/���$��]�:�͖���uI�q�q��Ե%����I	��:�P\���Öm}�^��0	w�]��:%�5H����9M�
��V�e{ۄA�(PRIc2$g�+ٗ6���I�;�f���
�mu���� �$���s\C�O<{c*#\�48y'��;�Pb��佯_\ir��<�������JO������"�����c��(*��W7}��y�ik��ҵP��\/�;�LLCY��5W�<&�@�=��-Z��j���a�[5�p��>4>pB'<�ħ���/|.^x�~���zI�P%�[�LbKNj�ԅ��Z�dnVw|����Wvg����<����w�b�������a�&�=mz����h��cuS�W&tv�Ic��6�r���ꁐזNh|�A�.���V�-]�E
���dN������ř�
��o(Zn�Ĕ�Kָ|�X-ԥg�:%{������h�Z��������RU�f$Ƕ��$��VE!�Z��ΰ��޺��[W��`	yQ�+�ť�9�.�ҬC�#g�q�9UE��r�F��e�7�"5[Hc^ۣi|��w�w�o�dHw�J�.�����b�U��>���zdm�)��Lt�6I���w��MI\�r�)�����EnL�I�~t]��KhI��]���e���=mߕ.7����qE��5�/��A,�M�c#!�����+��1db�Y��}oϙ$�ir%-���ȺF�g�R�d�^�X��4��%��j��[�2��J'��E� �ܔ3= hY��y��~Sh�v�D{496���e6�^�vN8�������d����R��-yF�{o!ç��ͪ��+P��ȍ�̓*�ҵ�*8�r:��.�N��H�i��6�'c�������h���gӪY��>l?��Ϫ�i���\�Ąb��b[/�<
Mj,������<����3w�~�����a�o�2峏6���F尫D���SM9�� ���q���zCɌ�E�#���t��r�*�q�6h�t��l.t��;V���h�L,���Ժ���
eC�3VHS�2�e�A�K7Y�l�z�'�$▭:\�t8C�$��"�r��YZ��O������vKB�*'Ȓok�|���j���a��i�ꦂ&�˔��C�ʁb!�l�,�(<CIpl�I��m�`�ض�H��v�q|��K��d��}�\�J�7:ɫ��B&���}D���S�4�;���ico9K:�V��J�l���<'�*X�ps�ۚ���w�I��&ɘ4;��Awj9�b:=���uP�>s�3���Q�;��d	�Akι�� #Q9+�:��\�g���T@B��F�ޓ*��B�_	+�*W��h�R̝���w,h�"�9,�q�e��gQ�s	C��v�AP~�m�?/疔���e��NVr��2[�{2B >�l�wFA� �7��e/Fk ��|�z9[�q����������:���Q�]p[�]�?�{����U\�_�}/j�U�6r���q��R�f�Rc�,�#��S��'�`ԺWM ���qSw��Q#ڸ�ޔ���12G�0nA�,���1�F��t#�c,�O�Af`%���d�Z�a��*h��J���?N����(2�%���C`"��ǂ��A�(d�1-�k�o��*Q��@<RJ�5����2c�E��aD~h. U)��U��N�
��.���O����f1�%]��C��=Z�в[��v�I��$Yk�4��n����bm�w:�U�B��f1�������a�8��xC�ߏ�	V��ٖ��9�bR��7��ra�1��0�kѪY�屧,[�+7���J�ܼ9�v�ބJb�9�װr�a�Z�,q݁�A�YQ�4' J�'ae�K!�J˱����K��(��#4�Xs�A`K��^U[�vtTN'�9�i��`����,��M�=@�[2[��)%�(M�,�n�*T���AW��ؔ� qd���hb]R�@�pJR۱�T/��хp��H���Cc�����a&e��"��5OĿ�mВ_�K�*]$�x�h.: ���:c�)6�K��PuU��?W;O���n�M\Vc�xI4�ڋ"bJ��f�Tʂ��U�^�0Q�V�|F|N*9?�9Y�0&}N���^7-W�C���R�Zr�/�/��������gg�����n'�V�N���O�+_�2����E��e\��qH���&+I��<��~�Lw*��Q���x).ҏ*��FLP�#�6^�i��1w���ܻ�@��1��ݫ�d����S����-�iK��4�^�OU���*l�w�=���/{��Cę
Ӓ���j���3��� j[�<Y��a��Y#u��뜅r@YHTz� Y{��G,�K^���J֨�-��ф�]	CHc�n?�۞(y�zt,�m�h�JYS�������.��H�5I��+}��_�x���f�cܲ\��W�/��W��QQ��V�3�7�2߯�,�uȏ�˙�"�}�ʥ�\�0�"?W�N%��*8�R���{��@�R'�����V1�<��mɸ@�.��h�K|��ǵF=kV�i}�y/�v�:s�N�b�oUMΩab��Ɇ�\�.Ӑ�=g�'#d�ܕ'��S�똊G)�(:�ne�]=���ȑc�n�{j�+�,��%�R���v.�o��C �qD-YJ@��u��I�Mq�y;;"UR�kQش�,X� ���^3X��}(l_���i
�����PY\�����N5�ԐJ����E��CX�u���r��zE��F���b4q�y�\��$�X�պ�śh���P}�'?����9���x�O�k���������/�*��&}]$Mo�DX�轕j�4ԥب���:l�K��]Ǐ�#~��|����	#�}��V+dn� �{%i�aZgb6W�4+���|��.1zq�rIP]+!NZ�ir-٫�h���l��R����Cd8}d�DՒ��?2�E�!��?k԰X���͠*B�.�����{� ���$$��������u&���z�ԉ�a�Ꮊ�i�A"mZ�^����J�-m"���Xيl�|R���C(��+3w�`8���J��-�
�uގ8��T �+�_�n�.1�~�h��3�T���+��}>]�qK�YJ�wb}$�2��Eʍ�%{���:tM��9u�WAz�GU�J�@I�,T��^A^�P]��-�J�L�+�QsRc�2fA��ɳ��9�|�f��s�dM�������HF)i�:mV�� S#�r���G�^.�dܩt$�FB� ���i$�Ž6�3B���Tz�_�Z�S�j��щ)򽤿���Q��T��<LZ< ���-%���0����Z�(be�q��i/�s9�(��Xʨ�u�S3 ���&cG%֪��}n��` �EP	2���%���Y�W<�3�g�Z=Wt[C9 �+P/1����m��w�=x�����ے�	=����<��|�կ��O!�ZF����u)�I|7K�G�SѲ!�x���N�y��jY�`��;R�7�]1M*�Uʁ5IPE(�N��2����^�o��H].��$F-/r�U�.B(e@��TTg�6f)z�@b+��`]�Q"���*.�����u�ЊF\�M���x�D�CF���R��PVm�l��*4G�{Ɏ�����<=�M�ǣ�@n��uL�f;��;J*X�nzq-���C�1�'j�E��w�v�����x��䚫�L��o�H�b����� w�+XU��ϟ�2{M�-F�FTմ=�����|+�^�q�&�g(Jb�t�Dʺ7�
�J.�rԎx��3�lu��5V�2���U�)�D�٢\,�}�'�,'h��C�3�!��3�f��B"���Rڎjx�n�l/�qWX�%Tu��ƽ6�[���ɂ\����i����F,��5�?d�
��~M��fz�,��(�;��K�,"2�����J���-���RA�����o �A��	��9潑-X�5�H�Ѧ������_&�Q�&���(�%"�=9v�NUVQ�ίT�؃�=���.(�AcI����N�µ�=S�ሢ�{I;r�4���+(6N�-syZ��j��cH�7��_�����6�W�=�p;�%�z���ϯ@����C�?�/���?��gC�|��ǆ�� 
����$@�����֮d�W6�>N4e���ׁQ��Xڧ��m�wy����$��..A;�j�f�`����ԗ�,�`��3D�����*����|
��$ӂ�_�7��SR����͚`WpP��Z��%V�3�CT�!m�-��@�XIR�t��И5k��HV�l�CqMN�IcW� ���hIqRQ]��%#�ѦCa��~p0��t(ܨ��%�d����IHl��Jb��t��Ԍs��E�2�{��PB�^�����\��Z�J�eܧ��L��]g�k
�7���0�F�������ⵃZ6����H#y-�$�8��Ϣ�d��K=4� Ւ�փ�e�t'7gn��� �0�9��K��5%&�Ui֒�~�	���19|ڗ������)ד�,�O��19�^u$����T����j�������^嘵v�:�6���E��	�=,���ZR�j�O�f�	�LT�C���Ʌ��a
o���> "��I�8�4KnJ�� ,��D@���|ǩ�3UO��q�G��fYy�dY����?��-���\���@5�6h��<�|%��cbŻ�F1m�7��vI|[��ڠ���ј��a���7ˇd �m�ۖ�Y|�y8^�w�}.����I�^jQ��HO���C�Ƣ>��?&�$ǉrE��=�荹���d��n7���D����`�.��h��t4�¶�*JҊ�b)�RwwaWq�	���I	'$��͏�Y��5g��T�����,�54H�Q{�S�N�U^_�c^�Ѭ�&�����3Z%<a��W2�tDx�;�噄N��TŁ��� C񺌖7e���V���	.�3��I�Ww�( D���d0Tx�U��� �*B��Ư��O-�0;|��]�d��m5%0�2w���q�P��!�g{���d�۾�mkC�w�ޞԘs�Lً�uk��F��6I;��Z���{b͉�����L9-e�"�n��HP�ӾZ���Ui��@�A�#���A88#V9�zck-�Ӊb�`��i�&͸&�ǀV�M���U�v6o�H줎X��������D�Ǜ��!-0/Tֽ��}���G	��-�m���j�35�$\RI�'
/� �6�l��x 7��v�B�9�aG���r�q�*J�8U�?a��3 xhL��@��A	m���P}`J�����X�)7�ph��qw�����XVc�>�J��_�\��e��be^�M޳h�ǦfoFl�ȑ�c���j��c��w(�^�f�����O}nWܶ�N�z����P���֟�ׯ���M�#A����EU7 Iz��%���Y�>ђ/�]i2�%�A� L0䱄l�v��k�6uф-b��64 ST�byۈ�8r��q&�;+Y�pbA�d.1�ʬi����c�f���$�O I���$�
����3H�-�zm������ɪR�z���3�*Q]��#��e�o��hw4�ɯDC.J"t"\��G��A��*����RAM%y�mwx.����h-�C��H�ڎ���p�~ 3_$�ɵ�h���j��!�۝�}��ys48�u�y�<>�|��3�D,,��NvKj9������
E�!�CY3]Iι�V=�<�i	�*REԵ�h�!Y�e-J���F��B�Z,`���A۱��B\f�myźi����Tޟ�J�z��2�%�H����� ���b�ɉ�3iX��QL�a3��\�O��'e��7({/G\^OϬY�Q=2Y�P����
!�\ͻ3�sȹ�p��DJ-�zɌ�G���˝�}j"e��j��=��{�ۭ��P2�%a���R=�$����/�+X"m�Ŵ[�I�9��b	�lR���;}w�+0z�FQV�h��M������cA����>�0>є$�Už����TR02W��p�H�5��|�z4W��r�B�.�D��oլ�/:$�\U˟�Cz�r��nw�քn���O3�߸�\���g��������!4?��Ie�S��#$Gc�<���9�b� �U�U�2m�-��!Z�n�ʈz���Y7����J2vp�;&Vݧ�c��ц"p��������~G�+'j�]1���A\���k�߭UI	�5Qc�Ԓ�s4��F-
���!n�v��V�����غbwk�b��+{���'P��.^��=�q],ީ�0��ȵ�+ֳ�ܐ�̍I�\7H�[��\Ԇ�h��.�0Z-Y�H.�Z=��s���`��jA�׀\�76'���X-8Y�d�w��U���%T��ג��sE@b����"-��Y�GgP9�a�e?�d�h@I���n�0�=6Z5�	�L<�5���ֹ���s�xr� ��:ƽ�
�j��O-�$|?���Ru2��C��FؤDp�ZK��
�J��l������ZA<<i}��׮f���^k8E�kU�wH��a�~�C�!/�hF�Bk�#�2ds��W�ְ�Gr����V��\�����Ӽ%S��D�y���I�,I���
g�:Vd���Ǧ��G�RP�]σAHq��O�q��'�-�V�m@{8�~$��C�A��-�r"p��̳0���kv�x�H~�"4��EA�KaHN��*S����*�n�TH>����LHk\=�&+��
���aYD�?�"?�'�j�0�2��]Q<���V��Gqm��\w(�i�������	<��!�	�#�@���g�����z���C�Z]���B��'��-����J&�����"n�G$��PmZ�.��`�m�\�<��S����jYVy.����r7�:���TTy;ZU\sJ�6j�H�s�� �vF�>)�UK�k �:r������l���H���G2'�Fk�}���9���X��Ζ��Zk�Ce�N�����oL�Wm���X;�B�AR�
��E��p������.��Ξ�g�(�q]47�b�~␥��NvN�oT���5s�k�ъ	h=-�^���.q$�6���E�B䤣�	$vj��F�v|�Z>xz]���^Q$��T�E��zy?z8��q�,��Q���e[�1����p�)F�R��Qq��~��ِ�k_�U>��t_�}�d������<��T�f���M���O
MF�A�"�E�t�%O��uK��-��r-�w^�>[�k�Q�q�k�G \��Xq���Zs��4����j��p�����S�9��%��W�R�{1w�ZH�hl'��&q7�hw�bFY�I��d��6n��^,4�Uh�u�%�tpB���Ǘý����!i�y;�%�����Xն/���|Ơ�"Q�[i����r>J��
�j[��Y�:��CDJ����l�C�|4����=U�%ᶳ|v��	W:i�f�QbŀY�0�H�玨S�Ԭ�gMA�Q�{Z%��C�a=b{!��G/ʤ�B��0sJ�kv:{���5؜��j���nu�9Y!RWr���]��l˟�o\���{o�'��?w
�B'<��O�+��[p��5��ۻ���_T!��!�3�.rS��I�[�Q�vu۳�*k��ˤ��n\M"�Q���z��c�C��E""-�,�m�V��e�ns���� h�%)U�M�� G��I��c��JL�W	�H��Įa�~Fb���fyJ�9r�#*�X2�7p� ��~�]���#�5J�.����]6�Y��D���c5�HDQ;�|wH�<�hN�(Ԯ�G���jl7��k��*�u�8���u8IC7p"`�y�(uӲʋ%~�~�3�U��9��<Z�QP���w&��A&�H�Y����Q��E4�A�Ȃ�e��(�"�����mW�t��G����l�Ӿ�4��%�dE�p^���t�0����7���AY}=�(�.D]�&�Fk0AVV��aZU0L	[���1�(�$��p�uv�C�l��5D�Vl״��PO��!-I��Z-�;�pDb�j�"*��rW���B�ˣ���2�Y��� ������#!$`�d&P�~5H.^'Zbʽ����Q�V����U]m�.Ħ���#�-���)��7��v��+۴��Ks_]�����JH��Lu�vx�jT�������TNH��j���zsX�sV���Ð�R�V��W�\.q?��=4�q1�:=�\�Kwy#����Q41q������ቅ�����9���k�.�-d��iv$��<��*fu�P�zr4���H٠�<��5^a�B%��h��F\*��(x�{�ʆ����Xvb��.�ZF)�g"���J�ь.{��g�Wb�V���Q��Q�X�bY�I|�+�BI|!^�f���,����1}�������ٳx�"t�C��,o�7��ē�_��O��V�O�e�yLÉė��Q��q��D+Oba|��Lgس�'km��PJ
��Z�Z-��>Z�&2o]�&��nQ�p�8$��e��]� vF+}�b��#�wx���-#J<�i��sſsc��<b�H� q/���%�Y����Z� '�v��AK����+�~R�e�[�����n�����W�p�����5\���/���2.�U$�׸G���]�X��B}[/:�h@7�Ӵn� R�p�\��U�w�C��v((��t�׳�;��.���>���������^v��� �n\l�M�����nׅaP7"+����!^c��~��u��w��Y��M����e�J��A'�U�S�H�BR[��s���a���FJ$h�C���z?Fϥ��xS��ɾ<���$Dݖ��&�
��޴=�yy�=�+.q��?A�B;$t��}�V�uw��D#��<`�/Ń�b�-l�lmqQ��X]8�;T���0��AJ���G]\v��h[�K$�x�kz��^�k��P�����2��w�ڽ�_߾�� �u�&$X�qs�r��'
���?h=�m���u^>�_H�[|�v���&S|��^��>8�͡AM�;�Dhq��M�Vx-*�^ց�N�~�q��H�UN;���5\�}� �����ݏ��}H�w�НG�=���p��Н41w�#��q)���%en�zt�ā�Ns��Z�T���z����:����{��w�No�c�Q�5I�,T�F	u}�D4�@�X�6�z���0� ��!�� �s������h�{R��n
�O妍O����js'��Z�|ܰ��(H���Ԩ��2��k�ѧ�iE��2G����-����x�?���7��y�ﵗ`��rG�9�#t-�~�wP��p�Ƶ�;8�s(L��������5�!"Yǎ����L�x&$Q_�@B9J�hr�es�I���d�����Zp��y�S3�\H���r\��[��	ʞl��O�to�X܊�FΐM%Q�c�<@�e�)���>�Qk���J�
��@?j�pnyG�#~7���Us�(��j9���oT�����[H�#���/���U<@["�����W]up�{�׿ԟ�A�Qfi�K�_3��?uir��iK�5�U�<X�Yۜl�dr+c��%���������ݠ �"4i�^���~l�K��\���~�#$�����n��l6��n 5���z�����1?�-���q�h":_��Q������M@	����|�1�
:����n��Dj���Mlɶ�f���py� .��.Ƹ���N��,[p���~�|�;�] �P����:U�m���&��v7(�#�B��琻���b�"j4����6������q�9Uזg�_Y\�pyu�~'��o�@}3ԋ�B�ڰ�ߣx�f�}Ŗy�4^�!���R1b;��_L�K�Hx�,]r'�����Ac�T�-c�Xi�m8����w�F�;��&�L�{AO.���UؑK`��:���Dq�ł׏�B��h�{Y����vp������\�w��߷�ۑQ�ˇ�Ck���=y��:�wᛞ�ϵ"�?���,��!Y���q�d̮ǟ��S�n��c����F���e`�@��<}���ND��a�{�q����[.��n��Jz���u��$<�Zb�[��l^'%s+k�����v������}WNy��W��/+�r;��V��Wi����Y�F��پ�󲺊���������=���O��w��HB'|�G���߅���~m;�����PX�d����Ń�ڡX޲�=R�&��(]��еW���K6�KLJL�=nM�y��ꂆPb�c��>b"l��*��)��ޟ:`��6�a���
�#�A@�l�d���[�*J)	�&�Y�4U�������A��H�0J�_��K�a�d~����g�:����VF��hӄ�JU-�@�~ַQqx5ٯ���Z���^����������HG���hli�~��m/]z��o�	��ٿ�����ݖ��+W�c?�ɗ�{�꿼z�$�a�D�ۊ\���=���:,ֹ:��!�� ���dǡ�Y�f��F	�A¡(o=�+5K�0>�+[��*�'��"IV��K0���4b�>����R��R�BIh�i�D�I��`$T�2��p�Bi�X��}�2O��b�\���d��B�H���ˉ�(u�'i$V4Gc�3�EB�#����;���v�:i�o��^Ajg�8�:���7^�]?��uj����Q
�uj���9o���~t,m9!Z�v/g넚�7p�#gҺ����vB�r��W�n���.�;6*���oO���z���owpR�~�a������Ο��G�k}/��9o���_Ev�P�n!+�t���aN�woK��q�\�DbC'������͐�7fb/�8
U2���w�d�G4j�G�J֕�E���Yy���%�4��/�p~���I�h��_F%j�ʰ�%)׭J'�`�K��?N>b2�ѧ�6��L�d��߬���@��+�t�R�g`s�;��	w,�z�3��W�
���`5|#�.~%\\���
��>4�^�?��8�Q����<�O$��Y�͙���'���2�lOg[Z��ru��%U����"�ٲҿ�	���F�����gPK�̽Ρ'���.o9�k�VC�5�T�E�	:��)�V�~�R# �Q(!d�u�H�+����� �����M�x}h���������U��.�on��-
��,W��/����?��
\{�X<|�¦�s�>?h�s�={_E�z����ۗ�f�u<g|�RF��e{��1��������֕����Cv�$��H!��Ą#I��=>A��k�xf�'j%�T�eXw`�&�Hڿ2T�I��Gz����m��%>ߴq�*�K��5͠�1��F-5�*�!*�\8�2��@zcw�M�7�|J�+�DCjC�6�ɐ6'h~o�t�z�h7�]}m�߻֋���$}���,shW�w#�k{p.��:}�����/����+��e��[�%��
�~x	"��;���������;o���Ґ�7��sz�܍js�2Z��'�6��u����G��?��~�nG�P����r��2��8ԱC��lJRd]��N|��4�r�* �I�t�����6��dH\���k��l*��ȵ�垄F�)_V��:���b����J+dU.UG�=��O���!X�t����K$��ߝ�KnO���m_&$�o���l뿎g�J�!Oȣ?�����;��	?��q�~#���W��r�8�%H7�L��O��~.��n�f-���dِ�HIEÄ�7�5�3��57�F$�U6�&Lc?'*�;&⹲֖�
%�!@Bo�^�c�t���I?�	l8Q�`����T�R���)n[hK�,R?�0�S��-�s�sp��\::8��^���ֿ�@|�^���f����=���܃�!/�5,P8����gΜ�����>��0�k�������j�.s~)��K���%�N�ڲW���TJ�n\`h�M*��U�'�Q�"HV6?��9.��a��!<�÷m��?��Ko|�k)�T���1�_�����.n��a�1<���~�$�\��uX,Z)���$���8�N|����u�Է�ݓ"JCZ:ɭ��J�c��IR@���Gi����q��km����3H�<�+E('�-e�e�����H>�(P^�^GfPJ���_+�#��i$Q�t�fGTy�8�8���"��b�:�T.7������t��>Ń~���쳴U�ͻ�����ڍ���t��:}	�"n�� id\�H��Y��u�41���btO">Y|����ӕ���!
��՗��jާZodͷ��fj�X7�ȷ${9�PʤB�2��ي:�5�*����w�"m{�!�Ԗ�X���$-O���s�5�Ggw���}$�g�����h��[��~��k/�CIM���
.�}8>Xܩ.@ǿ:�}���{~��Ǐ^����w��/��������'и�h���3�$�����Z-������D1$�b�b�Z?*\TRB@y,�X�r�k���ٚ���+�d��/�v)�L^+�8���<bd��h�`��`Wy��r��1h5J�<k�]F���,L|Z8�]z��?�FJ��f��|9�����Z��̣�l��yl\�;�"t�O=���<�?��|��+9�r����ٕ����>R��'q��萺�����4,�Щ�$��H	]\�b���&�b�2�hY�v�K�����3ژړ�T��5ר���j�r��~♭�ƭ�7{��ó8�x�")d������$C�tc�8��ษ��98���s~���K��w��/��ڷ��wp�O���1�;w��ӟ���������1ʧgК|��}����z���Ç�j�4��g}�m/V�_"�י�Y�Չf$SZ����X���)oП�2�M4`'�(\6f8LYf2����ÛF�s),E͠�w����DI��F9Zd����
���r���Bo�3וe���;d�kh��j����WQ���ܝ\�t�)��k�|
�Y:ᡇ�m,m��~�����{��p?�,����a{W�ǐ�?�W��H��"��C�z�O\DH�B�9Qt�i����Y�Kq2}|��5sR3�?��Y�U�mm=ZWK<;8�jNT�4�Hڌ�,t�~�עl�m7�*�s�,Z���耖,�1�%F��`}p��ѽ/�q���_;sp�6�o�&��;����p8���������y�m��}���s��j��'oý��O�����w�ǡ���L�|h�Ȣ��{�d-o�zhTlHy!֜u������B�y�|#�2�����[ו���9��N�0-����9j��t�Ci1�ڕc�A��$�)ɓ�Q�	ߏ2\���'U����_����0��LP����;ys�{N�zl~�l	�0uURS���z��2R�ej,������_�{C�°[��{���Cx���^܄тG�χ1!o���?�c������\*rB�9k���E)��[[�ɐ�=�h;�4��l����i_iz��[TR��N�� ����j��q��qLK�:����"�`��{��їV���}᥯\=\���K?��t�; ��'�����|�$��}�8��<t/T����rN'G9ԗ���c�2<����!�=(��#C@�-�|[�����]�=2��c	&��A�zγu��ReI��)�|�&"�[Ge��X�6�Mr�Ř 
06�	eh��:�UT��>�K&����->�?�5�
�ĺz�m|��R׿c�^W�Js��;��g�Mf�>�0�����Ԕ���K�C��}}��.�[H�oqV�嫰~���C�o��S���U��R�8��de�zu��zf��7�7�7��q�-mkf[���1�1p���)Y���#nY�֋o�bt}r'�m��]�!"�䦪B��h���n����i�r������4�����/_���g�y�_<��'O?���}�U���08�;��G��dI_y�۰���&��d�7��_|��?�{��Vi�[P#�&��������Q�܅�~�:,�a8LCZ#!���u��9СT�ID�Ȃ�
r�'9^8�$,iD�!C��F5�q%{��Y�Xq����ax�o��ȚjJ)��O��N��ŚH�*�N}
�B��F�����Fc�*�G�]l���K''�|��q_ ��ݯ�Ï���o��?�y�3��"�)��'���{��p8�=��V�M�"8f�m	��p8�9�	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8���o��<"�*}    IEND�B`�PK
     $s�[d��   �   /   images/d3b73945-fe79-451b-b309-b64aab767520.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     $s�[��RL  RL  /   images/f093df24-6efd-4d47-a863-17c5645b3aaa.png�PNG

   IHDR  �  �   ��ߊ   	pHYs  �  ��+  LIDATx���}�$w}��|����͌��F �%�!!�aa�`־[{msqwqq���ᇋ���%��?6�6�ݰ��q�F�= �H�f��a43�~�zȇ�}3�W��_gfUO�H��KQtUfVfV�П�=f� ��{:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:�s�������kk�V���L�8�?�t�n7��$�$	<��i�z���AN�i�i��F���Zi�$�,�iD��T�۵kW�̙3�{�7� �\ Ё�!O<�D�+�h���5^���|����˭���w,,,��t:���K{WWW���u._^]��eބz����J� ȼ,��,����Z���{*��4Ra�6MՒt��I�S_]���a�m�Z�;��δZ�����s��S�3�v�;��ҕ}������o��N��m�|��]��x�;vl��W_�������������������io�KZ�׵��}������M�q<��ل
�VE�0��N/T�H���*�*����Y�Ga�gY68��L^eYV�h5�2�K�12�H�EWm�B��Q�[m�k�Fs%j6&[�YU�?�љ?����{��z�[.]z�[޲t�7.z �:�8r�H�l��c�ĉ�ӧOO?~��O~�o_^Y~��ss�w��=*���z���FS�[�z>��5Tx�Bu6��S��4M�$�yi{��ċ��f]��,�T(��
h�rW�-����������q��f�Z]a����o��uUI��v�~��+�V���Ԏ3SSS�������|�e���ڵk媫�ZU��e�G���s_r�%Ӈ�>s�̾O��o�=7�����۝�>U�ާ"�
�iU�PAۜ���[�V���*�����a,��,��		ky�r������ײ�\��������A�/TǕGK=v���j�:����bgaa��N�<����#���q.lD�&'Z������������yU��x ��l���?�������C_{��gߵ����n�sy��=�6�VA8�~J(6U�;_�Q�����PGQ��E�`��:�=i4� 6�@�?�t���m��m�z������^�o}�(
������b�̓Ϡ�5�Ӧ:�i�����:��Ͳ���l}hv����>t��h��{��g>�'�x��^����n^���;�mt`T���x�{_}�ս����'��������+T��k��;�$��&n]�֥o]
VA��,�%_��,Yr�������S�\�W�{�s����\��[_L蒼�90���+���4�[�v{��|W��7u���S�N�w����|��C�NL������w����S��~�Z� �78?���+��r���_����N������ޔf�ժD{ M���nwR�0�B�T����[�SWk����z	N�z��/�f�jz�f��ܼx��1��/̋	��܇Y}o~V��'�
��^�򪵵���kk�;77�/~�ԓ/�����X��u��2���]5O�y`�t`�����z���_������F�X�ߢ�|F��Taˈ0i7�f�m���z�Ts���~����ҹ��,��c��(;O�t_�9�����T?�j�n���N���^;u��g�{���~r�e��3���/��s��K�/x �B�c�җ����矿�S��ԯ����ވ���`�����Hg1�6ץ�ͨ
d{�ӛ��|oY8s�����û���e����$���'h4�{�˫��޹����W^=��������ƭw�u�W�����Z:P�����#�\�������t�	�覉V�,KvJ8I��m�:��y�������
qs;���i�eǳ�S�O����P���:^o�l6��I}��MK�C=�K��V���u���Ͻ����w��?��}w���{�9]L��F�%~���������?�K�<w�z�*�_��z�h�u���l�mY/Ǩ�p�̼h0k�ڿ���j �R��ެ	0z�ʎ�����>��Y����>j�t��h���z��z�-O=����{���{����/?�����}�0�@�j~��߿�o��?�ĉ�l�������K�w��_�h'�ҥ�>&��;���eʪυ]-��a�{�WU�WU�ۡ^u�fo���S�ň��^�cǎ�EJ�YR㻓cKg�f�9��ޥ����sw}��c��ğ��]��{���~7U�@�����W|�3��#/��k���wOLM^��|�Ĥ��j�A�$���8S%I���2{��Ϫv���ef�\���|�qmf/��P/;�8���0��=��b)j�/ �"=�/M%��F��E��N�s��O>��#/~�S���_��}�9�d5 �x�=����>�����_����݈�k[3I�x���`����Lc�7gk���ǀ�u�xviVO(��/t���-{^��>�ݮ]�ٮ�B��u*�z�y�����w)??ʗ�w�/��+++�z�_-���?w̓=��S����#�<���q9�/�˗}����3�>���v��V�q�
?M�ي�q�E(�z�)Xu�7�f'0sv����v�1}\}��/*��5ǂ�G3�c.7��Mem����m�e�vU��rL=&_���ˋ�����)%x���q:�^_��C����ĉW�O�����{��
c�q�"�q����?×���}nv�WVWW��q�<�����Y=]�.	vs�7s�z�e�W���9/��7R�/6[j6�g����W��}��bng����f��;��ּ�Q��=�N睯�9si�{��mya�O~���}׻�=�"C�����~��o~�[���k��Ue߫͢W[�t�J�znt�K��T��z}�����������<���lg�7����ו���V�,�������z��C�z��ceuI��V���/��<�ē�--,|���z����i��踨�=ȿ��#���?~�_��;wO�.�01�,&!���PP�U�z̹��<|��^�u%c{����#�^_vsU%~�|ƭ��zǛ�q�J_z�?�ϯX��s�vv���a���џΤq��������\$t\4T��g�?x���s~~���.��1��u�Hov���X��?u��l۶{�[�S[�����Nj��QVk`�7�e?�F��^7�#w�+���韫���u�q���.� ѝ���N���'ON}�ۏ�x��O�ʯ�{�.:.����ny���s��ݣ�3l��n�
6���*s��\�;��}���BϜ �JU�{��ks٨��	����Û�}�sn;
zC?��+��F���?2�P^�D5*ԛ����_�x>|�����~��?��#�qQx�����_�׳�gߧB��#]J���~� �wB�S��R����Ӳ\�K����d>ь�[-�>===8=��,����e����\�fn���}�ەmSVCPVBץn���dN�Zv\�������Is��~��v;�G�~��(Z]]��_��f#\{衇>C�:\G��y���7������>�x�����`6��l㕐�	�bv8o0w���,�u2ۙ<$\�d(:d���������� ��X��voQu�Ӻ��mS�Uc嫶���1t����.ɗ��,����.�J��C~��,ߩ�G~�&9ҹQ]Pi|��c��g��?�я�p�m��x��t8�{�;2�ȣ_����'��
۫�T*qC��V%��σ¬6kkk޹s缅�O��� �0�a!��]�釐��s3�eKKyo�|?�عsg~ ���<ץz30�ڝ�@�O�:x�y��'�џK���yOOܢo�"�|ֶ(*�����f�KY���Z�������mc��|�~��z�����U�+Ȇ���8�|��f�7?�ʿ|��K�?��"�ᴗ^z��������47�^���ٳA...z���y����K�v�Z��b�)��տ�:^.�)��%���o����z�N_ }��:�ف�k�-YOJ��� }�!ǔ��iAj�I�ں�g���J}��/�=�mS׿`p�Q�=.I{^���X\X�����k�>�虻���8�@���z��>�͏--.ܪ��B�P2ȑ�����q	h]Bסm2��uۺYR�%�ݻwB\B]W�����ݛoc]U�z�Ym.� �	f��0��钫ty���ϩ/*����̟���ݸ����dW�^��uA���ߊ�Ԡ'�Y]]9��+/dzz��O<�ķn����a�#t8��ї�����W���<���os��I?��;�I�I��Ozf�Nm��b�lP2�a���幄��V����R����	󩩩A�Լ�Ъڣe��/����l^��;��9hf󶯯��z~�={�x���˃]�ؓ��7�啱;���5�d`~�QC��jR�־�*.ڊ�e��	�����+/�����~A�~�C��I�����t����A��]�jׁbvJ3Z��� 7�gס�K��St�Vw���PzzX�!N�Ζ��������GYxM�9}�t��NJ������x�S�n?��R��s��+򋎲��=���!N��l;�}�v��싀�k��Q�8�z~�س������E��U_�Z ��p�
�����z�Z���,E�CW���L���XC�a�K�z�����r==��&U�C�.�� ��m�,���/4�����R*?{�����/^����5��t/��t�^���	N_?/�_�����T7��f.6�9��W�o����N���?��w��p�'-,,�\[]��z�f)ۮz���r��s�����rI"�U��7v��Gs�y�.y��C?�hW��.ƴ�achJY=�L��9�'x�\���Mu���8\M��{�yEQ3?�_+B=�o�CW����'�/t�v��]�j�׮Z�nc�Z^���ř�ַ��Wu��������^Թ����	�@�ct8iu��CEь
�PW�={� ��p�:\�2K|�R��U�fș��*z��\�����z)K�\w�~�p�nfff0[��޼({�nz��m�t.�$�7���s3ü���8��m����Ͽq�|������9��������D�߷��8��!��$UBW��<-��[z��q,�W9� 0K�e�t؛��CQw��6h�ä��-���}̺[�jRe��W{gΜ����y��l�6;ەuJ� ��t����iB_����y�u`+��n/��nw����J��j�s/~ͨ�,-O�Ξhx�ct8�ш�8IݎlN�2|'�d�}f��d�Io/ᧇ�	�'���l�e����vG�:zr)�K�y=����f�KX��={v�a.%}}�2�0ѽ��q�湛������o�/g^�=�Y�^��#�/dt�}�K\]���"��43���fI[�e�f��:��U	���f�4s�Y���U�2�g�q�r\O.,�,�lV��;��Y�Z�F^�/���>Ϫ��^u~v��k/����C��Q���m�y�u�<��xȶ��EE;����pR+;�~,%3��&��U��f��y!`�Y���u�tU)\?��d�]@�*��6~���\J��g�ǰ�)�߶<T�7�F��g~'��MU����{�wQ�㜃0��e��v��O��!��$jq��HVW�7T�c̽���e�Q����,����Qð6S2�t'>�֡���ef�����3{������Qm�em�z�f�>~U��f�2\�o��;���tv�Mf��st8�՚H'[����biI׾�IY����X�l�����<ި�e&{;s�u�3ꐮ��^���P��U}��{ٶU�1/��k����}�}^{��w������\�$I693��'��C��ISSS�Ԏ�����g@3ǡ�{�m��s<vYռ9{�]��;���e����m�J�v�u�s����o�t?܉l�tm���e�e秷��g��¢�v �9���M ��[�^�Lϴ'&&hC�st8I&;kM�s�����Rm1C��N_�µ��m�q7��3n W��y[T;�˖��/�[��u��_v��6����� .����g~�����X����.0�9�['�&�i��p�'%I�޵�_�_���^���a���iY#V�$�Bc�hUU�e������jC���c�풪��*���l����ظ�TE�{�?�g�����?�V=mzQ�m���>�^��Ȩ0g����Q�
'��.�%o
|/f[�z��	���'�ɞy��C�u��p<������M��ћ��$���j�?�j/��ס6��/`���y��Ԭ�ׯ���OBf��2���J�)���m]M�ݴPwnum�v�z��T�G];��<Ɇߓ޳>P�����ȿu����U��)�ʢ��d��<�W;�C�T]2���S�ykT[���k������s�'2��
F�yY��f�����a�nc�ۖW���wC�W��٧����w-�^L�SL�#��$ԩr��t8I
�Y�������%�Y�-�&U���X�J7ãl�Qs�9���nm����U�Wu�{^���Iy-Cչ�Ǫۧ~nN_[�}U�A�yV_TX�z�������@WxrŶ~�x�!:����_��>=��k��z+����q���g�>�f��C[�w%���mlf�W�@�J�e�<N�Q�m���ܟ٩N/���/ۦ�V��}>�7__L�oP#w��o�in%��$զY3����!��$��S������LhI�h�ց�o!j�
7��U�8���˪�u-����6m�8C�6"��J���q��� /kv�{���ng����u�{݈����^�[�¶�V~����ɿ	�N"�᬴��[W�K���
�P�i�4ﰦ@��%������0z��xY��0�c��n�7Յv3��:���൫�͉g�Ϋ���47�g�*��j�������۟b��y�>կ������E	�P�p�'��܍�a������Ef~:����3��f�i�J�uA[V�����xu������vv�z�~�:����<e��2�C蒸<:�n1��?�P���7��U�zX���P�Ԏvz�kt8I"\�叿�a��:y`�v	�|L��L~��,������
�8�����J��n^������]|�����~���\n_��~�}xTi�|��1�7��n�7�c�w���F2U�oC79��mWe5�~������g�bŲ���j4���w���Akb}�8�O����.�u��q�:Dt�MJ�z���K[B@�u5�پ��Y�!�̇9�[Y;�8%ٺR��9���4�[w[U/�����h޼�������>��w�7A:��/~O��;��;>��a}���N�d�����~ճ�����e�����]�[^B]C�����PU˫�j�.[�v;yɴ�#{�W����|����1�k������|��#�9�P�Ό2C\>��k��zcJ����C:\��Ü�Y%��E���rC	t]�U�:�%�V�����t+c�ʫ�ū^۟�j���4��}��S6n���8��ì�/�Qѿ���%si;7����@���C���E:.
�R��,��0J��5$�ԨK�L��%�Z�Aojs�y����0+_?��<���ju��[�������i��W���Fn^T�5��9�}�u�G�8="A?�u�������|�߆�`����pVY�	��זu�wt>V�_2�!���{Wײ�,dz�w]�/cmϾ=�>O3��f]3�k~F�g]	�V�f��2e3╅�� ���F���n�9���n�~�}�߭}�;��_:JN��p�'坞2o�jU�]�+���W���ɫ��ޠD���g&ӓ���m�u�������m�e�1_Wu\նnԁ.I�M��f���߿n7g�z���?>�����@��Zkkk:�C��Ii�S*0������.�m�Y�t��f~'����R�������.a�2�{�W��y>v	�*����.�b��.���f�u�9��	}�c�����t�C�{��~nf�:��5��6g\(�ȇ(����p�����4�#U���p��5�r7C@T��%F=�Z�IwZBo�{fO4[���v�f���ߊ����2K�2�:�՝������x$I�Kݪ|;x^ƜD�j�y�3YY{�ݛ~��Y���F:���~��Y�s�=a�u}�T��M//�����gC/�ׂ�C�y�%�}?Lӵ��� ��$�'����߷�fn���p��)�mn'��t 钻9�JB�<�ّKLN���?�ݬ�th�������6�j�n�s���!o���g3C�^&�1ü����d�3kE��Uu�2��a�{Y��L�s�@���4ieY���i���׺*W�r7�[��'.�׋��0+J��P�T��ץRU��<I��z��Jٶz}�o����M��N�E�nZ0{���2���u��"k��[V<��D����|�1Y��S�"�Q������ovP�n�y�k1�D؋;�烱�f�}��K}t'�4�{��D�K��� ���yu�_^ʵK���t ��<�,q�jV��cٝ�R���yT���0����(����}����z=J�p�W�R�U�Z>U%PaO(c�z�n.b>�x�^c�����뒲�6���uS����C�> ����U5�v�쳙�/���um��q�Σ�	��Ϊ�@/+��}�Y&]&�X�!��@�ҽ���.v�T��.+�;�t@���b�K���������1��Y��!a�zG���p{&6;l��(;O]��۵�>�}�dv�3_��,���J����U�-�=��N��9:����/���벟e��"Pҡe�D1�qs���m)���>N�.H�y����?"/���w�Ҽu���c���a��7����������]m_4r���o����`�b��>+>y�O�8�~O���lx��.A��J�9��R"b�!��$�G�5�Y�T��O�z{Y��A^�-�6��-E��}��*��Rh�[VV�.U�uwd�;�Y��������M��uh3?�]�7���)[Wv<�=e��?�$`:�C��I�4	�(����dNR��=���6_�w�
�����{������g�6�$-J��nYQ<5��Vv���.���l���wT�V>�9J��P��Ual��.on'/�^��=؍&����2�!��"U<�N����~T�p��R�Vj~����J˛=���j��_�166A���n�p���%|)�AB	�!��$?�>����߅����s�}���+EN�(W���K�1����jtH�n��}��g��>�n�8������n�F���*��]\�P��z΃=u9m�Hg�T%��T��s/k����x�)�PUPW�_UB�:����i��k���}p���"�ݮ��ن���7�T>���\]����i���M�i{�z����c�3�]����G�;�C��E��ݷxe���B�|.��/C�|��~~U�u�ƫ���v���q���[s�u!Qv,��K�x@�MB��9�I,�^XVB�S��r���}#J��÷t���w��������6N[��0���`]p���ZXu���2��9�Cw�oS�tS�c��@�s�G=?�FU��ެ�v{H�`��]J�U��s��Н��}WQ��W���K����I)��"A��9ǃ^7�0��q�B�E�ǥˍI�dh��*�+f/��U�ö����iQ�^�_B]B?��3#�_���Ƥg�c͘�ǁ�c�������1��1���]�
v���X����A�P���������� �3]P���O\Ŀj8'C_u0N	}��:��
����u7x}��Z�ý���8�����V;�](�j�����a���o��?j8'����GI��cYY�����o�{�{�cJ��Y�ު6����Z��n�X]���`�N�:5����ajz�?������t�z�ױ8�@����v��_���uPY"��K�v��3^�{�������ɬm�h��	��U������o!\[��z�����p��׵^�V�����B��>U�K])�.��Uӗ���j2��c��$����>G3Х��a�$�F��|���mD��9g�#I�ָ����*�:����wv����6m�ㄵ��F�kX?���r��V��k���@�St���iƽd��Ӆ��[��l�Wm�/ަ�\54���ٽ�G����gܡ�r��uҨo���7��E����,����笭�I7�5x�0�Lh��P�6��Y�-k/�0(s;��}���noW��jf�LBq��WO^c�RdoF�#����D�l�:^�tjf8��溺�+���ڙg����^ƓۡY�k�l6ϧ�4n.�:�����;ם��q�>{��ap����+AW�*�mk�6O��nfX�߅����۱c�>':��9:��X��S�ڡg�v]){T'����� �L/w=�NU�}PqS:��_�z�lWUU^������m�?�u$ц��pN���8��?�U�6��{t��i�MTF%FY;qq��������Bw��]E_��[{��"��f����o�Uϳk3��!��Ή:aЍ���?�ڕ���oD'������nU;��}{�%\3�SkJX���}�~���f�׾H��A0z��9���*w��@�sz�n�&is;Jav�U] lf_���9ŪP�K�fsU� ]�^W�m??���sd�����<?˸e�C��9i�Di�5���*󪒧ݩL/+���C�n�V�qIU����
�q��B�Po�;,k���EUII�@�st8g�kK�z�8�4\���3��:ם����1W��5��n��n�Y�����};.�~e;�cT�����?�Y^��7�Z����e���aT�E��lU�7����U��7s�� �ϣl�fj=Fu���g�}�+�8�@�sf���V����d�5�����}�=/��c�?��m�v�ږmƈ��+�#;����T���O{�Z�{������o&�떗u�+[6h���c�[=��r�;Y"?e��f���k�'�C��t8'��bU�j���ó���o���������U�U����~�����n�:�Q�s��_�!��V���ܟe�vR3��ڥ�J�S����ۮF.[VW5=�٠�������l�}+�c�_��?��3��9B��9�I��u�SI��U=�A�՗4�v�^��k�zU�\WB�k�Q�޶.��:�������7���x���"Ή�8���ۣ�8U�KWm7v�M��}�u�Q����*ԫj%�>S�g����ۼ1n绺����H�ڵ�D��I��F��NkV������ێvk��_]s�8��}�ǩ���of?e��>?K�*w��@���,���Sܸ8*,�J�췪��r�~ͺ��nf�-㢧,�G��@�L@�q��~��߄��QJ�[t8I�D���C���B5��6���Ԭ��=��<���,�WU����F����6e���/y�Fc��kp
�����2Ը��l���*.�b/[^V%=n)u����o�^�*����n~^}��S0���[�z����a����F~��_ϲhq�*w��@�s�N c�T���*Z��L�v������l�Q!汪�����j?�7�;�f#��j��ϒ$��yn!��5��*�Ū�+��Fݶv'8s����,VY5��>��ZW%^v>U��v�qFͫl3�ovgr���ߣ���=�%=&s�st8'��t���?��8ۏӛ�j��v7�6�q�n{�6��v�����R����#���ԍ��p�JqU ��0�GmkWKۏ����4��q�ᅮ]��g>�lS����U��EJ�R��oK�4�����d�B��9W�޽:15qxmumM��5j���k�>_ea^W`^P���ou�V�W���f1����gn��=/�v�e+�ι馛�����?������e�����Gm��*������mʪ�͠�S��߻��~]U_7�m��l{�d���ȗ���Z[����� ��p����W۝�[��^M)}hL���lhօhK���0{��\�u�����M�B��|��뎿*��G�z	��h~��z2����gfff�<�1:�tٮ�����#�p���w�?��j5�n����<�q'�?v�-��73��T��Z�=�7�G�/Қ`'4��Λ�� �y������7����=�n]v�`��1�i�u�m&7:W��$�~�aC�GJ窔6Vgg��������~���=�1:�t�~������g_�z���{��zؒ&��SYi��f�'۽��sU�P�)p�ޚ<ޮڋ�Ie�4Ο�o慏<VW���Ԕt�K���������;^� �p�}��w�|�S���O^����˓S������?�;v���y�ũK�{y��wY�v��I������7�����m��������D*u��_g���n���̮o�z�ۿu�o�� �p�/�rˋ�O���ǎ��_����TImJ�R�ڍ��voDǯQ�3��Q�������٪�����}�z��PFJ�kkk��q�;w�q��/��W=�Q:�v������o�8����G/i�&ޡ��7󹽷�ڽ.�֗yo
�<.��yq�=ݷJn#g��r��`PZׁ��z���k��������ʿp���s�=�����^;s溹��I�G�`��jlWzU��<،eoFI��M���+ǩ��w�Ʃa(:#�T���̶۝��-W}������Ep�����>���������������ٳ����ĵ��˓�ovu�8��īT�r��GU��xS�W�Wz�K�������BM�ə(j~��W~�����q洛�y:.���p�����?���}ciye�Q�����ne�U3�����6���d���u=˫�_(�a�z���J�����;Q���]w�����=�<�"@���[��['��կ��c�}����_�${�ӹLB�
�b\z1J�D�ݹb�|�]ֺz7N^2,��F�{���כT7\�r}~v�@��7��k)A����7�쒻���C~7B��(
��2�[�=�q��n��`5I��&���r�ͷ�����#�,y�E�@�E����x�G����^��w��?%I������]�Qnmm-���	O�}>i�,��V�Id�,�����e-�fV�޲s���X?^/z�f:���-�GQ��JF)�H~?r���8������}���=w|�w�w��cs�T\Tt\����_������o}�{�=r�����v�T�!��P���.��=�u&�\f�eUښ��}CU�gͼVtu�����6κ��{�{ǻ�h3�K�cd�|�rQeV�����f��n����G���������ɏ��������y�ņ@�E�c���C�=�կ>|����?�V�~��l^�J��%4$Lt[��iNBEJ������y>���a�.���1�{�֗����w�y��$%ty�woԔ����� 🙘�|��w��������P[��������7���������W�������*8ߪB��*�O��J���*g�br��"�Ǩ�.k��+a���^�u��H���di���DչI���0�^�{��ϥi�S�;��m������sױ_��_?�o���z�Ō@���~�ȑ�����w���[\Z��n�sK�f�T�L�%uy^�d��Y7�jU�������P�����|�9V����}�]xLOO{�v[�n͢(ZPT'���n�ᆿ�����w~�wN��/�����o�/>��O=��|���?�����+�Api�ј� ד��,1�+>��}��ᠴ{�W�j��U�^V�-�^�����>�3�a�k-꿀���l��=�|?xmyy��k��������w���w�~���= (q���ۋ����<������w�:�ꉏ�q|����U�H繡<��3�����T�U�7�>U�fvU�u�{�~�ھn�q��G���i�{�Pe/���Ν;Nu:�^rɾ��k���?���?|����m�:P�߾��<>�ٿ{��'���_<����[TZ]�f���f��y�{i�zaP�n��>���=(U�rG�~�m�*i��KӢ��ш�Ҹ>+����?SQ��s�g^q+S�N��@3�?��=��C�F�����W�)P�K�vA� dy�܏\:A�D���ey���8~ٯ,�l�!�+q���hM�1����~��}���v�:����{�[�1:0&�iN�8���=������Շ?��s�f�Z\�G��\јh4Z����u����U���B_��{��|+Řv�lz���ev�3o*�u�~��4K��������r��BBj$�嶢�,׭�r�Qצn��7�:����v�c􋋁�����I7���7ő�2J@>r���k���={��}��{���=w��ڭ��z���?� �F�����}F�8s�ȑg�|�k�}����г����*����v7/���4�li��-3�I��>��R�zg;݋�n���4袹<��;,*���x�sʗ�r
~�3)�����7�G߼����Q��:�C�Q^ji��?�u�@:�u�ͩ����w�ջ��n�~l���~�~���8x��O^<���:s��.�y�[f2~�%ռ�4�j	4	}�3�.��Z�r1�N����½h���ot)�+J�z��n���שg�lŪ��&]e��]���D��ЋuM�y�$�&��W����[[��:33;�e7�tӑ_����/����= �@���n[y�С�o�����s{Μ}�u䅣�s�Νm�'VVV��V&�W�w���L���T��z�*`76����w2��T�kK��7$��y(�IU�*�#뇻�%`����~����ӽA;�9�����p�`Pj/^��EI�η�.�'{I� ˒ �:�3�6�����PF	4���5�\�]y��ށ������=� ́�!Ёm�������ۿߕ��۳c���������z�T��?~z�ɓ�/=q����O�v��������4Nw�i�����P�9�v�R%[U�UڏT���O�f��G�)-�!L]��C������Л7o�?���j]"�(
cuы��'qG��Ν;v�^�������}/_y�UG���K/ݧR?���[�M��>��O}7����q����6�lEo����+3�����v�={��j�Zs�_��^�G�d���ɕ'�T��������������/_XX����z�Z�����M��ܭJ����۩WJ�SI�����L�%�U��ϲ�/�ȇz�^��uM��Ey��4oF��Fo���|ԩ
�D=�4M�Q���z�N'Q�Z�h�vL�\hM4�,X��5yz��'ffv�����������k��bi׮]k�\rI��K/����������굓����}2
�5�S�������:t����v��W�a��TS�n4�ׅRGm��F_�屡z�رc���-y���E���拇ʹ�xoG|�ӛYYY>���|e/�'	x?h�AI��
�@����@oPtf���m�;TRG����T��Ժ%��륙ڕ��˂�*���M�ԵZ7����;�v̪t����;'^qp���n�i��ɩ�����
�v�OA��k���.@�F���L�h0O�:�=j�[�/= ز={�D��7�^k7�(���lMD�}c�LZ��?aJ�)�����V�
U�?�Z��4I�ιsa�q��z=_]H�Q���Q��	Μ97���MLL�vRr�/���;��
�$�Չ�)��*\cu!��ϕ�߿?��>�ٶ�Uo�f����{���	?����A��= �@�(I��^��(���1�����wE�h�Zt|;�ӟXe�����.T�?�V-�ߩ���j�y?��� ������*j��ݯFN=n���R����=��4(�������F�[�q��ɲz�^�Cʔ5)�{ȥi��~�VAދ�f1$/-��z��تkU���~�����˄-~1����SN7Aڈ�D����y?
�v7�K7�� j���,�q��0�F�wa�C]޽��ĹO�УL"<���y��Q�֖�w����[��lQx*����*q�2���{�~�ÀL�d�Aa��mr�9��"Ё� Ё-���zdQ�rC�<���gb���b'�ߥ��P!f��]���ɳ�Y��*��X�kR/jE�P�$�{�,��W�y�OF�0�\��FV�ԛ� ��z($Ё- Ё-�^�~��L����N� �Nrmϧ�W_>K���i�"�,zU|o�>��:�ER��RUo��|�, �J�����H�~����@�HơY��i�M4�[��I櫜��O5r�
pp.My��;��b��Q�l�l��̀�����5t�m������U���-�2���s�`V���
)�[C�[t�7�?��sk�,���A���,�Gk&�R�C��<��;j�������^|��ٰ��O�$�t��=?hqz�e��>?�<Hӄ�ܽt�@��@��Ts�\;Z\���q�
�a�J°�!Wvm��8���G���D���y#Ёm�B���v;I/ɢP�m^/��v����������O�=M����K{ъ�B	��� �@�*Udjr]��b�$)��x�^ѹ���w��Ǳ�4ll�m�DI�dYҐ9�e4�]β(��������|�����>`�\`�t`DI$7b��3^��m���%�?!}��\�9ܳ�o��y�O��{i&��~��y�-!Ёm�l&I�(������qdy���_�a��*5�~C.p��jy~Kw�_	`+t`�i+Q��n~C�^QM�8T�P���_�O�>�-+�t�$\� l�l�D��T�í�(M�*f���k^�QpГ]W�K߸,���l�l�b4����/5����K[�GX��+	�T/�@ς �� �<�R>o�Z=I����8^���V��*:z�(�(SS�����jrW:�.Ͻ���թt*� �7���8��e]�4����͆J����ξ=D?+�o��]^��=?����p�t`̤3�Bv�����Q�o�*w��,����+����ߟ@�<��H��ďO���x ��lU��|�O{i�7����$ɲ����7��q����O�O0#U�A�)�/���H�[@��@�н�Sy���Aѱ]��7x�n�����l��m?ͦ�����m���7O{ ��@��ҥKq0לO�n,A.�^���*�w�T&�o߾αW^9ҋ��a�O�7��{Ǣ��`�:�E:�n�n�=:����^7�:����td[z3����w�=��N��x#�≉�j����T���믿~��%:��fk��~U%�b�׻���zk�n7˲�ZM;z_��y!���Lοx�љ�駯��Y����6��T'��̻\=�Q�K��u	{��o�Y��}����{ ��l����WT	�ө�uZ�
u/x�oL�������K�ی@��W\�z�ر�MƓO��3���r��Ox � Ёmt��Ai3?���@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�@ �:   � p � �t  @� �   �  8�����%_x\�    IEND�B`�PK
     $s�[2)h�V
  V
  /   images/72f663bc-d85e-4d27-9085-2f4219a623d3.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��+  
IDATx��{pTg��}�n���	6$�b��+��_�Hg�qԡ��mi�S�L��R�h)"��2V*4>�S�MK���S^�-m�1P$aw�;��s�ݻ��������w��{�o�s���� a��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0���~�6ml۶:Ν���0-�up��AeU%��� K�>
��)S&Ík!�?��=�qg>p~��ضc+tuw�[G�O�x�%�U�(��!�Lo��L�S�߼v����,��X/���>�0L�0��RH[[l޼�m������K0i���L�lTU�����Ϝ=�w��n��$DU��欙�4]�PQ�c��kh����g�LUTV����,\|w>Lnjn��q���ǟ�ښZx�W����pE�������X��ul��<��+���SgZ�%|^FU��'��)//�g�u�Л��:�6xj��a��M�زe�	VB��	{�_��á������wE��w��B��8��CH���m��t����^�[��h�N�e�߫���]�X=����W���n�GY\`%��_߂,��`pt���^���,�.	2� ��{�D�V�:+LAy	,w\k����3b�M������?x���+!�550n��`K�kͦ�n��A*�#����c�EUWW���O?$�IԲ�2�u}PpEF�a�:6�6��d>���fBc��HOOgK˟���tvvB4�j:��� 1
!��2��
���>���n!��?NH��[��
9$/������`4�Iyy��JH"�Ŀ�����Ax�B�t�J�ES\�8���<B�|�!0��Hq ﯋]�@,.�
�0�a��Jd�x6��\��iT�=�5�s]�ؗ�5L����	u���.�2|����4.\���u�>��@~fU����	�
���[z�{�4QF�Fֹػ@(.��d�%����/ �H|��0�>�p]n�[,�(NK��4z��X��UʃA�(�$ܓ�6B(�+�\M�f5;c&���x.wuc�V�,�h�(G��HQ����"4jH��L�a�`���D�mۂh,\`#�p�(��X4T��mB*����8���kΠT�Jͦ��T����
/���TQKr�=��?�D��K��Κ�N.��H�{>�'��t1��[`�u鴅�~K\�b�W1�:�Ғ�=�j�
�MQų��	L%��6Bz�-/��A=���'���bL��������0h��ˎ���G���M(p���t�
vݘ�]Ǡ�i�f0`%CK5tF�v.��fY�{�EZ)YVq�M�>G�?��%�.�M��
,���E.�v(�s����$��Y��4��4��CE=�������;��:.�7�-]�ua�Wͥ+77Z@���K�#�U,˼�t�z�F�B���}�﬽U���2���
��B�N�s�4��8:��J/�FVo�<;�-�n#�=G~T�q ����M�t�����K�����_O�I'S8mUIH�;�(P���oF�����ׯ�)\.�G���k�\`#$�Aǂ�13-�k/�N�ϔD��_4��y�?�1�=�I
��?��e�Ce�6BLS������8\[S�ö�{��?8�q�*��[^�*�����Ϯ[���+V�r5�a���c��ѣGZw�ȳ�Tz=v�cr����4卐�R\ĳբ�A3/����?�ŋ���r���p���.�BlX�.Zw��h;s�Պ�ʿ`�� NM�Vj�X�����(�⬐���^C�ͲM��}�4M�3�,�|<�ױx�#�EaƜ9�i�F�+!�����e��ɓ����US6~��i/�nrߩ�g.uwE�c68�[���4T04��(�8�͠���Q<�qUMe��o�ؤj�WZ���;�	o���.�=�w����7��{�O������So��=x���k�n��j����N�c�]kg�e�EB����8�M��ب[n�����V�������7�k߀��m��{�¬Y��#,�xl޼��������c����>��eۮ��IwY��E��b�^�O)bi>����XCǿ���E#Q?�6?۹Cl\a-�� :&8�O7�e��a���ߥ��׬���+��oD�Qx�����|vl����H�T�CYwRrK0���O� �fu-����7��5njƲ첡,��T�A!��"�`/�jC��It`+����$.��`ِ�~���J��k�v|`d�S��ʧ<�LQ���k�Zj�{!i+�`,G]���~�C_�bO���>�C�� �/�"P��y0t5-����勗K^O�:��^��ѣ��{oa/��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0C
a��)�R3�fH!̐B�!�0��}jS�R��    IEND�B`�PK
     $s�[
�8b  8b  /   images/a7e3301e-fb46-458d-916f-a05c0bde95f4.png�PNG

   IHDR  �  �   ��O3   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���]l��}����%R�(��(�"mY�-?(˃���S�$]Ңht�:l��u����C�m�i˴�Л]�z�a7	$C
�hs5�r��b9�]�ReZ�����"��8�BQ<�����z��s>�o��/S  �laa�G�"⹈8Px� ����N�*=Z�7�7�^(=   ��.Eę��}��� "6K ��T�  ���=�"�E�gC�     t�LD|:���^8z��J ��� xU�s���C      �ӓ9�?>z��ϖ  M� ��������K�      �!�9��>??���C  `��  <P>�R���w      찱�����=Uz  �� �I�."z��      �TUU���8Qz  �� ��ѣG�^D�.�     `�����ߔ  �"p �����8�s���w      4�_=z���G  �0� x �u��#��;      ��9/�  � p �A�"⟖     РO�����  �iw  :onn�q��     �&���Xz  �4�;  ��R�g�7      𩹹��,=  v�� �N;r��#)�ϖ�     PBUU���  �Iw  :������     Fק���*=  v� �NK)���      JJ)���  `�� 謥����;      JJ)�Å��=�w  �N� �Yu]���      Z�@���K�  �� p ��r���     �6H)���  `'� 褣G�.F��K�      h��.--�(=  �� �N�9��     �6?_z  �/�;  ��s�L�      -��  ��� �E���'K�      h�g���N�  �C� @�,,,<ӥw      ��`0���  �~� �ϔ      �R�Pz   ��;  ]���      Z�������#  `��  tʣ�>�;"�)�     ��R]�~.  �%p �Snܸ�LD���     �bw  :K� @�|��      ������  �!p �k�      wwpaa�åG  �v� ���     ��L�  �w  :c~~���8\z     @��?[z  l�� ��H)=Wz     @���9v�؁�;  �^	� �ӥ      tD������#  �^	� ��;     ��?^z  �+�;  ]ы��Rz     @�|��   �W��  `+���zO�[UUU���݆Q��������p'ccc�k׮�3    �j}}��az�ȑ#�o�����C  `�7  tB]ק�z�~����1111>>����v�~����cccQUU�z=A;���<fggKπV���?O>�d�    [���q�֭�y�f���ō7�ڵkq�ڵ�~�z\�v-rΥ�ދ�~��\D|��  �*  ]�����XLOO���t�߿?���SSS�gOg�     ;dll,���bϞ=q���;>���o��V���ƛo��.]�˗/G]��ݺ���C� @�� ���LLL���|������LLMM��.     `D���8t�P:t�����|�r\�x1.]�/^��7o\�#>Qz   ��;  ]PE�������Ǐ�������     �]�^/>�~�sׯ_�.�믿���zlll\��7B�%G  �V	� h����G��ޭ>_UU;v,�񘙙�4     �199'N��'ND]ױ�����Z���q�����,..>�ꫯ�m�� `;�  ��`08���RJq�ĉ8u�T�ݻ�     `h����������ӧOǕ+W��^�������J#��pD� ��;  ��Rz_����8p �}����      m355SSS��OƵk��ܹs���/�[o�5���9�DD�ǡ�  � �;  ��s~�n__ZZ��~������     莽{�ƩS��ԩSq���x饗��_����}��҇w� `���  `��^_8~�x|���     �6==�>�l|��}�C199��/�����=;��  0,w  Z����c�؝�v�Сx��g#���*     ��ؽ{w<��S��}.>�āv�e����x!  6g. h�7�x㉈�u���>}:z�^Ë      ����8~�x?~<^y�8s�L\�zuۯ�s���x~� �p� h�������gggcvv��9      �{��cii)���ę3gb}}��_#���� ��� �vO��sssM�      (���x�������g�Ɵ�ٟE��^^���  ;�*=   ~�������ɦw      �{��x�gⓟ�dLLL��o=y�ر�a� ��"p ��N�      �6�����?��1;;���ҿu�����  ;A� @���x�N_�r�J�S      �eϞ=�O}*�����|J��C�  �M� @k-...Dľ;}mee��5      �������x���o�q�;  �'p ��r�'��k/^����&�      �RUU�},&''����  t�� �6{��="��_lj     @��޽;������9��GDjf  l�� �6�k�~�ܹXYYij     @�;v,�����ȁ������  �!p ���q<��󱶶��     �V��*:t�gRJw?�  �	� h����������矏����     �j9���SM�  ��� �VUD<������<������-     �k0ĥK���L��Ɇ�  ���K  �;YXXX���[}��W^����|�#����5     �����o����]�I)�� @��� @+UUu�^�+��_���bmmm�      Z���_�o~�[y��� �b�Y ��꺾��="bee%���/����NO     h��^z)����G]�[y|����C��  �%p ��rΏl��޸q#��կ�ٳg���      �s�ʕ��?����7�qO'�����,  �/��  �NRJۺ�~[]���o~3Ο?�=�\LOO��4     ���_���ַ⥗^�ֱ������/��2  �w  ����._�_��W�G�~��111�/     Ш�s\�p!�����������>�S�  `�	� h�	�#������w������O�O<�w�ީ�     �����p�B���k�ꫯ����N��� ��� �:���;��q�������'O���'O��     ����f\�|9.^�.\�����x����  ��  �N��{h�����/��b|�[ߊ�z(N�<��[     ����㭷ފ���������t�R\�|9�n������YYYy��7 �{!p �u��Zl�}꺎s��Źs�b߾}q�ĉ8v�X�ݻ���     F���f\�v-�^�������o��V\�r��������c!p �u�  ��R�ox���8s�L�9s&<KKK�����R�s     ��X[[��7o�͛7�ƍq��ոv�Z\�~=�]�kkk�'���"���  �&p �����^�|��x��7�^�]�v���\������L8p �}�F    �����X__�[�n��������vȾ��7n܈����W��GJ��  �N�9  �Q��������{��^|�{ߋ����bjj*���SSS�o߾����ݻw���x���^     �����9G�9666""b0�����u]���f�����ǃ� ����3d���,�?�Qu]� h%�;  m�Tz�{��:VWWcuu�=���z���\���c����X��J_��W��ٳ�g    r;Dg�\p ���  �Qk.�o���/�hx�(��ݾ~   @+=)"r�!  �NU�  p���     ���\\\\(=  �M� @����싈��;      F�c�  ��	� h�~��z;     @��� ��� �*UU-��      0
RJ���   �&p �m\p     h�#�  ��	� h�;     @3�  ��� ��Y,=      `D/=   �M� @��     �1}�����G  �;	� h���      Fŭ[����   �$p �m\p     hH����  ���  ����̾��*�     `T���  ��� �������      0J\p �m�  �FJi��     �s��   x'�;  ��RZ*�     `ĸ� @�� h���      F̱�H�G  �mw  �d��      ����ѣӥG  �mw  Z#�t��     ��Tz   �&p �5rγ�7      ����  �6�;  m�;     @��  ��� �6�     4��룥7  �mw  Z�رc�1Uz     ��I)�� @k� h������      F�� ��� �
u])�     `D-�   �	� h�^��;     @.� �w  Z!��;     @�=����#   B� @{��     PH]׮� �
w  Z!�,p     (dssS� @+� h��ґ�      FUJI� @+� h�     
� �w  ��w     �r�  ��� ��p�     ��;  � p ���8Tz     �� �
w  �;r��LD�K�      aK�  @�� �v�-=      `�훞��*=  �  ������      0�v�ڵXz  � (.��;     @aUU	� (N� @q9g�     �[*=   �  WU��      �� @qw  ��9.�     �8Zz   � h�;     @y�  �� �6�.=      `��gKo   �;  m p     (,�t��  � �w     ��\p �8�;  mp��       bbfff_�  �6�;  E9rd2"�K�       b||�H�  �6�;  E�z���      ����gKo  `�	� (*�$p     h����  %p �4�;     @KTU%p �(�;  E�u-p     h���l�  �6�;  E����      ���  %p �4�     Z"�|��  F�� ��\p     h����  %p �����      ��;  E	� (��k�;     @{�� @Qw  �r�     �U<�裻K�  `t	� (M�     ���͛�K�  `t	� (M�     �"9���  ]w  J�     �H]�GJo  `t	� (�駟�{K�      �/�z=� (F� @1+++��     �L��w  �� PL���     ���  #p �����      -�Rr� �b�  �$p     h����  #p �����     �}\p ��;  %	�     ��w  �� PL��@�      ����H�G  0��  �R�*�     �16==���  F�� �br�w     �;Tz  �I� @1.�     �SUUӥ7  0��  �s�_z      ?*�$p ��;  ��]p     h'�;  E� (&�$p     h!� (E� @Iw     �v� P�� ���      -T׵� �"�  �ҋ���#      �Q)%�;  E� (�رc�""��     �	� (B� @�n��_z      �I� @w  ���zS�7      ��  !p �����      �%p ��;  E�     Z�PD��#  =w  ���J�     �^c333{K�  `�� ("�,p     h������  =w  �p�     ��RJw  'p ��     �M� @	w  �H)	�     �M� @��  �;     @��u-p �qw  ��     �ޡ�  =w  �H)	�     Z,�t��  F�� �R��      �]M�  ��� P��      �&p �qw  J�     ��� ��	� (E�     �b)%�;  �� PB{K�      ����  ��� и����J�      ��  ��� и��I��     �o��G�]z  �E� @�rΓ�7      ��]�vm��  F�� ��	�     �allL� @��  4N�     ���@� @��  � p     耪����  �h� �8�     ���k� h�� ��      �s� �(�;  %�     : ����  F�� ��UU%p     � � h�� ��      �R� �(�;  ��9�     �A� @��  � p     ���  0Z�  � p     �� h�� ��      �R� �(�;  %�     : 缿�  F�� ����      ��;  M� и���      �s� �(�;  �s�     �3��  �h� P��     ��'J�  `t� (A�     ����S�7  0:�  � p     �]�v	� h�� ��U1^z      [3���  ��� ШÇTz      [SU��  4F� @�RJ��7      �u9g�;  �� �(�;     @������  ��� Ш��1�;     @��� @��  4*�,p     萔�� ��� h��     �C\p �Iw  �;     @�� h�� ���)=      ��K)�/� ��!p �i�      pO��^  #p �Q)���      �'w  #p �iw     �n� ��;  ���Z�     �-w  #p �Q)%�;     @����  4F� @��      �s� ��;  M�     t�� ��� hTJI�     �-{""� �h� Ш���      �R-..�;  !p �Q)���      �7u]O��  �h� �4�=      :&�,p �w  �&p     ��;  M� �4�;     @�� h�� �F���      ������  �h� Ш���     �{\p �w  �6Qz       �&�,p �w  ��;     @�� h�� ��	�     �G� @#�  4M�     �=w  !p �iw     ���9� h�� �&��      �"p �w  3333Qz      ���*�;  �� И~�?^z      �.�,p �w  SU��     ���  4B� @c�      �%p �w  �$p     �&�;  �� И��M�;     @7	� h�� �Ƥ�&Jo      `[�  4B� @cRJ.�     t�� �F� h��     ����  �h� И����      ؖ=�  0�  4��k�;     @7�N�>=Vz  >�;  �I)�*�     ��y�W�Ko  ��'p �1w     �����w  �N� @cr�~l%     @GUU%p `��  4�w     ��J)M��  ��O� @c��     tTJ�w  �N� @c\p     �4�;  C'p �19��      ؞�` p `��  4�w     ��J)	� :�;  �I)��     �]w  �N� @cr�.�     t��  4A� @��      �%p `��  4�w     ���Z� ��	� hLJI�     �Q)%�;  C'p �1)���      �6�;  C'p �19g�     �K� ��	� h��     ��RJ�Ko  ��'p �Iw  ��ha    IDAT   �����w  �N� @��      �R�(� ��� ����Jo      `�\p `��  4&��;     @w	� :�;  M�     t�� ��� �$�;     @G���  �� �&	�     :*�,p `��  4i��       �M� ��	� h��      �%p `��  4I�     �]w  �N� @��      �%p `��  4i��       �M� ��	� hJ?|�	     �ew  ��_z��Z^^���z����ґ�����@UU�1Q����R*��-�@D��Ǜ)�A�y="�kq3���s^����N (f}}�������g      �MUUM-//���; �aUJi<�<����kWD�RJ�rν��w5"���=�9窪V#�f]�k?��r���^�wq0\��_��K�w�"��}�K_ZJ)=]����HD����"b|0DDD�9""RJ?�1�u���V?       �v9�^���Z 5��~x�c�1��v����v㻼���"���nD�\U՟���W~�W�7�yT�w�o��o���깈x6">�r��  �w�      �)�9g��Q2O�������:""���W#�ň��񍺮������_����6����Ω�ҧ"��\D�� �j���     ���ATUUz @������^UU,//�DğD���9��~��^,����[�{��{677&��3񩈘+�	 �K�d     ��s� �f#��"��RJ���|!"��s�r����������:A�~��[�����?�s��`0�k)��қ  ��v     t�`0(= �K�"�SJ�86�����R�������7~�7^/=�������9��9����l���G  ;@�     �}�� `��"�r�?���������?�9��]�v��_��_�Rz\���#"眖��2��Ku]����(�	 �A�s����}�eg]�߳ϝ	I�$Pe����ش�VQ���"(-��ը���ҁ{�3#Jr@��9�d���j��"�6`*��,|c�l�4�,�$& M($s3q^�~�G��I2/����}���]k��������^��]:      [d�; �XT9��F�s�9r�`0�����f�d3�������������L)}M�<  ��4     ���� 0vgG�����8~�����ѣ���׼����2��<��녈�ќ�9��  ��     ��w ���g)���:�+���[��:����ҡ�6S����_\U՞�h�҈�� 0K�     �Ϟ ���~�h4z�`0xw]�����sK�\M���{����)�+"��J� �E�y      ��= �Fu"�������`����~fqq��5iS]pEľ�����
�       �V��t �Y�����}0�^J銥����4)SYp_�Rzm������\  �0��      �g� ��/�9�`0��N��waa�s�C��T�{������WD��s��� �?��	     �~�Ѩt  "���l4����:�������C�KU:�������*"���v �m&�\:      [d� ��rnJ�ʺ�?9_T:̸�~����r4��/+� �S��	     �~&� lKO�9�w0�nJ駖����t��h���s���F���v �mN�     ����  lk/�9|8�"�J�٬V��������9�_���K� ��rΥ#      �E&� l{��i8~`8>�t��h]�}8^RUխ���Y  X?�<      �Ϟ @k<?����`𓥃l�\� 뵲�����9����Y  �8�     ��w �V9?"���F?�w�ރ��G+&���:��M�� �R�y      ��= �VzY�ӹy����*d=�}�}m,��qQ�,  l��N     ���� �Z�����u�����N�����ڵ�@�����  �u9��      آ�hT:  �����~0����՟��zGJ:�m9���o|����@� `z��     �~�|  ��ڵ돮��'�r2ۮ������s�Λ#�y��  0>&�     ��	�  �!���cǎ}���?�t�G�V�~���)�E�SJg `�L�      h?{>  S�))�?ۿ�w�r�mSp����>����8�t  ��w     ��3� `��WU��~����A���~��;���xL�,  L�i      �g� `*�L)�z���]:H�6(��=)�k�C  &�b'     @��� �ZUJ���`pE� %/����F�J�  4#�\:      [4�JG  `�^7�*�X�}0�.�T�? ���     �~�|  �_�y�`0(6ļH�����"���z  �c�;     @��� 03��u��x����2�te�� �,�<      ��P# �ّR�r0,5}�F��ಔҵM^ ���b'     @�;v�t  ��?��+�����6yM  �w     ���� 0sRD��.x#)��߿���;#����  �~,v     ��= ��ԩ��7����k�b/����\PU�{"b~�� `���	     �~u]��  @9�s������I_k�����]�N���I^        �<C�  f�W��ͽweee�$/2��{�9u:�_��gL�  ���N        h�g��ͽ#�&u��������dR� �]�     گ���  (,����p�<��O������-��I�        (C� �5o�9���ྲ�rAD�fD̍��  ��	�      �g� �5U��k���x�'��zU��y{J���</  �g�     ����  p\J��UU���덵�>֓���w#���<'        �=�u]:  �HJ�[�=�ܥq�sl��`����q� ��b�     @��� ��RJoX뒏�X
��]w�Y����9�� 0},v       �T�����3�����~�ȑ+"�_��\        ��T�u�  lO_}����8N���p8|fD,�!  S�w     ��Sp �TRJ{����z�-ܯ���9�GĎ� `�)�       �T���_�����-�R�}uu�?F�3�r        �Lp ��y���Wn��.�_s�5O�9_��� 0;Lp     h?w  ��u+++l��M܏;֏��7{<  �E�     ����  ����z�f�T�}���ύ���E          �N)���:����{UU�#"m�X        ���. �vHUU]�s�p�|���`��ƍ �l��	     �~�|  ؀��n�m��~�7t"��7z           fKJ�M�^on#�l��~�w�<".�P*  ���s�      l�	�  l�����d#���6�}�F @��;     �4Pp `~f#S��]p��;~0"���H  �<w     ���� �&<u׮]�a�_^W�}mz��l:  3/�T:      [�� �f�_��I?�u�o����o)  3��*     �O� �Mz�Z'���UpO)-n-        0�� ؤ��|���p�����-� `�Y�     ��}  ،�ҿ���g쥟���s�=�H  �2�      ���  �UU���-����\/["  f��N     ��P�u�  �T������)���>77���1�T        @k)� �;:�Ώ���,��S���          ��X�9���S�8���D        Z�w  �����N��)�u]�|2y           �a�쪟�����/�X           f�K����O��I�v�zaD�h$        �urΥ#  �~�u]��d����s�d�y           �a'�?�����Ή�N<           3)��=�~��G���������1�H*           fN������G����{J�I        �Nιt  �DUU/x�{�|#���<  lUJ�t        `�9� ���b��
����9���          �z�`0���xX�����l           f�N|Q=��om.           �,��-'�~��~�7tRJ��|$  fAJ�t        `�y�7��9�⡂�w��8�H$           f�y��v�3���N����          `���겟Xp��Y           �a)������g� ��H)��      ��KG  `�\|�UD�u�]w^D��bq           �UO�ꪫΏX+�>|��0R          ����;w>+b���*          �6��6b���R��e�  0�R��      �i�s. ����k�����f `�)�        ��Rzz�?LpWp          ���+++�"�+
� `�yT%        p_y�uםW���=�t        �6 `R>�UU]�O* ��R*        �ƪ�zR�Rzb�         @;�� ���u��*"�          (�UD\P:           �-���*"�Q�   L��R�        �6�s~\�+        h��s�  L����;           ��㪈xl�           ̼�V9�sK�  `���JG      `��  0A�V)��S  0�,t        g��J)�,� ���        ���*�l�;        �. 0A;���+� ��g�     `:�� `�vTq�t
  �_UU�#      0
�  L��*�t�t
  ���N     ��`� �	:Z圏�N ����	        ���*�l�;  ��     0��  0AG���j�  L?�      ӡ���  �^�W��)  �~
�      ���  ��R�b_, ��g�     `:�� `Rr�_4� �FX�        N'���*"�_�   L?w     ��`� �II)}���ϖ ����	     0��  0)9绪���t  ���N     ��`� �	��J)�Y:  ��B'     �t�� �����4� �FX�        N'�|Wu����J `�)�     L�>  L�h4��ڷo߽�w��  0�,t     �_Jɾ  ��}���[���T�(  L=�      �g� �I�9*"���H)�U�8  L;��        ���W9�O�� ������_     `[3� �	�ˈ�����Y  �v;     �Ϟ  ��s�h�Z���ѣ�DD.� ��f�     ����  0!ynn�ck�}����.	 ��f�     ����  0!���𥈵���[
� `X�        N����P�=���2Y        �60� �	���?N,��L  fAUUg�      ۚ=  &�.�Cw���w��"�`�8  L=�<      �Ϟ  ������_<Tp��z�RJ.�	 �ig�     ����  0�����g����<  ���        �I�ɉ/Vp����� ��Pp     h?{>  �[J��'�~X�}yy�/"�F 0,v     ��=  ��s������7VpO)���F# 0��:�      ��� �����:�9Y����        ���;  �s~�#�{T�}uu��#��F 03:�N�      l��� 0.)�C9�?x�������z��w  ��b'     @�j ���߻������j�k�y  �1
�      �R* �)�R:ig��-�����E��D 0S�     ��w  �!�t����?�g'm�z�C��&�
 ����     �~&� 0u]�{yy���}vʖQJ魓� ��Qp     h?{>  ��)�ꧼ�\\\�����$�  0{L�      h?w  ��o�����Mp�)��O&  ���锎      �)� 0oI)�S}x�;Δ�["���# 0sLp     h?w  ��hUUo=�N{ǹ��xWD�8�H  �$�     �O� �-�����)��3�|���  0�,v     ���F  lEJ���3�����?>�D  ̬�R�      l�=  ��楥�������Ѽf�a  �q�y      ���� ���|i]w�^x��-� `���     �~
�  lҧWWWߵ�/����K/��V��	 �Yf�     ����  �9�_��z����u�q��Ͽ#"n�l(  f��N     ����^  6*�t����������[F�_~�є�U�� ��Sp     h�N�S:  ���^�wd�_�P���O~�/�?��L  �:w     ��3� ������[6r��ZF�^z�(�t��2 ����<     ��P#  6"����/���F���g��}wD|x�� 0��     گ�锎  @{�����=h�R�/"�&� `F)�     ���  �)G�rJiÝ�Mܻ��"�77s,  ��D     �v����� `���~c�s�a����z1"����  �=      �M� �u8�Rڳك7}ǹgϞ��9�a�� 0{Lp     h7w  �$�����Ż6{���8�;�k"��[9  ��w     �vSp �>>??�VN��;��/��hJ�#��V� �l��	     �n�{  8�c�c�_~����[��\ZZ�hJ�ꭞ ����tJG      `<� ��t����Փ��O*w��qeD|b� `zY�     h7�  8�������8�X
�w�>�s�ш��8y  ��O     �v���ԍ  �.Gs�?�����8N6�;���古�^7�� 0}Lp     h7w  N������q�l�w�|SD��8�	 ��0�     ��� x�]x�+�<�X�8{�^=�~8"�0�� 0Lp     h7�=  �����.����8O:�?�ܻw�9�E�X� �~&z      ��'� ��������{�O<������SJWN��  ��O     �v�� ���v���O�������Ɯ�oM��  ��O     �v��^  "�w����4��O�3���:���['u  �ł'     @���͕�  @Y��ܹ�R��&�0ڽ{�}�N�E��I^ �v0�     ����  ̴{�~��ݻ��E&>BsaaᶈxaD�?�k ����     �n�� 0�H)}��={>=�5r���vo����Q� `{��	     �n ̤QD�����MM\���Q�۽1"~,"rS� `{��J     �v�� 0srD��Z�����v�o�9���k �}X�     h7�=  3g_��}s�l�����|]����.  �UU㷟      ����\�  4��nw�-�0Z^^����ĵ (�D     �v�� 0r΃n����.6Bsyyy9"^_��  4ς'     @�yb/ �Lؿ��.��g�۽2缯d  ���     �^UUEJ�t  &(����v���P�O*���WRJ��Kg `��     ��^ �T�)�奥���ˋ�#"���)������  09Y	     �^
�  S�X��'�����Dl��{D���ү��^��� �dX�     h/{=  S��������_)�mSp��XZZ�ú��w�� ��Y�     h�����  �;���n����AN��
�{��e�ΝGćJg `��     ګ��]� �ͻ���|ݞ={n)䑶�]��ݻ�޹s�wD��Jg `|�     ��^ �������maa�s���̶}n��ݻG������)�AD�H\�    IDATU:  [c�     ����m� ��9�s�.//�b� ��-'��hyy���ƈ�t�,  l��V     ��aF  �R�#���۽�т�{DĞ={n9v�س#���Y  �<��      �e� @k�x���g,--�T:�z��A���7"�w8^�s�>"W:  ��     �^ss�� ��"b���t��hݟU.--�+"�6"��t  6F�     ����  �������m+�G�����vo_]]}~D�:"VK� `}<�     ��� Za5"^����M���]:�f���A�^���kWVV���t������ ��yl%     @{)� l{���v�����o�ݻ��q�`0xID\O*	 �S0�     ��� ��;#�U�n���A�ajF�n����է��E���y  x4��      �e� `{I)J)��F�����1�O���E���W_�ku]_?ST� h;��      �e� `����,,,�V:̸MU�����Ż"��~���RJWD�K#"� 0���     ���; ��������vo.dR���~�������K���3s�?��� 0�����     `�)� ����~vqq��K���h---�E<XtND��9�8"� hXUU�R��s�(      l��; @���{"b����M��4e&
�ǭ��}Ɂ�Z���r�?g�� 0K����hT:      �i�  �9����iaaᓥ�4m&�:>�:p������҈xUD\T8 �L���Sp     h!� &��9��r�Yg�e���w�S�L܏[XX�RD������9�����.��F�Y�� L-�      �d�; �D��߫���C�}���ե��3"�~>8p��c�����e���ʦ �.
�      �� 0V7G�;v����Y��~2�:am���Fį��D�Kr�/N)����� �"�      �d� `KF9���RzOD���vo/h�r�yk�8"��`0��ҋr���_V6 @;Y�     h'�<  ��������rο���|O�@m�s����=�x[�׫�9�g���=�������xlр  -��x(     @�ر�t ���K������СC��zu�Pm��	k�h����s��k��꺮����礔.���"�ܢA �!�=      ��> �����9�RU�MUU}�կ~�_��r�`m�s�~?��󶈈^�W���_u�ر����RJO�������'� �L2�     ��<� �AG#�o#�o"�orΟ��O���}��{����Jd�:
��������<⳹��?��ǎ{|J�	)�'�u��qVUU��9?&"Ύ��a
�vw,"��.�9?����D�h���	?D�߯� 3�ȑ#�O*�     ���9�N<8� fI'"��:�:᧳��s�{;"b5">Q #�s(�r�联���u�ň8\U�=9���??77w����{w��;V �LSp/`��sk?  3�.xgD|�      l�[��֟���?�K�  `�U�  0s(      �����P�  L?w  ����      �qw�}�}  &N� �F�-|     �ϑ�8V:  �O� ��=P:       f� �F(� Ш��Lp     h�C�  0� hT�Y�     �eRJ&� �w  �f�     �er��x  h��;  M3�     �eRJ�Jg  `6(� Ш���;     @˘� @S� h��O     ��1� �F(� ШN�c�;     @�b @#� h��W     ��=  �� @�Lp     h�C�  0� h��      �c� �F(� Ш��	�      �c�;  �Pp �Q9g�=      ��  �Pp �Q���w     ��Qp �
�  4j~~^�     �}� h��;  �:��-~     �ϡ�  �
�  4��[o=��9      �C�  h��;  %.      �1� �F(� P�	      -�s�� @#� (�(     @��� �
�  �`     �ERJ��3  0� (���      X?w  ��� @	�J      `������  �lPp ��     Z����7� �F(� P��;     @{�{���  �Pp ��C�      �n�"�. �٠� @	&|      ����  �
�  4.�d�;     @{��  ��Pp ��     �C� ��(� P�	�      �� @c� h\]�&�     �DJ�`�  �w  J0�     �%r�&� �w  J0�     �=� h��;  %��     �K  `v(� и��	�      -�R2� ��(� P��;     @K�u�� @c� (�P�       ��	�  4I� �ƥ�Lp     hw  �� @	&�     �DJ�`�  �w  ��tLp     h���Mp �1
�  4n׮]
�      -�RRp �1
�  4��[o=�J�      ��RJKg  `v(� Pʡ�      8���Lp �1
�  �r�       ���Ç� h��;  ���     �sssKg  `v(� P�	�      �_���~���!  �
�  �b�;  ��ۻ�9ӳ������n�7Yd��,k,Y���@H��D�!eI@BBd�a�r��d�'$�x�v������~� ��C���y��kg�]��޼���.   �w��ҲG  �>�  dq�     �w�  �^�  d�     ��N�   ֋� �,��      �J.� �Tw  ���     й�� �Tw  Rx3     �����  ��;  )�q���     ����;  K%p  ED�     :�Z��� ��"p  ��     ��5� X*�;  )�q�     t."�  ,�� �.�     L���  ��;  )�      �s� �e� �b�ϲ7      �r�5�;  K%p  ��      ������  �z� �b�;     @��qt� ��� ����w     ���� �R	� H�����2f�      ��Ο?�;  K%p  �XJ��=     �:���z�= ��"p  ӝ�      ����  ��;  �>�      �d  `�� ��;     @�"B� ��	� �$p     �Tk�v�  ֏� �Lw     �N��\p `��  d�     t*"\p `��  �i�	�     ��;  K'p  MD�     :w  �N� @�;     @�Zk��7  �~�  ����      <��  d� ��w     �~�� @�;  i�      ���w  �N� @�q�      ��A� ��	� H�;     @����ogo  `�� HSk�     tjcc�w  �N� @�Ǐ�     �Ԯ^��Y�  ֏� �4��̛�      }�[J9� ��� �f{{���Ҳw      �7�  ���  d:*���     �� H!p  ���      |�� �w  �d      ��  �� ��w     ��� H!p  ��     �?w  R� �&p     �� �w  �	�     �#p  �� �T�5�;     @gZkw  R� H�      ��;  )�  �r�     �?�8
� H!p  U�U�     ЙǏ� H!p  ��      �y|�֭;�#  XOw  R��(p     �˭RJ� �z� �j6�	�     �r3{   �K� @���#�;     @_�  �� ��_���     �/w  �� Hu���ǥ���;      �w  �� �+�      �� �F� @�      �� �F� @�      �� �F� @�֚�     �w  �� Hw     �N���  �� ��;     @'�  d� ��w     �~��(p  �� �t����      �֗����do  `}	� H�Zs�     ��.]z�= ��%p  ]�U�     Ё���� ��&p  ]k�V�      Ji����  �z� ��@      ���  �z� ��;     @�  �� ����X�     Ё֚� �Tw  �-�{���;      �]D� H%p ���      ������  �z� Ћ��      ��8�.� �J� @/�      �j�w  R	� ��~�      �u���)p  �� �.��\p     �������#  Xow  z!p     ��z;  ��  t��*p     H�Z� �N� @/�      �"b/{  � �BD�go      Xs.� �N� @/\p     H�Z� �N� @/�      �"B� @:�;  ]��
�     	� �� �.\�z�v)�({     ���q/{  � �E+��&{     ������ @:�;  =��=      `]mnn
� H'p �'w     �/_�|�=  �  �d?{      ��r� �.� ��      	Zkw  � p �'w     �!p �w  z"p     ȱ�=   J� ��;     @�֚�  tA� @O��      ���� ��;  ���)     @�k�  ��;  9::�     $h�ͳ7  @)w  �"p     H0���  tA� @7�ŽR���      k�p�X��  �� �+�      Kۥ���  J� ��;     �r]�   �� ��;     �����  �sw  ��Z�     ,��  tC� @W"B�     �\.� ��;  ]�     ,�� �n� ��8�w     �庖=   >'p �+���     `��� @7�  te�     ��p�X��  �� Е�
�     �g^Ji�#  �sw  �r�ƍ���{�;      �AD̳7  ���  ��z�      �u�Z� ��;  =Zd      Xײ  ���  �h/{      ��p� ��� �Nk�w     ��� ��;  ݉�;     �r\�   O� �#�;     ��� @W�  t��&p     8{����F�  x�� ��D��     ���K)-{  <M� @wj�w     �3��  �,�;  ��q;{     ��k�meo  �g	� ������Rʭ�      +���  �,�;  ��      g("�  tG� @�Zkw     �3�Z���  �%p �Wײ      ��Z��  tG� @�j���      V��|>��  �� Х��<{     �
�*���#  �Yw  z%p     8;�f  ��� Ыk�      V�� �.	� �����     ��� �� �.-�{����;      VQk�r�  x�;  ݊�y�     �UTk�u�  x�;  �j�	�     ����� �.	� �ٵ�      +ho�N�  x�;  =��      ��~�=   ^d�=   ^b�Z+��� /t���rpp�=���ѣ2�c�    �Rk-E� @��  t��6?<<�]������׳g@��Ey��a�    ��/}��R>��  /R�  ���֮eo      X5�V� �� �n	�     N�� �n	� ������Z���      �""������  �"w  z��      �
"��Rv����do �� е����      �
��d�  ��� е��V�     �U�����  �2w  �VkuE     �<��.p �kw  ����     `DD��;  ]� е�l�MV     �S�$p�8{  ��� ��=z��'_�	     �[���������  /#p �k7nܸ�;      V�/J)-{  ��� �)pI     �-DD��^��  �"p �{�֭�      S�����  �*w  ��Z�${     ���ZK)���  �*w  �7�k"      o��Zj�>s �{w  �7�k"      o!"������;  �U�  tocc�W�=     `�"�J)c�  x�;  ݻr��^��a�     ������  pw  ��E�N�     �)�����G�;  �$�  L�V�      �)� 0%w  &�����      Smss�g�;  �$�  L�0���      0E����u;{  ��� ���yDdo      ��Z�G�  ��  L�0��     ���(�0|��  NJ� �$���Ok���w      LI����x1{  ��� ��8��ne�      ��Zk���d�  ��� 0�q�     �)�����ٹ��  NJ� �d��Q�     �)q� ��� 0%��     �$"��Z��  ^�: �ɨ�
�     N���*�w  ��P 0��엵�1{     ��Z˹s�~��  ^�� �����zW�w      LA�u�ʕ+��;  �u� ��a~��     `
�a�Q�  x]w  �惈��      еZk)��w�  x]w  &����'o�     ���w  &G �������     ��axx���w  ��R 0)����Z���      =����ҥK��w  ��� 05���Q�     �^ED��~/{  �	�;  �DD�     �.�P"���;  �M� ����Ok�(     �<�0���d�  �7�
 `���     <_D\��緲w  ��P 09���G�0<��     Л�(����  oJ� ��\�x�q����      ����R���  oJ� �$E�k�8     �ak����  oJ �$��~$p     �]�0|o>�?��  oJ �$���'_�	     @)��g'���  oC� �$]�v�r�u?{     @/�a(�n�  xw  ��E�k�H     PJ)�ֽ���f�  ��� `���     �����RJ��  oC �d�����0d�      H7��J)�;�;  �m	� ������#� {     @�Z��W����w  ��� 0e���Z=�     ��Z�a�ǋ/>��  oK	 ��E�{�0d�      H�䳒�d�  �� p `�Zk��;     ��f���Rʻ�;  �4(�  ����݋�0lg�      �Pk-�͝����[  �4� ��VJ��'_�	     �Vf�Y���g�  ��"p `���     XG�0�r{{��;  �� X��� {     �2=������o� �� p `�vvv�R��V��     ��������7�w  �iR  �*�9�Ͳ7      ,E����wׯ__do ��$p `%Dķ�a���     `f��8���d�  ��&p `%���܏����#.     ��"��f�o���}��  N�� ��Qk��l6˞     p�666Jk�w  �Y� �2���{��̥     `eED���������-  p�  ���Z�+W�    �U���qw�?��  gE� �J�����l6�u�     ����c�  �IDAT6C��/���v�  8+w  V�q��/�a��     p�Ν;�㝝����  gI� ��������s��-{     �i����Mk�OJ)��[  �,	� XE-"�l6���     �f��݈���b�i�  8kw  V����s���iq�     ���l�����{{{?��  � p `e���~kss�K)7��      ��Z��l������������{  `Yf�  �,-�*�|�TJ���X=<x��͛���:�[Jy�=  ���ZJN�Ν���͎�����f��8����儍Gk���x*��g�M�^��~ "�k��[��Q)�=��G���q)�w��a~�5#�?���Xk�=����s�  �v���R�y�L    IEND�B`�PK
     $s�['�Y��  �  /   images/4bf63cb1-3675-4452-8ab6-1403298522d5.png�PNG

   IHDR   d      X�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  SIDATx���KA�_�&�Ҕj�PZL-1����?�7O=x��[�ދ'�{�xl=x#"�P"�ɖ�T�[b�&���ݢv��xa��o�;o�f&
I ��ё��v��F��5�M������Yj�ۧ�����ZZZ��v�����$��\�v�T�)�Q�Z���?�;r�V�B�x�1E����� &M6���������FM�0��UUu���[�;<<$��K�Z�L���B�@�LF/_7Ft�o}<YB��.��Ȉ�8��p�\�b�hY��|>D�A=�\����l!�>����=�����y�ϐ!v�[V�������ѓ�=��a��ò���;�\��)�mr.�&�277'�A,C�d�����ƉpF��F)�uI�
f�`���(_���X��N�ǐ�v�����4�q$����"�q�	T���.�[�$�F���E��:MdW���a��n��4�'�b�to���f�����<��.�1L� �=�%n ���r�F�I�wQR�V!��{�G"[��Zbh_+���Ol3$����%��;�'���������(Ϥ'�0�j�����U�99��Xf{Ƕk�Cv�8����
�����v� ;;;����W��t)�x�D�ֱLmll ��PX���ښ^����.�P̂(p$mP!��/eqqQh��!Fk�\��jX� 8.1�d�"��{�n��Il�~�&#��r���>�t�z�JE���>��-��ޞ^�n�a<I��+nDE#E������O�[V�0��T*u�pZl�k'���UV�R1�n�y0q�<��>���$���I�"�t}�4���������J�u�    IEND�B`�PK
     $s�[Vm�80 80 /   images/9ce856c6-be81-4769-87b3-53be9928d02a.png�PNG

   IHDR  �  A   s���   	pHYs  A  Ak!T�   tEXtSoftware www.inkscape.org��<  ��IDATx���	|e��_vs���@iI�3��5�X����(�"ʩ�R��'(�x������(7価 ��(Vc��&)G�+M�l��/ݩ�4��f�wf���3��M�����;�3�;�[:00 DDDDDDDT\�BDDDDDDDEǀNDDDDDDd t"""""""0���������� �DDDDDDD`@'""""""2 :��)+S�L�v����/))���X,[�-��?'DDDDDd���QW_��r<\��UX��eq__�;�l�͢��
:k�ĉc***����Xf`�K���8��8��o;k"""""2ˆu�����tuu�ٶ݊��[��簞��^�`/�w�I���8��e����}���������1䀏a}�x˲�a�������sZZZڅ򂡋ֳm;�՗���e��l�p~8և����!���>�������ΕB9ÀN���d2y.��0 DDDDDD�@8��+**~�,q+�/�F���F�ݧ�Kjjj����z�8Qt��3�>ݶ퇓��O�īBYc@�!<_�,���Q������FF{�j���5�CP?A���1��H8�200�Gl~^������rK���
����9���g���N�Z����l^�e��O�oVTT|ɲ�����Bia@�8۶w��N,"""""��	���܈L�5k֜�t��B�ŀ�a�e���/ج"""""��8nԨQ�'����ׅ�Ā�A'NSQQ�W�����������G>yɶ��b�+�6��c��p�����I�������Q���,�@H?g``�_�C�=���v2v�Ǳ9E�������s�[�Ue��q��B�1�{D8nĎ�6'
�َ��Ȕ)S�X�hQ�� t@8���al�""""""w�Too�3���D"�����|*��}�pNDDDTp�@@���&�u�mo�x�O��D�k2�|��������U�s�.
�l���|k!"""��C��RRR��ߕN�O�B�p?K���ƿosx�6c�����q���O|�ݥηE8����P�����?�V6���{}�qoo�`e���ȱv�Z���Q�FIii������"� rq�����P˲���|�?`t�N[���nl� Di��y���M��p���������n�s2�ާ�l�u�e8FVc{%֫�W��{�߮�z��,���}�7��J��ƿ�q�;v�{���F����ܛ�sGṣ���K��c�g+����;��ߴ�1Z����x,~>F���>�R���]K������e4O�y���|�5�6��#��� �Z_qi��D۶`}���a�����
"�H6!3�@���e�);�2���ë�/�;t�>��l'��Xn���?_VVV������e�|s�}��H��oTUU�G�_ZZ�->������zBj{[���mɺYLʄ�ȴ�����=z��t�6S�_�j�ōP��ڲ����ć�]&;�y�qZ���\�ز��������i����,hӅ��Dj�m�mQ��P�oO$��>ǟ~~KS˰P~�L�4i��k�v|���5,,��B�YK-�m�(ϴ�r���RVV��t*87��2�۷۶�[,{_|��E�kPѸ	����T�F��VsJS;��X���.���kjjښ���
D�~��Բ`��W__��5kj�&!�O��&�"��}����
Q�.�AI/���lM�B�@8w�����~���]�*����v��K�"FTH��t�m�~��wP�� �|1��Ŝ�}����c����uuu[���=6�l��z{T�S���i@_�j�`��ޟN�/
�P�n��)ؼ^|��%����$&>ÐN�����ؒΏ􊌆�P!x����o�B�N*БO���%�|��ɓ�C9����Xvďv���I�k�hz~q�M�-u�k^���� ��秮��.
�*Q�_��!�
AOjzr#_�{��@�����X�USS�_vG��,^�xp0?,����<n��i*6?��IC�`x��NqZ��=��W�y������,�	�.��{����)_��\��s 8Oґ��-��G~娆�18C��ڧ�!���1�b�����#]j�|���@����4�p̜����h4:O|��puuu:�����)��pR�m��0�'�y�d����z![ũ�P�l�J����ik;�����`h���S���X'� r:sQ�|T�	����������8ysD��t�N��z�Ԁm�n�2������|�DFK��?�ZM�2e�o3�/�~�;��B��LǦ��q�ʄ3ی��iYց�x�)�8t��`4�
}C:��Os��(_�w6��x�4N��	�G,Z���'R� ���7��}�4`ߟ��GiK��oؚN�к�ޞ�7(�:�s�b
��tʔ�R8#��K�X�����X,��_�J�{���"'NS^^>��~x�)Y��^)�Nk:�c���k8O9���=�����a膪������!�ҥ�����jn�B�\���g[[[[��>���s%VsS�L�:���>�о7��B��\L��t��B��y8���|�c@7T2�<Ax�C:m�r���	���D�4���b�"��u^���_��Zj��4l� Y��>Fȕ6��MG{'b8_�P(N$Q�(ts�$��t����L�R�}��)�����I�m!��J�2/���������sO�����w~�����f���Ӛ�������C8fb}�x��,��;�t��9]�9�(�^N�VlzU�5,O"<Y]]�,�;#*��1���~���^VV�G а�K��+hǹ7���Uw�a8�(��Ot*$�<Oὲ�s�13������I�ӧE;ʭGQ~=���	��Nd��=��w�4iR��Cp�~�Jk4=�ioA���z�0�i�p8<=��b@7N��e�!ݿ8}Z�i+�+������D"�`�>�k�c�J�P(T�s��@���nI�uڢ���q:6o�E8�A�>��s˟���p��ߠ�u1�S��$�qL�BYcH���T7���� �sR�@��%��X=�Zt&��([�q~(�wl���DÕvyשش�Cޓm8�@��AhO��f ��G�NZo�[���?+ŀn�`0��� �F�!��j^�by����]�t�
!"O�D"���B۶���(*��?��m!dWNk:�c�l¹~��Q��b�}��^��ߧ�������p8\���t��/�����F9�J���#`1�{�O�/|��8f����D"����u�&����b�c5[����-Q�jH�"ʅC�Ӹ��*��M�:��ݲ	�#�]���t]��Ч��U<�� ��X��)��z��W�6�7�j��+x�ޣ����V�`�/h���~r*����(,[��h�v�q�n���ekl��u�m��e@9���5����o�+v7�5���'4M�{X��ywj�=��{xK��.�ﵷ�������XݮK]]�(����wp>�c�m'T4z�ZϏZ�ak�;e��{���r1�֑u����:��|Z�)��������`�I(vZ��*��`�M.0�{��n��k�EX��ػ+�����&��q��#�9��Tʺ�=�	^�M7\hy��u�\]W��qއ�m�^����w�bݒZ���Z��[�D��z����h��ǹ�e��W�9)�g*0���̙��)r�Lù����A����.
�b@7�'� �c$W�������0��Ő�nz�FO\n�?�PQ,�᳼��5!J�^\�m�����L��j��t�v�7
�[k���^˃0�5֓������@�k��5�o��obY����߱X���cV��-����������3p*�<�M8׋0��)�!]_�%ӻM�2'u��3��m7Wj4Xk8��� �]m����OX�ߗ3��2, t�ikk{�+�������	�pUa����*���Zk��	��n8�r�K����*�����>��������㳝��q��k��2��(�]���7�s������x�t�8ӱi�'��è8���ܹg<��w�{s�9�Ǐa�P<�G�Ap��^\J���2�;r��FOVZ2��O+����s��l�_�C�������f^������W竮�qR�uH[�u�e0�c����y�����F[��4�>5u��Cp}�_���Xkh݋�=�7=�Kmm���G�o=	�^�O�y�G5l�5�<N�4S�P��+W��a?�A�)�v�_����w�g�U+�S j�Cf��iYӦ�gp,ތ
�=�-�r��S���X�B�`��w:Y�S����T;��oWѺ����v����w׏�������g0��D�-����f邿��I��8,�WNK(�c3��E�i|�p^���SJ߫�R�S��R/.T��h-����Uk�S02��E�^<1�d` ���Hohiiir5˲G�����+/Zy�ܲ�.�����b���x��}/VVV��JO�X,֌���~
�>��x2��/	�X�ݧV�^��5��'�p�
=���>��d(?\�y(��I�����e��B�ۤ'=��
C�Y�� i��'����S���C��!��:������Z��7�'��,//��#�ʭ�u�8q�9�����Щx���|���UgB�Ǝ|2FCI8׋���Μi�M��Ὅ�a@7D8���u��BB�\ޓ̐n��H�4,z6ʋ�%�w�<��-eee�`��$цth���b?�F��UTN���^YY���[�;;;�f�u�.�X��u�O?k�G�Z�j�ᣐ�8����sG.�;ϔ�s�:��a@7�1n��Y��'=�68�
�ӧ�mN�7c}u<_ �i���^��;?L��6���Xסּe�j�7�y!�����7u���/_~����� a�zN�X/Z�� ��a��%X��H���4|.�����kA׮�.,�՝�i�eH/�hW;ڬ��܀��� K���iK":e�r��t�����.\�'�;t�m[�R:����PN8�霎-8�m~�se@����s��L1Z��yA�!�0�B�^E��iC�
�|NI$/�Ҹq����z�����
F�AX���}%B��8�>��1�����+�V�e˖���l<��Јq:���e8/V�w��t��.��V�<���0�痶��j�<Z��j��yo9i�!����<G�rC>��.�[�Ձ���9�� ����V�9���	�o`9A��9O#�LǦu�b���5�n9/FO[}�.���i	Љ6�{l5� *�O���B�#��6�}�F���M���X-��a]R#�WWW?���d�ȝ�X�_X���~��T�,,uBYs�c���8[��ѭ]�}�B6�i�m�]������6��{�6I�܉�h4�/!���<t��I��K�K׏��ѡ����
M$Q1X���2��kjj���-<��pP��i�7،���g�G_��#�>�W1�S֊�奐��!}d�Ĥ��,�?�ȫ����f7vJ�����v�?T�a}��k]��	S�_O�BzR�����~�����D��5�ӱ�/ߍ���7��LݖL���P�)kz���M��Czv�K�8�V��^������٦Vl�L(_o�qt��k�$*��X�@X?����Oc�|?{(b�H$�&VgTWW���Wo�e[��9ӱi]ȍSJ!zj��ߣ������ߢ���9����}N�-9��dC�B��BcHO��GZ����#X.��b�
Q��h������Ac;���D[صu]��nb}���4�,Y���B�Х����<�"���c+d��-
y;������bI���ѣ���D�ǀ�szp����n6�J���)=��u@3�O����.K��è����&!��`q�d�uA��C������!���;;;W�!��j�����/555_@�G��K(#έkZ�tl�z��B����;p���%}���h8���S������r�`�4\i(ӂ�\���bH�4-ȝ���i��o8~����*D9�c�>����"����X}U�����p8�2�_h�>�� ��t�����M���ʥM�}Nk���~�M��:>���s�5��E�������Ӗt=��`�4�k���[��J�v�1�;C����|�r,7������%B�c�X�۲����=E�ܣ�����u��ض�ol?��L�
�D�����|���r�p���8��ڋR��ck���\�4gB�^z�$W�׹ؐ�p���y��i�[�3	�z ��*�ô�Y��u8}��c���������UB�G��܊��)B�^����,�z��am]G(x��ehj>��jjj~�c�G�>NXGN��4��-�;�;�:���K6�p��@����
,�9>�!Ε�LC�3G�Cz����!�ӧI'��a��2uO#Q�E�ѧj�	����r"�'���u#�?����z/�zg��T[[�[X�TWWw!�q:���)چ�qk�י�7�Ы߁.�],��̹Mթ��3��yv��#���i�uW��g�h�~�>o5�ptIii�5�*�
M�#�ߎ��\!�ђ�s��p8���9�SܓH$b�xC�qD��c�2s�������!8��h���tl&��i=M��k]ܙs\��t��z>ourD��<k�I��gҝ�6z�N��dspj�����k�SH�6����ZA��,�X���f,��e��[��m��Q���{R������[UUU�B�滺-lQ�,g:6mI�z����7���b�td�yn0��feҕsOG�t��l�뻆q�>���s�Tz�[W>q���q\���l� �[�
�#�,��T!�>�44�nD�������I�V0�n��B��������X8�f8�4{�5�M�X��K8�ވ1�Ӱ���ٴ�j��{=p�Bz�6nNW|��t�o3ȓ��\��Dƞ�QQ������e�(?/"���囨3|Ӳ�V�kX�F��(P%en�3kjj.�?�uSʱ.=g*0�ic�[1���<�X�PZ�.�#��A<��鸼ҝy0���>m%�?����zѢE]b�I�&U��s	N��ض==5�0�r�-� ���o�"���I�EYxo!�z[[[�3Q��Σ�5��l��,�aݍӱ1�O{�j8��a@��iHׂՇ-�is{H��i����y�����x<��
�^)*��`��X�L������ݛ��|98�i��s����
���z<
���B������ά���#��(��$�[8!]ot���i8מ��[�8B�N�dH�[C�3MJ>G�4�����<�%�`�px?T<�,��xZ{{��0�.��r�0�m�6��������H��X�rz��K����G8����LnMg8�^ha8�tʘS����5#n�>�>m ����F�����؜)�L��-?�m�vu�����;Q�\!���hc�sP�x<���O#�%�.�� �Nk����Ŵ���p><��2j'4�tʊN��!]�+�MsCH׫��H�>�
���!�?'�;�Ptvu�#��퇱�%!���0�=��{t;��:��EX��>�iM���Iӱ1�O[�+*��K�m�)kΈ��C39��l��(����M���^���'l~2������h7wt�����8���Y�P��@ �l��8���tl�tl��Ӌ)�yǀN#�!�iI��<�iѐ���I]���6υ>�rIii�---F_IB0��_c9]��ξ9���/اAeRg`��h�x$yS�H$Vcu�eYע����;ʼ~�E�L�V��t���9cP�1�ӈ9]]ؒ>4';��IP�'L�68 >����;�`����B�����K������p8|�����BD�11Xj��o���!�^8��8��ν�@��|xl9/,t�	�%��Њҵ%�'�=��;�X�Yg��Ζe��{��%�uvv� �_	y*��cŀN$�ǃ1��7'�H������eԛ.�v��z�W�Z5XW*�tlzA�u���`n�8~��N9�iee�`A���V������j����Pщ�o=+�?(��B��@@��ޓ�ӳ����gWw�þ�$*��Cd��������{�ԩS����:K��7�i_�=�ӵ���p^�S:]�Ή�oh��dS��B~h5�Ae�����ϟ�p~��ج�ӯ�3��������m:U8����5�����u$�+&M�tg__߯P7�1�)� Z_�u�W�z:6���ic�3 4:��[l��`�ǖ�M����~i5דǘ1c��1��Ϸ���b ۶CX]�p^���weWwHusg@'_sK������.�ꫡP�O8G\��݅i=�@.Wu&���1�:�Ӫɐ>�|�t�⬭�^����1v�؍Oc�������b���Ʋ���s�y��B�^����F��<+�?gYV����Iӫ�D"�x���d/��X�?/4H�L�tl#iMg8��X(���44~��7���eH��X[���Uzk�s=y�流A��i8��fC~}9����Lf���%�w�D@���w�ȟ�O�0�e�=���=y���p>��O�,���"��u�l�f8�<�c��v�:商t������J.B�3
��/����|�Ǿ���ojjz[�(5܅X�'ŝ�v��w��Lȳ��ݎc����)/���x���N������3�w���{��@��|��si��t�;=蝖t��MIH���|/ғŖ[n�����X�Ķ�ϧ�!�� p��EMM̓mmmo	yR4���N��"�A�	�0���o�Ͳ�s������{�ʕi�+�p�yl97:C��2�z��.�^�<���.N�r�����ܹsڭ{���ۭ]�V[�O�T��7|����N���n����x����Iݦt�m�wa���Gr�j:6���c87:�ҵ+��G�V:!]��;�y�^7n\�'��+V��CR �e��[[ͷ3��x6��d2y�t�w���"�X,�����t�z������ش5}��͜��hӜz�ގJfa@��ڰ%�!}�4��紩.��Z�'����IB�Mj�t�`qy赵�����u���7x�G"��B���0ض�#�O"�@����P"�x����9DO"7�x��#����N}i��o�ַ���pn&t*
-�>��H8���t�O��'T��<'T��e�]&.X��S� �_��P��B�aTX�ы	��x�[,�B��誥�eVg��������B�u%m ��Ou��4�ex� :�sϋ^�dH�4'���`/_��U��F�����w�c:u�y��N�l����	y���P!���5�����s�s�H�����]:::t&D.���<&��p+Cq�@f87:�Ӓ�W<飜ڽzX��y�b�U�a@שӂ���^�!ŝ:mD�/]��F�mB���/ض=�3�����b1�`�i�.���0�׋;/ S��>�LMG�ÀNE��z(��M�b8�@���G2�{>9}�����{e�/�p�7��u�.���
�,��"������ۇ�����eY���ϰ��$K���s�p��d�t�ЮU�j^��Dj�������v!��㡗FR�B8>.��&�)���s���.vs'�{T�#RS�]���(γ7b{!_Ӗs�{�{0��14�khs�#o)P��Ǝkll<���)�IP`��{�6�ŃP��r���O/^��C�3ZZZZm�~U�ŕ��9��WhH�x|�T���tޛ�SN�vrt2��ҽ��9�Ǐ�B�ݷ��z����9�'8����Z�����8��y
���q�1����{{��t۶���4!��9��݉���!][ҝQ����C��X,vgCC���^耮���V@�ßE8���k�������h4z��g�{���/"�b@� ��o����f͚�d��g�tJ�a8w7t2����!]Gx'�z�W��xBTTT����{%6�*���tcc㔦��EC�T\�ľv6O�ݻ;00�׺�����%@e�ٶ�7���yϚd2���477k�ǏP6�+�.ZLȓtz��NH9ƀN��F1���N{�#�?l0�/�Ѝ�|;6�^�����d,n�����x�:��-�T�v�Zmm=[�K�t�g�D���:�X�������E�3�<E��ݏ���!�iI��\��2��Cރ��z|�����c�9�gw�yg��)S�����T|�j�1|/g���ۢ��sB��J&�?"�a��jnn^����Ok/*)|�6��s�`@'��}4:�{ww�����ɕ�ƍ����O�$oll,F�[kѢEa��>�m���^sKHPI����n���vY�H$�eYo���|B���=G����P�@ 0?-�Z��N��v��n���OƉ��t�?�x����O������珲��;}��k׮=���B���I^�H�XʙD"�y� ˲���ګ�ӱ��s�����+++C:������X��p�n���+������fA/����~�|w��IB��J�y�P�T�^������!��K�sEmm���d�Vlo/�
��ĀN�[�W���0E�ݠ�C���@p�x���khhxa�KR +W��}���|X��@�j|7{��r�x<����w���y �&�<�D"�'N�؀Ч��� d4���P����\GC:[ҋ��[X���l_C��*����_���d�ڵBi�
��������X�"�[��?�W˳��ΕXʹ,�q�����B�a8�6tr%�%�!���	���XlD�L�<��ŋ�$�S�龱b�
�Y�w������#��b!W�wy7�t�'8�e�����8�O&�w��B������I��o�\�iI���ay���o �_�����o��$�P���˗KOO�P�*�9^�pw� .W�F�M�m녖�B�n��^`�H��(?��,�**�vXù������������(/���h��7r�������$�-{9��|͚5����r�P(4뛄��,�"����^�R=�eYVS������p�������\�	�ڒ�`�[������t���~��^{�����yl�;���F^朆/�P!�}UU�c���B����n|���Z�_�F�	�����7�B�y�s��éBÖs�a@'Op
/mAՁ�h����'�K��K��w7�����;إ��{^�/++��p4_WK$/[��fX�\(�L�{�P��m�����¹����F(���:y�b��qk#������������  ^��-�y~j�4�A�_Ǉ��;����B����R}��Rr�������~*ʔ��'����I��/��)NaƐ��G���p�~!~قV566���e�<����tM��|w�	���V*�d2� *y��FK��+BFAP������<��)�щ�ܟ��sҳ�MЗ"����mA?4�|�GxH;�s����5�W�Xת��~���c6�"�9�a��`�@�h�9�-����ގ���cul%]�?1��'9���9��k%*?_E8�S�_��+������6?�����\�5�q�(α,��B��@���Դ6?�������s�-Y�d)�\���K<��Ј83��:y�3p�ڵk�6i����U�7��p=NF���z�eٲe�Q\|G�4�	����b@'7Y[VV����P�hK�y�m�t��`�ʘ��V�sb@'���/���-����c�XA�7�T�f���.�e���]��;utt|�˄�H�҂��~r��[ZZ�	���Z��&�JY+�6�s�O��Z����N�E�f���sRW��^�hhhx'�Ý���ڥ]�72�O������*�*z1ζ����� �	���2�[�^]]=����.aY��s�:�FEE�`K�ϻ�w�pj4�C���3е��|0��8[���և���p���L���������}�������际��$�!����s�1���hww�ç��K��pn�t5cƌyhŊK�����圌�9˲����rT���)oQ 7X�H$�r���f�h�l��?���0s|�9��Nyy���g!���������"b�����@ �noo/�Su����+�����������
������!�K͗Щ�8�c
�9m:���t���'Sv����3���s�
������$�U}}}���B������;W�x��GD���jjj�
���a��\YY��m�DCa@'��Ry<��1�rco���z����+�ntvjn��\C�CǊ�L�����B������m�{`�,��Һ��nI�9��kZPjKzww�xL��oE�ѫ�Px��900p�>r#��*,�M����ǟ�,�=l�"�Ly4u3y��$Q__�5k��Ù�3�{�-�t�=�> �t���K�ψ�&N�8a6B�QBn��m����r!W�q׏��Ql� D�>z��'酗����B�P���'t*5�sJ:�x'��Rӊ�D"�
'e{ԨQ��}�&�	�.>iҤ{Z[[[�\!5�:��/<,�Y:��O����9�e�q����S�j}�h8�K�R���+�Z����t>�'�P�{��uN����ǍN��y!W(++{��Y.Df�G$�@�����e�Pw�);=?��y��[�ZI�9�D)k׮um8G�}b���_nnn6vq۶OG8��0x�!������2ޢE���}=����,���#�x�����}�ɤ��_+�t�_G�a@'���.��D"�uS����B��eXW���X__�����Ct4wt2J0���>�D�=iҤ=���5�O�� �ɮ�9�;�d]��u�D��%�X�<1�ԩS�-˺���Aǒ΍�-!�������8��?�{_2q���***���ϊ���;��|O�f��.�o���Yb(�'Z���`!?�?˲n���/	-�,�m�Ml�(D�_ȷ:;;WN�:���˗߄}��(vu��0�����k�*,_F8TUWWW��C�ݗtn���4pnt��;z�:��B��p��^�IǇB���>K<�]�is�W����k��d2yh"���*O�J?6?&�W;�r��/d�@ �8�W�A&H����&�{(�t�޳mێ`��(vu��0��o��k{;NZ�C8_ �B8����69��ϡ��3T���b�N�G�r=�r�������p�`0�8\�zEgj�t�evu��xng'J�ۺ����"�|6�7��jjj>����pN��~�[��2VKK˚�tk����8�}D4�!�}�On^HdWw���K.�ڮ�8���b(˲vA8��
QJII�W�o\�ǟ2�'��΀N��5v��g�h��m�Y75�X�vu��1��︬k��d2��D"�
lW�T���>�ƕ����655�2�cX~+DE200��&DC��bφ��Sc�l#®�1t��um��f͚#�.]�B
�v�=u���ڱ����X_&d�h4�жm�c	Q�<���hX(�����/�'����;m�{������7jԨcc���WP��/))yX�ixb��ƙ��8�O��[�}��iC�,�D�U�O��3�������|�E]���n��7�Kp(���'��hxc8`��Rӭ�"D��ȳ�H�!Ʈ��*--��:ҙ����|����x�����|�-]��>�H$3c���W���'��86k�(M0�l���O���i�"6�PA����iH����ƍ;�'������`P��zk�ZHgWwR����е�F����}{���rKT��{��e�ƙ����Ӷm�1�BT@"
�Fv�9�k�3e���ҷ�f�������Ů�ĀN�璮���b�3|�b(T�u�Q��d7!��3�\a@��z����U�`�=��u�� ���e�t�ַ��y$���;1�����k;NBW#��mr8�{Z�u'6����q�Ҁ�BT8�����A�ԃN@}c�L��Őή���o�<����xo���������X*D#�����P�@�K���>򞞞���u��f̘Q�L&���i�����Őή��ŀN�ez�v����b��ٶ}��U�r�ƙ	���8�bsg!ʿ� �-����Q���ˮUUU �����,���k!]/ZhH=z���0��'��k��s~�.���_	Q�����qg��΀Ny���!ϛ2e�8�S-������Ɩ[n���結��.���/��ɓ��~]<?��n����-�(��JyPRR�	g|/sq�K�����B������Z�b�a�`����ޭ��wwwK2��q�����B:���:y��]�u*�X,v��©������f���3*�Ϣ�ԩ�B�?-�D�5!���tvl�D�F��ƴ���筶�j0L����}�ϓή��ÀN�bx���DN3=�WUUM,--}'ح�(�t��˱���ZZZ���C�E����=dڴi[!�z�ױLs~�bŊ!{3jc��u>�|А�y����_�-��ܵ��x<~ޛ�g����2���&	Q�2w�eY�8`�9𝼈������]�D���a/�OD���Un��&�k0���-��ҝ��!]/��Ѯ�nƮ����N�ap��GF�u���\utt\�է���8`�AP�}Q[(?b�x|��+��!���g���EV�\�V���f�%��,�����-�ڒ���ή����N�`p���Ώjnn6��mȶ�bu��3���Q�����J6u��򊊊�����(&?h�I&u�Czyy�䃆tg�87�tvu�~��	�vm'�/�b17��C�өQq]0iҤ�[[[�U<��eYK�9A�r������]�����X�2jԨS��������Li�	���VC�����_#bWw�c@'�3�k������Εb8��ۅ�6Sq��q���*TTں�������jokkc���>c{zz�J&�'�8(��kx�zY����d�رy�ƭ��5�/[�̵!�]ݽ��\�Ю틂��g[[[��UWWO(--}�[
Q��2xrmm�#��|��Jusg@�\�c�L&~�ӣ�3����c�m��{�GB�u˗/��W �n�:��t�bWwo�J�f`��6��>�n�8�-˺��Bd�@2����޼G����I�����1cF��c��5��;���]�zu��א���kW�|�n�ҵ�ޭ��ݻ�ɵ�ھ'�/D"����m_���Y!2˞�7��x�PѠb</hM���P�t���煊J�G�>}�8�u�#��d�t��V��\rF�3f��èQ�/dsϼ	�^��w��0��+ص}5
�C�����pX�d����eUUU���綶GiCY�ڲ����B�ؗ������U�،3l�S�ohh8����0����5�k�O�Kχ����������U�͝]ݽ��&��a]���#c��?�l���k��\VYY�����P� P�Gt�	��^x����ƍ;��3p<��/�vk�������!Z��烶���www�����0���ֵ]o�==�<!.P[[�5V�`��M]D��Ú�����"BŲ �qB4r��X~F� f̘�I���4<���6ҁ���4����0v��d�����iO'g
vu�trӺ����$��(.������"D����BE�-���r�^�K�\Y�����q����q{&�V�߫�&�A��\�9���rKii�����~˾�2���-��U��~-�����P��X}^���+�e]��#�*����D9���y�����D<��ue��C�XC�4ҷ�z둄tm��ɛ�L���w޹~l<>��Yl�".î����N�aX������G�����vے�cٓӮ^{{{�eY�����-7n�SB9��n����O��)�*5jݬ��w�����!�C&O}��d2yݫ���tS�aѢE](�E����E���;����ބ�r�[��B�p�n���Jn�;�ᣱ�S��R�,DY�>t�{�F�c�	����ӣ�~�P�/Ľ�C��e˖vw&�/�>x���755�5�_���������.O�����+Ե������X,V��R&L�0vԨQ:(��N0DB��7����577s��G�%�42��>ӧO���S���1����:z{1iu��o"����6A��d<�Z4]h۶�y��,/�����j�#2�k��(�?�x��q�lY�u��Q�ܭ�����'TP(���G#�AEE�cB�k��F������Ѳ�&����C��{0�A���gvͼy����c��#�����"���~�d4�����{9&��G\'���,D�3&X�u#����
�E:?0Q��fϗ�5@ 8坶܎5��vm7�\Ж���{o)ʫ�[ZZ���k#��	���a�[�"���n���hum�?���8�|��	�wl����XW��	Q�p��Mh�v�y���ʎF?�.����aX����ۄ���'C�Ё�D�\�6�ߵ,��G�����{1�����~I,�%.������&lf4�)��P;Ƕ�p<�W� ��hE��U.D�iGPzV�#tz��ӧ�����!.:�
=�Z�B�@�8O|�7r��8�$��c�,3�%��ݽ��Hum�7��fz2��KC���Xl+D�S�}�b��*�����F��1!�������{X}}}'444|�|�����zz��cA�{�����H$2?W/������>�ӯ�����N���H�tm'��ʩ��eY^�"��q�����_*��΀N�b�v����7n����.��sZ��O&�Oڶ}0��+�z�h4چ����u��-�%���}��8�tmoG�~xgg�k�F8}��	��i�R,�
Gr�,,���9Fn��n��NB8�n��cHC^���k+,��n��\�t�ׯ�5O��]⒋-���>�dC�����8*�H��%B������"�� QP��GBD��Q��Cٲh�����,8Fo��N���8����O�q��x��Z�74N���Z����_�sq�-����.���(&tmǉ��(|_����q���;'?����n�ŭ��Q���.>�L���P.���s�L�V-CNH���/��E�Z�B�����`Ww�`@'cҵ��h4���p��*C��RO���Q�:�;��M�҄��[�x�_�q����XiW��x>6��Z/3qZ�iH,�!]/O�8񄊊
e�� ���:����O�i�veY�P1���K(7~�J�=MMMk��&�L����҃s�l�c�9&��ں�N���G���.�ھ)9�:NQ]]�a}}}��%�簫�;��!#е=��8���7᧋��I}GG�)X_#�7�������+S:�5y�x���}�W�y
���'\2�Z&r�[ZZZ-��JII����\Ů��sŎD�f@��nT(�Z�d�Rq����2�s��o���E�P�D"��>���
�о+��&ڜg�4�������V�Xq�ۧG˖���`HG��\<��xCx���z��~�{qvu7:�	]�Q���
�k�"����`��QM0<�˅�i�0��0p>�I\N|�Qر9�6~me���>wM���q����۶w�����n6~+TT��ڮW;����"�p�|f�"���G����477/�(n!ZwYY��Ņ�M��U 8u����*>���U�V���<�#���c@C�'����\�T4tm&��@\���nN�׋�s�����>�_�Gr��ܳhѢ.q	���������?)~?-4hŊn�V-ҵ��������B�З��ι>VǮ��b@��(v�v��������4(��w��ȭ��Z��Cp|�;a?-]�t�PΡ�\�V��to�u�]C8��lhh8!�����������Ȗ�m��L,{e�/�H$���'����$��\��n&~TE��ޏ����%�"8y��ٞBD�2~ԨQz/��B9�xu�g9��e�����+ƍw86OB9��&-_�\|x�o��Գ�GHc�/�F�,��n��]��ÀNg@����\���4>�������'N�x��M+�S��hh���#����'#��i�6K{6����Om��ɚ��O����5�K$?DHo��~b8vu7:�@�Gm��U-l���ڥ}���?�p�E��'�S(��g�
m�l1�{�e���d�D�	�Eoc��ꪔuӐ�Մ`0��]�E"��#y!�`5y��c֮]�*ֈ����,����ܵ=�E�r��'�\�X�����������P诜=�P�'D��F<_P�7�ӣ�3P���[��RZ��y��g5���cg�"J&�skjj�kkk���/^�a۶�O�Y����T0E�ھ�񨴿/.�p�X!D��*T�O��
��a:E�]�~��3�pn?���}L�8	�z����]�`�����������a������������>���b� ���?ñ��9Щ ��~.���"(�wxE���bu5*V��8�؂NCX�}��B�Bgz4s���H,eB����` �5o޼�6����?`�T�a�}}}���Q�N<��eY�`�@1�����>D���߅��Jq�=Q�5<ae���X_+�(C�QQ�
>犦��D>(�/�6mZ=B�	�"����G�k��ѣo{���?2e8>�~�ЦhC��&L��H���[+Q~���ױl+�cW��c@��+r��8�3�e�yi�ܝ����=T.�sӘ.��H!!���������Q+V�8���`�@����ʿ9�d�����r�0�~���6g�ѣG?RUUup{{��l_$�%�O��Cb�����^|�WE�ڮ�G�5��P��3��Fb˲>���B�����ɱ8�?����05�hO�mؒ��$�\O� k֬�o��Η���Nߺ��f�sݻ��������577g]�E}��̏ή���O���]���s���ඊ9��ǜ+�䪋��_8�_;����iӶ
���u,ӄҥ=o�����k��֚�B������Bi�>��io��h�B-�ש��:���cOl�)�cW��a@���n���ڎ���сo��u��BD�p *����kB�����чpw�H_D�{{a}b0���J�th+����-]x��J��P&�D=�6�_�Gޟ�455������L&u~t��gW��a@��ЃZ���2=я�
g1ض}>���BD9�J�v%<Q(
2��h4ږ��w�u�Pii�L�s��k2�GKۛX�B������Et`8���ƗүҞ�� �D"�Q�;�7���ս8�iS^�k;
ͳ[ZZZ�Ejkk�y] D�kǆB�'��Ј��Zή��������9S�N-���8X[�Q��p�:hz��݁��&���G�b�=൮�3p^Y��O�}�X,v����/�cW��c�H9W̮�8�\�B�6q����-����=s.W��+�Rq�Ј�r��4C�)������vhll�8V��5�T�'
�kpz4ԧnY�`A֣�o���K{� 4"(�G�~7��!��@��,|�{a��i�ս��)��ܵ�������A�{�ꅈ�崺���ZZZ�V8y�tvE&��p����>cQ�?*�L���� �t-�2[��?�s�⩁h��	|���#mCH�3��㜴,
}-<.�O�Ʈ��O�r��]ۓ((���ٹR\$���BD�4��c��V~���-�ԍ�ມ�Q�GC�8��x<�.�i���5Wgp;v���Ν��.��n~��5F(W��nB]nY4}<�H$O��W�{���]���r��]��2�ω�TUUM,--��Q���>"lA'�-�h4����k����/c��?,;qI��\�z�/��RG��eY�aB�����
�>���j6/PQQq����YƮ�ÀN9Q��o�w��N�%8Y���	p8��F����L&W�������Kj�>}��'t�#�c��G+J�dz�l466��;�R(_��;}���vo�=�'777����x����]���.�D����s���-�m�l|^�
*?ڊ�U��p�8�{����a�g�x�J�|,7������/�_�_����}�;
�S��ǫ���\�d��L��`�o���K�p���4b��ڎ��"������|"^*DTP:��eY�߸�.����@@ȟ����>��A��̹S{���+��M �}�!���(#SJKKﮯ�����g�d��~�S�as_1���:�H���ϟ8q����v3C8��`+��
m4�N��[���c�O酙��ʩB�I�^�4>����������~Cx?W!��*�}���o�g~\��0�'�O�s��������?U�"vm_���MMMk�E:;;/�j�QQ���:*?:�qR(#+�RF��p.�Y	,7���_~��1�m�3Q�}F���
�t�3}n<�O8����p��?�5���k;
���:�"�e�B�BD�4�V��>&��������?Z�=��Ƽb�.���>rӔ)S���;�� (���r���qs�}	�3}n,�=��%l�!cW��a@��8e���H$�(.
�*Q�ծ�A!�b��0�g���m*��e��%>��f>�-,7&���^}�Ռ+ �p�P����(3�ҟ��y�c���x
��ׄ]�}��&e��]�{Q`}M/q�g=Qn/DTt(?���������)�6�-���^lV���Z��u���755=/���:�g�(>��n���c��3yb"�x��6#�cW��c@���k;�_��k��x�g��N���'��j0��_��g��s˂V�L�:����.��������{477/���x�2�������`��{蔑"wm�ז[ni����2e�8���'J"��,ӑr/(RW �Q��	�����P;��y��-�����V��� ؗ>�f���K�P��7
����nt�eW���H)b�v��~�{�Ez{{��*,Dd�l����҆��1�CEE��*��ط�bߞ��{�6C�eZ=V�	��H˲.��g�<)�H��/���s1���oJ^�"����x<���
�#�:Q��T�	zFP�Z-�>�������c\7����������-�>�S|Go�>;'�'i�Ѯ�����=#��=w�)-��ڎ�����{��Huu���W�̅������oG"��҂2m�
�����ţt����y��=��\l�>ʁB&��(���Y����V�O�ޣ�p���~��o�dW���Gi)b�v���uvv�A�f�d2�ӯl'Dd��(׎��*��hw!�3f�x�|,7��|�/��x�eY��.r���`pN(��H$���F��m�Zl�.�cW��c@�a�k;��ǟ��D"O`�Smmm����>�x!"�������4m9/++�X��p'��7o�k�Q�@�w������(�n�J��������j1���:mV�Gm_ .���W��O�:�{|����{N�gz$~�����x�Ͳ�]����t���<�z��d��c{6����7���O	ǻq������{f���E�u���6oñ����S��*b�v�s^kk������R[[�u2�<�g`i"*6��\�a� q�ݳ\�z��r��[��+�,������s���ӫjjj�er?z,�!]{e~AǮ��c@�!�k{
�Y�A���o����I�umU?�W'*{3�s��J��������p�s���8��cǎ��ܹs�Vi)�������[m�@��u޴o���?���>_Ʈ��c@�M*r���@ ��U���!����.���8�_��9,A!�B����y��m��^��x��Fn�k׮�~����Czk��
��N�/��;�>���-���b<�Wb8vu�?-ڤbvm��R�n�F���]&M�T��߯]nu�	��;=�Ї�
![�=���+p��g���+O���8,�m�:|������7�}��ŞM�9[m��o��������]�3ǀNQ̮�(�:���.K�w�.�Q��^���LD.wX(�6�H�+4$���J���z>�ݬ���[.\�)W�Ų��� �B^�r�ĉwNwZ������~��]�3ǀNR��zu�---˄�z�9eʔ������$|G{�Zy �9ѯ[н����۱��h�655�Kh=۶w��GB^SWQQ�]ֿ������eݏr�p1��g��}H�Gm�g,�M�#tj���r;&�I�֤�7o+D�+'�p�=����ۓ�<������堍�]�Ȯæ��hD�϶�.�L�O��A���4�y�]��ǀN�y�v������gX�H�M�Ϋ�����e�tm�	�Y!�T�vB�-vC@Ū�Ŵ��z�r+B�_^}�ՈАP>���ӳz�vu�[UU������yꄋ-˺e�b8vuO:2�k�5�h�I(m---k��U���3��u� D���X82�8͚��=�X]N��q��Y>o޼�xq~x555���y�䲲����~�O@���8�N�z����N��O�y���8�\$��x<��Ϋ���iww�������@a�:Q�N@%�G8~�B���3KyGFn�`�qο��_~O(-����ݘ)'�m���t{s�������]��9P���ݵ]/\����.4b����*1G�P(�����{Չ2BEx_�Ӟ��O؂��z^�Jr��w�njjzU(c(���Q�/4�]��f�t/#�ߍ��	<�3b8�����/44t�ӃD�d��UUUʹD"�U�(��&q�5o��0���k�x��l����͛�Z(+�Ph7��ٵ�f pk#���}B0�v2�\ .�w쉵y���_�l9O�.Gjͯ!Z�O�2^�hS�����f�ءp�5o�������mXn�����	|\e���ߜ�I�=EZ�fδi�V:���_��z�媨W���uAq��(^pd�ʾ��M�a�m�Y�$�t�6s��{�IIK����d�9������3əI��9�����@�����X�'3��*��Gŝ5���nݺ-���$¶m_��O\����tS"��UP1C��z?=�;_ۧ�����f����U���1�������d�Ymƌ׮^�z�?���t:}�n^&�C�����o�|7@�3�E@�dI;����(-3��n.5����H˲>��k���A@�2��	��Ƅ�.g&�+Q����boڴ�KPRzm>V�N����s?�p������g�����h4z���$p-:&��8.H�RO
&��6��%K�|��������^^*���q�.=&fm޼�[0�ۻ�	����|�{ˣ�Wccc���ͽ�L����8��vYL��fV��~.���G�D@�d��(�*� r�^.\�`������T��5������[��4A�6�L�^3f�(����zp��)S����v	�*�N�FWx��H���qf����==Ws�r):&��XV�z��XeJ4]��ͧ�L*��ƍ�N�@���T(������ޮ��5�L�7�ׯ�$���~H7�@?�3g��m۶��Y*�����/�������{���񸙅�[���?0��}E!�?���y|��s�����=w����f�7�V_����/���.���ox�yuuuf��o峳��Ķ�k����QQz�8-�O�P=4����,�r�6 �;�s��O�RPw�2�t:mf�=W0���B555�eI-Wd2��mذ�UPq�X,���˵:K��}EC��Ds>;�~��o���W!����J�Ry�?����ֶN7�,^�������k���{��]f�;�9t�>}�H_��rC6���%KnY�re^P�<:;;�WX�c3�����?
xη��]KI�n@e�Q1�@�[�`}T�زeK�nΌ�b�ttt�'7���x˫l�^�o���]fʔ)���q�7"�k׮��`�E�ѷ��k��.<�����|v�k�?�v����.A@GEhx�?�_'�m��f�)���_�}�p~�W��3+O렻��q?��Z�֯6��z��k=eT��ŋӿ�%jȓ�������ܤ���}O�}O�jX�
4�Qz2����r��OZ�h��3��)Z7�^ w��Ї��]dʔ)[-�2�|^�iӦ=�����jhh��n�	��Wڶm�G�2��̈́��H�B}�}V�
tT�]�dr��7Z[[[t�K��ooo�'d��=[ wza4�i#g���������^��SO̫���og���(��o~�lٲ���B(�Q&���V�
�e�������ܼS7��b��ttt�[�&��� �c���}@w'k�M�����T=�Ϋ���XC�(����n�#��$����[m���V�)�zt��-�x|���r��_c�6J^���/jy�>
��~���Su�����Aw}��O&�W�Rcc�"�q�$\11�]�d�%�7o��g�P(tF:���VT5:�)kY�i���f&(�϶���Z>%�B������F��%>��/�I�0龜�R�,��M���/Z=T��9����T�~7��[ZZvD��s��xAU#�����M<O"���n�4���B!���)s�Rڨ6���:�=�UO�W����kUJ�#�տ�Q������D~�T�����{nmm헅������{�1��[�n��鍍�g��i3[��O��T�w�b���n��+zu����T%۶�2��ẗ3Z��|v�����F��6��U�����e2��$@�ZZZzus�^h��`��wX�e��[!@�xAgg�1��M|�uЫ��}��si���h8�n���>���L��Z>;��֞�����^��E@G98�`�O�P��}�7���P��Z��:�(>�Bz���dg]]ݙ����se��� �g�W�S����lV��@�z����*�Qrf򓶶����܄rǙ��8�Y�ZX�	��=˖-�l�k�z�JY����Җ�"����V���L4lD�kg�R�'��?����oz�g�%��O�QRC3����(m�����m� �7�������^t�A�Z�ĥ��bfl�k��B�+��5����l�f���yZ�����Qj71s;�%�J��͉.<\����?�udQy~�Nz�f�_ՒT�@ `E"������j�>#�H�#��kjj~����E����QR����r�P��A����w�1=ꨔ��q���+^<cƌ��޽[PU��L&W������ͻ�+�5�?��ι^�_j�4AU!����J�R�P!���I�h�,ݞ��f�'ܣ�����6���*��׾vJ��zl���c�� �Wu1��Z���s�n� @����H$���t���j�.�t�ҏ��x�I7�נ�L� ���ʲ�����!}8c�s�X�:�&�fA����u�hBL=]~���䳳�?����zn���j�Q*�A~� �hXP_��@z� e� 3��g�4���x��p8|����[�+	�Uo[MM�OUc���qs�p�&�	��m�G���q�s���9�����Z�����1�Z�e��)@i�a����q13�Պ+ެ��5� 4�\C��i�RAU���k�zs�Vk�\s~��;��9�4�_�����*�Q
Mzl�uFcT�T*�J�rm8�O�?�/-�Dr��]�_��WG���/_���}��U�Q=�](�
�H��7ku� ��x۶�-�H�=��3�����0��*�1a�`�Y�V�T�yM,���������`��}��e˖��a�K�.��5kֻ�z����8Kjp,�����L:�/�}�.�P]N���|vL�ROF�ћ���W�;ʋ���j����R�*�v�Z�,�אrUOO�i��ڟa�W�cǎ�t{�T���:�p˲N�p�I}x��Z&��_�����kU�s�T�����[wj�}Q�ޢ���x��|v��ӂ�^蘨���0ܭ��y�n�n���uk֩}� E�ƹ�^u=��Ҡ�aޟ�r���6�;�N��^�{��`�͛7on8�C�Q�T�^�c�����@�>�u�IE@�D������Pni�w444�S��&�/�@ڐ9�onn���m�S4�Y[[��@���آ'�s~�J��I�׍C5�߭�Pݎ����u�׎3�Mt�`R�Q4m^��ֶ] ���˖-��������GZf�����3���J�P/�s�i�U�}��i�*�=��Ϻ���L�H$�=�Vi�e��Yi������~��ǟ��K����be�Q�+< w�ƹ,�.�N�T0r���е���1z�5C�џ9�������d������z=�̄p��=�η�L����Z��L:����5mmm[����6ݼM��I����`��n�@:�~���	�0����}pC2�t�~^�;&�=�1\F�!���=���8�E�e��iM:���9x�6�/[�x��g�Ï
0�Y������D_�h�| 'h�>|��zơ��}�u��Y�dɬ\8_!��9�H$�m�<8޾�Tj��{�>竂IA@G1����a[�l���I�X��[�70:�荍��r���l6�F�r]��}q�6������~�9\O�/ߐ}תq9�s^0��V����!�bp�9|�L"�!j���3�᧵Х���[?��05�f�ht����~X�+�טm��ߩ£�s&��p�*����,���M��hn��m���W�Gi�Q�muuu�GZZZv��H$r�6������P}�^F�ǯ���n``����9I�MB��ׅ*}�A6��jGG�A�����B8�w���M��ֽs��>)h � z`��Yd�W�d����/�jC�]�4d�z�m�G�y�c��}�p� ��[�9| >	.\8�q3[;�^��h4��x<�y������Q�G*���B�����c[�nݦ�r3��F����?�=��9s�L������G>���p
g��_T\.���s�9���w���䳳^�����E��"�#oz��5�H$��L�[�u�>\.�H�mۗhc�L���4(�^o���!��ŋ���N��\ ������Z�#mӧ���*��LXr���(į�~�T�ImH�:�|W��l�>����� }u��Ԝ.�����y�tz�V_&��՚�-t���v�ߣa��Z���b���cz�� �����h4z���E,* P�on޼�[P1Q˲�����@ p������ݶ7&�q~����Ul*����h��U�u��Q���{�,Y������� 
�`*��LP1����4|�m��Ǵ`0�ݞ6ގf��m��j��	*���|�����L�W x$1�4���F  ?��/�ax�444�8�s� ��h{勍���䖒��$��^!t��L����^�q}n4�_�Wk}� ��~�H$T�mۯ�pn&��+�?�J��f6�3��q֬?www�B8^*���qiȸP $��]�t�}}}�1t� �(��K��F�j�h9T �JCC�y�Tj�X;555��UJ��A��1�'��� knnީ���E�d��R�`�@`���"������5������w}�Vg���e}R��QƤ���q��������^�.�~8`b���.\�63�}� ��X��+m�^m��Tj�������wl��u`ȩ�X�wk׮k����-�H�.=���c��� �0���kll���isL/ 0�7Y����+���7[[[�
&L����B�8����eV��r�5�_�z�q�¨������ ?f�E���+��{�~�%( �|f�G3��{5X�(�L�L��AQ�w�yݜ+�F��oj���F͆B����i3qt��l���������F7j�
��@ `dӴ��D>���D��7%�Y��{eCCÛu{�X;�����1�R�'ʆ��Ѵ����- �"�߮�#-�2B�� ��0��i��w555�ټys�`L��
����Z�� �2f����/��^���ˈ����w�G �M*�J,]��������8�I �3��|N��D"_L&��(���wt��c>" ��۶_�H$�1�Nz�yP�{R�/�#2] �]sss�n>������{��X4�8��k���5��a���khh����vP3��k���x;j[�2��eA@�HN�RO
���>}����nڱc�d2�`l�@>Q�Gk =Y��7
d��������y� (�;����~c���t�#a�۲ �c$,�T��ŋo۲eK�C�������_ `�,˺޶�������յ[|*�.�pq�V_. ��s�t���vJ$)=���[%G@��������V�\���b������eϞ=� ��rrmm�.�X[[�}�3��><�m0Q�,Y��'�MF.�㎀^t@�[Y���L��`0�-s�����z��s�N�t yX�8�=�m�8�L��/����U��Yˡ�f|Z�?k'm�\oY��3]PRt����$ٰaCs,3�_G��uuu��]̐w�K�s?��#���/^��-[�t������@ `F�M %��f��lٲ󚚚F��.�J�m���!AI�1\�^�n �F/�������a9�C�L700  ��c�|�v���w��s�� �֠��8w��\iY����D"�# &M:��FC��Z�9�5���t3ܽ��C@^"�x^m������ϲ�WF���5��X���������:w̞=������*(:���R L�M�6��b�X���ߛ9s��}�w��t �0�4оv�ܹu�,�B�m�J���r{�o�����v0C�u��j����!�cȿ���j0�,˺�q�O����S�{7C�u�<���������w�����͛7oZ$�*��/ *B����=�ϕ�@��^Bt��/z����{����bOh��#}���۷3y�|�<�N?b�������E/^|���n�jL T�[�2�mmm���C*�Z�Dڵ�@Ptr�P5��%�l��Ѿofw�/���O  f)�ۣ��g���%��o]b����RPi�_����%m���V�((	:�m�T�U��^���t:m&Au�b3yܬY��I߻w� @j�A}�6�O&�ߪ���#�ȫ��Z�# &�G��Y�_��瑫�X%��o��C=���n��	c�ǯ̘1cp�8ӛ y:U��?����+Uƶ�����
�N �iJ04=�?m���$�Ո`��`x;P��qzq6�=A�0eʔ����q 
pB:��u�ҥ'477W�'|�͐�s�X`�i[俗-[v���}��g���^��Lfx����L�>��]�vm���|�g�8 Excoo�����{{GGG�d�C*����o�j��������|�4�_��0��>��_�T�իW�W�Xq�����3y�^�������~�<,��ڶ��D"����,]������R�~@ T�fɵQ���*�<��&���s��^ T-�q.֋b��0�����ˮ]����G  ���MC�[5����?X�!��N�]G�����h4zt<_3����o����	!����P(�Z T�u��=�bŊ����B�gB�̙3�K7A �`�1������T*��?pѢE��1b�D T5m��^�5c|�Z�����j����r���!S�N\����N�q�猻���q�x|m9���z~�Q�o�	 78A��%zn�<�7��qGoo���!(�Ǵ�~� �z}}}W��ՙ���|}����� O��F���!=���ܬ�<M ��YY��Z�2�7������q��?�/(ݿ��p�����Դ;��Y�/�5��@�LH�c�ǵ���+�k8���_i5( \E���;w�����v���uZ�@@������3��0w˲>>��`�w ����l�>&�H<:��-��}�|_ �լ����t�������m��șE��So�e�����b�'e�)��{�nٻw� �8ղ�����T��b_d޼y�4��%��- \�q��k{��&�ikk�n���ZeU�"�}J�����u��z��d��cB��3{ԙ�@�X�u����iH���h4� �e]c����R=�Y�w�������^$�?=�H$���d2�KC���D�m�����- 0���/n�m�چx6�'����͍Z��34�AF�7k���(t�f��
 �ٸqc*�ݮշ��5��@^��憆�cR�Ը��h8�n��2S x�;-Z�����r�7��?��o��BA��>�����+����l��14û	��tZ `��,�
=�O�E�.	���/��,i	 /�2��gu������,�A�����8�}��zzzn���ۦ�9�|]Ӌ>{�������`�D"f��5��Q����V?' ��S���;���c��3��Ћ@@��{�D� p������˗_��௔�����&��ܹ�|  0�������x��C_�3g��fH{IG� �Z�����t{������K�׫�:AA����v��4H�a�%�CfΜ9����# 0=�����d2y�����άs� �s;����U�m�oZ}�� t�q�6�j�<�H����	+��3�O�.�P������П�n�����Kz� Wx�Y�!�H<z�7���*���D@�=@ZS��S����w�n��3���2l��`f��˴�����-�9=�?:���J�/(�G����v�;���gZ������H}}=˰-p�?�\��d~�����X;�R�M�H���z�G��,���k�v�b�k���r�,�a ��z5K\�m��ZZZZ�y��Հ~w �� ot�p��W x���E���`6  |���-g%��T�O�v�]�!����zplL$� �X�~���˗o��J�<s?��nBz__߈�d�Y�~3  \o���C��O[ZZ:�}}����+�'ǹG x�:����L�W�g��=k�,�V����/��  �����זe���ֶ}�/f��۶ݢ�FA^���Z xN(�(�N���`�~f.������w��Q  �]B����~A*��[��^��ӂ���!S[[�F x�C=���b�������~衇&�m��_�b����	  �cn��e(�}KKKo9~��=����D���o޼�[ x�Y]/|����~������������  �b��~�J���m��?H��=������퀇���������3vh���z���� p�@ p&�9S������[�l�m�Y�K�"���=�������/_~�^t?_ɟk>׋��  T3G�-Z~���>��l6{��S�y �{_����>�uh�X@7˩�ܹ�T�  ��dƕ_��d~�����d�C,�Z�m�O�E@��۶m�% <mݺu��b�Z=�?o���º�  T�=Z��8��R�TB���A䅀�} ��X*����e��R��  &h��_k�U2�|F�H"�h�m{�V��D@��@ � �����+4<��պr��]�� @i�rn��0/����O0&��e2z��x���]�b���l���{��ah;  �ah��?��g3̝�>���W�}' *�q���@Yz&��  `�L�Ri��m�5�e	�F@�0s�
 _Y�~��˗/�k5Z��6C����  ���J������#�B���"��n�N����a��0���N,�T��+�����J__�  ��2��"m��<�J��Ŵ���m{�V��`Ttt��2��E�`�;Z-�82m01  �ե�Z�K$ϊw<,�1н�w֬Y��lذ�5�ݣ�7���̒j&� ��۬�Z��`�#��f	��нk}SSS� �%� ���&�M0g�s  ��,�|v2�4��x�S�p8�������]k�o��������|_?��ٽ{7� P-��u�������F"��@ p�`Dt��}� �x�'�]�����n39  ()3�˕�^����g4��Y�����Q�`����^ /֋���s  Jj���-�:���m��}to��ǟ ���#�<��6i���>����e�  (�u�l��T*�'�r����1
�7m��`�Kͽm�>��� �����nq�\��1�������v �,˺,���T���>���  (�������`Έ�$��gl�Nh�<݃� �������,_��&=/�G�ϡ� ��qya�-x��=��g&��M^��s  �����a��_^ �]m��ō���==�d�	��ŋ߶e˖����ݻW  ���/�`����I0"���'���p+W���b�˵�?c�gzΙ� �Quk�4
�����UP4�,#"�{O� �A2����`�[Zu��={�  x�Z~�8��T��f%�L&7G"3��t����f 8Ȇ�W�X�F�o���t��s  �3��d2�LZ�i{ım�t,�Zp ��Ѓ`D��\���:�� 0;�Zy�^3��<!(�=o��7� t�ѓ	�����5�p�\���u=oHoo�  �cf���:yYKK��`��нeg{{����ٶ�^�,��Z-S�=6������@`��K6������su�i��9�����R��ڣe��T����}��ߥ_K{����_ۡ_�{<��e0ܡ�&k�����ݖe9����P(��w��ئM���b��Z���p��_ �g��]w���=�L>(�4n��[�����M��m���X/=��}9���l��Z!��F��֡����6��>̗wiIۚ�/̢�{������[}�W�g��kݺ�m�~m�� �ɘ�{����� JE�S��쀀���#  ��V-���_oݺu�`R���?�"�{K�����2#��}�7����v(�m��M���� vju{�<;��=��o�3��.a���ӕJ��%�0?���X�	���<֋��q  x����׶չ�>��e�'_GGG��o����н%�a"Sn43W���{��z���gz����x�^����ڵ��d2�`0ؚH$:�l�_0�����LSgr8 �ǙQ��k�U[[C����]��6����=DC�y�J��qCr��&���ۏD"ZR�=3�A����۴����Z[[�
<C������;�6=�  x��c���̥Z� �?+�J�wzR7�a�200�t���q��^��֔�����d���?�+O�O�ן���y��N�硇��b�������p  ��6ʍ�]�*O	@@����[��V#C�Q(3�>�+����=�Ng4����ǵ�ӯ?���gI~UM0����   ���5�o]�H$����8O�6%�C@���{��W7��@�Z���C��E"��կ�C��^��.�J=Ƅ,գ��3�g(  \"�������Eǀ;i8Rp �w�;����1��V����No�s��ެ_[g�������<����'��)  ����_7��Ommm���L&�hѴk������%�c2�	�ϕ������޽�7��Z�nJ"�(佌"h�&��	  �C�Jm;�>�J�xF6�5�K������ޑW�6�-m��	��T-�ɕ/�/�I�[ߧ��	۬Ujz������%����< �z9�xP��i{�r��Q�wޢgz�;���i�������ғ���=67i����LBgz�ԋ��z��~�	����C �Fz�2˽^��d.iooox���[��="�Ճ�����1)}Y�|҄v�]Z�_O�k��}�Db��G=�H$� �ztk��q�˘��L@���9to����֑ώ�P�&�&����jy����c��8�D�эZ�������ݻy��n��ض�:�=�  &W��;��t��?3�ݿ�￙���7���Ic���A��x�n_g���>7�<���ӯ��d2�lݺu��,�wA �$2���1�N��k3�`0� ��н!��sB�P�̞x�Y�}p�x�'����o���k��L<��������>�)  T�Y�����w�^�0L&�٢����A�'�I/���t�t���\\�M{R�k��Y���~�x.�����
  �g&x5����H$�+	�dno�D"]�&;L@@�y�`0f	0(��Cz<|�|h��N��k��{��� �|C��+4���`���tC@�'҃��d�AF`>�5ˏi��\�V���=�{a������ %d&v[�ז��Zys*�ʻM
����^��;����@>��`0x�=���[�J\���a���  &ƬY}�� ����֮���L��pd��>tH��yt�q�A���v���LE�wk^F�X0|��[k ����r�^�̈�[�0g*O�(�At�K���o�wgzЁ�1a�d3K�n���8f���}}}�V[��^��$  �/�e��Uz][5u��5���}�WJ0���~)mx���Y�C�G�����:J��������Z��F�5n�ϟ���k�L򿑀 IF�_��:v���X��ѱG��"���]NO��k��3IPvf��X��������h��������U�3gΜuuuG	  ���߯ץ��]xW<V��E@�!��_A�k�!���7]��cu{��3���[[[�M����o��� �?��k�F�ͨ.��h"����$�ɎH$��}��F@w9=�v����C���n��L���˾	��2e�����O��� ���<������@{{��z}�P��{T�C�Z] >G@w9=�v��eYAzЁ�b�U�����z{{��j���6w$���g� �E{�z�A��LyMMͽ[�l)�mT3̝�.p�B{�e_ P��jy��o14�wi��o��ܤۛ4�t��>'�D� �ۙ^�'���ֲ���L��\�xޓU��ք��zzR.�SRݟ���\3^s��h`� ��Fu�C �6f~3��:=��g9�����Z�܊K@w�`0X��R���2�0;��{���x�-�J�~�6�s���7<���M�����m�t	�n�'񂆸g�� �u�3�k9�m̙���~���8����~MSSS��� PM�}0�J�K <# ��\v֬Y�
|C��z�)ʿ��ݽ7�>��� �,-Z6�yy��w\�Z�802=N�1�5��5=d�<�R��_��[{ P~f>�f��3���ǅ�q� �L�_fD���ݭ��s���   ���-m�.>VSS�����' ���h	���s�    �/
�kkk�" ʁ�.t��Q�s7  p 39գZ�b&�ܤ���Tj� ��)S�l����#��[1=���  �2s��S��+N�8P�m"�m����1��Й$  ���m�{���X0|<�?�uG T+3̝�w�L1C��>  ^��r�ƛ�iںuk����U��v=v���.fYֳ�>�q   ����~b۶m���iV��qL@w����=�  �c���L�ۣ����N�ߎK@w7:  �=m�/:�z���]�q��"��  ��h�~� p=z�	讦o�=E<'�ew  �!ڶ�# \�t�����q2��  �Ĳ�C��iNٕ�n�o�E<'#   B:�z,��#���eYE�,C� ��Ѓx =�tW�70C� ��5T��F:��Uv�=��]lڴiq ��i$��֚5�%
��[rp�)��H�Hoo/��Bߗ����+>G@w�LSSS�Ob�; `<&�O�6M�N�:G}ʔ)�eƌ���#{��1� T�!��	j����������ݽ
�=7� �	�ӧO�b��9��&��ܹs�G���E�f�v� p�l6�'>G@w)}��� �	�3g��^�ך5k����Ȯ]�������!��F@'��Y��q ����~0P���I7a���s�A��: 3=�$qp�b�@7� 8��9/u8bz�����'('m؏?i���׋���B����R�����!� ���,����}�}}}���eD:�r�p�I��T�,�q gf^��K��3�0�e��-K ���A�#��WQ�!� �!��RC	��1��MO:Pھ�w��&���>����^E]�� R��a> ������^��~;ݥ��l���  3��\Í����K&�����]�؞p�xe�>l ����4��M���= \���^�~J\���  o��el��%��� p9˲|�]j���~:  @5c�8 ^@@w�b�A��� ��&k>��o��!���{Ճ�2z� fN_�\x�ԩS#�i ��cǎl�W�6t�*j1sm�L��@ ��a�7�ٕ�8t�g��m��M ��Hj.���m۶mo$  z{{M�����E�F�{����Օ+W2L�k�]*�͆�|�c�v�VY� |n�޽tx�	�}AKK�����J��@@w�b{�s�Dqt �9s?xOO�L�2��?kϞ=����f�:�ZӦM�})N�K�h";3Q\�  |o׮]R[[[�{�M07(�@`��<�[�t�盛�������Ԅ�E��{M� ���ֺ�����~x�)��o߾}Җu�?���~֬Yf�����B��9�{M�%�Z ����o��)yH
�mG�4�s'�.��r��?�%��=� ��1!��g���3gJ)��{M�'��������y��6l�! \E�5ϾC@w��ރ �L�6=�ӦM�ݽ��t��a�773�g֎
9��.
�W�	 W�c�!�W�F�D޼�� FdB��ݻ���ݔ|z3����`�I1�$��)t�uL@�2�.5�5q�A ��q���pSL@���ܚ^u���M1C�M8g(;&��"i�MGqD�ƍS�5�ZRS�UE܀��R�@�6��Ӄ ���z�@��Ao�B�����qj����5U���lqc@�A  �aFq�����N@\D�a�A���D꤈�p}���r   ���;wʮ]�oŨ�����:��9�U�z��~����+hF�^��>݈��b��a�t}��   1�f�BSL`7A=�9o޼����� Uϲ�Y&��[����~�d
  x�	���px�m��~�6�olkk[' ����st�NQ���iG�!�  ��r�Mq���[�~��o�?��֮];  �B �]�Z��b��C   ��Q�-��bgg��h�.�7���^�y��n0i�A'���D:C�  �m����������������T*� ez�I��Vz�(�&:  �󄴍�:ݾβ���m�q�ߨ�������,��f�����]L���󼚚���tZ   0��Mq监H$��L2w}0�[KKK� (���stw+*�+�A  ȟ>��f?�N�{�Ѩ�Q_��dnhooB �
=�7�]̓Z[[wF"G��j
  ��M�p~�n��gض�E��Ds555wһL=��
Et��8z1yF�s   �X�ɖe�<�w]���T�IP����;���   �R�߻�������S������' ���9��M$�w	   �i�zoo��h4����2��u���m`����:�L�#��[QC��8t��  @�Lv�YƭI���n��������_ 8�|B@w��{���O:  ��Yf���N����]_eY֪x<��u��C��n��mB��>  @U�߻�8�D"�.��M6wk*�J�}t!����X,^�v�@�O4C�   �h���N�퉖ee�px}|g �s```MGG�<F��s�@$������efbo/���  ���)���v{�n����7ɾ��͐���D� �G��]OO�󥈀^�s   0�L�}�)ο���ԩSװ�\��.t��d2�y^0L��i  ���{{{�h`�_���~��ٳ�2C<�@߯�ŝ��z�&.*����vF"�^��	   �b��7E�twwh`T����
��kkk�.@��\�@@@w������;�d���   ^��z�M/eFۀO����9x��{R�T\���  ����T����ɘ�  �A-��N6C�5��S?���Z�5k�F��cЃ.t/(j����>�}   ���\��y���m&�{Zr���`p]<<�@(�$�H$2��G� ��\�C�s�e8   f2��^v�qD��6����i�dY�F�-�v����L�cP@@w;='�UB ��S�ȺGYO��� @a�hyG�H.����^W�2ou�Qۦ��.��{ t�a��={��|o�0��|ֳ��"�������
 �J����{�eYw�����oض�	�,  &f�^k^�[S$��ڛ��Oh�l��O���=����%p���F��S}��#fi�ٷN�!Շo_��Y��п��~dD0���~5��6CBڥ@�P�I�B<c�6����*����@�~�a�� P!��T���vS����x�~�Y���݄���8�ZO��;�2�������h�����i�ޟ����`p��j����w^�[��v�~}�n���}�^k^���_�f�W��L�C@��L&�H��---z�4�`� nc>]3C
M/������m�ڵ�<Q��Z/��  �e�ߊ\�C�N�H$b&�����Vm׭	�;�Vﯛ��s��=�����kU��d�kx���נ�z=�L�������3;�5��/Ǆg���c�ƽ	�3rAz0t��fj1����w8��~0���C�{��=>��X��kS!��s�W�C@� =1Eu�@�OR�k@�3��l�b֬�����m۶�*�R��S� zT��  ���&f-�ֆ�Ǒ��i�����Л�	�Nn�Ѳs������'Z_/����;�L��}a�yL�~��L/�Tٷ�t�o
�C��m!=���v+(�믮Q0���zp.�����At�:��o�c�v�pݝH$�-���]��K@ x�P@>d�ojKr����OtE@�!�{����Z�hp�?���'�J-?�}��   J��^$�h��耮m�'���T[��2�����֮��ݕ���7۶�Z�o  ���I&�[��Y�#Sts�`�&�7Ё�z�,���ǹC/`������B=� @)=n���wg3�u0$��н�耞J��mo��|P��Q��m��fΜ�����mZ�#   %P����>��ϛ7onGGGW1O�f����.P*f��[��nzѹ���m�T�����h4z��;�,   �Q��L���G��־H7Et˲у��L��Zn���x<~�%W�L&�{�7� @Ih�B�w��[n�C@�=���"��� (�^-wk�Q�͉D"%.�J���m�Aa�E  P�`pc!�����ޱ��'�A�p:�6�}|t�mp�u�qn�:u����}��:  ��m���[|���="�;��綴��m�Y�E��Qf2�5�@��7&�ɧŃ;찫;;;�ը   I3I���V$)��ы��1�p}����X�mz�����,�83�|4��^T�  �"ijS!�k�c�����#�{��'P��v�|�j-���6�s�noJ�RO�8r��������}W��  �8t�/���S,X�m��'��ՙLF ����4�ߨ�Z�]/Ķm�vٶ}�V�.   E��U�C�_�e��н�Q/*����q��V_,�7�h�Kˍ�p��-[�t
�8�y�e}I�a  (L�ܹs�*�	��!�{H04}U���9H�1����.s?y�_���vF�J��m_�Տ  @�����צ��1�� t��l��_��gp�v-��d2�&��r�F,������T   O����C@?�C4\O(����{��0�Í���K&��s{{��~��T����m�J�~X   �W�q��8D7s �{��'�䎎�.=Ṕu� ��̷p�eY�������0RJ?���  �W��/�v��@4���>�����h�!��Zm��g}��YC�ZAY$�ڶ}�V?)   ��j�~��'��Wп�|t��s/:��۴|[����z�+�q����LW+   ckmkk�^�s^!x���a���D"�@$yV��0y�	�&�״��ߪ�<-��T*�m�B�~N   ƶ��'h��!�{�D'�33^G�ѻt{� �գ�ߛ2��gϞ}{SSS�`R����\�	�N  ��е��D"/<�{&�sn�B@G%���6�q�h�y<�T�{�۶}�VO  �QX�UP@����l6;S�<t��7��t�Y�9ޚN�Yn��������%[�l�T��M/��W	  �4;l(dm[p��(��S�F_��Ǌ}����}�z�%@����Ӳ�?9�si2�,hL�D"��D��ի  ���R�Կ
|������A�Lf�L ����է�N}?]6o޼�֮]; p�d2�Ҷ��j��  p��'�fp݃��	�M�5L@���SE�?O��|}]�H$����M��O��|P   r��@@/!�����!ȶmo��b�ӯ��3������w�^���9ac4�P���  @N��566�cTt����B];Z_�}�/0�f-H��mݺu�������ާ�  �X_��ڞX!LF=*�7M�F�/��܇N@�H��h��	���Tj5�����7�V   ���A���W	FE@��RL�L&�D"3#��K�����<.����ƺt:m�C��   <�����+�"�{T�&��D�ћu�1���{�U�S��B�oii�!���4^%L�  ��@�P�1�=���\����_i8?'�J��|`#�H$r����hu�   ��ܵmќ�@0*�G��rD)&���������[��~a�'��q��j0@�;K�,�����;=�|P `��4%z> ��� β�S����]�l�>B��;ٯ���/�^��I���*�|;�?"�%=o��[���˟ (	�9�M��-[�t������az �V&�s�s�n�f��������a�/�{ �D�$pgk	  ��*�9�>��i�z�nΛ��v�awvvv>#�}�9�`�]����ŋ�p~�V�"   �)����NK�1�����kK�:k׮�m�:�~R��,��mmm�	|-��{6�5�|�   䯠􆆆��Z����mQ3SbRM�4�]�8���ƾ�J���e�_[�timoo��Z=U�%   ����yB 8Z0.���^��}�x<~�f�.���ѳZ�
�B綴��
|Ͷ�1sK)   ��Ph�2�;�I#�G@�8˲�}��f�h4j�����M���N����$�C�{�ߣ����  @q
� N����"�{\n&�R���q#��ǟ5�����U�{�!�gi��  01����ظH7�`\t�;���aj*��;�J&��F"�v�.T�����������!�f$�  0A�`��B�O�ӯ䅀�}akf��]}�l6�hC�/Z����!�g̚5�MMM��`8�n� iP^wky� �����֖B�`��3?q~���&)A@7ǹڲ,zuq�\100�����.dp(Y]:�>S��̴�}g*�z�m�gk�+���8/��s}3�牀��@�M�z����"�H�V
��#z��b2�,�D	��c�Ezܛ!� (#�=?`&�����4����	 /�{!;��n^*��^5gΜ۶m�5�2kgk��/z��`2m�r��_�[�ы���i��� (��P(���VsMl#�b�Owvv�%Y�& ��Ў!�Yh	�B@��Д)S�l�%�4L�f6w��07�\�N���u��m�h0����|J ��z5�����P׮];����`0x�Y�X x���bm!O�s�1��?�O�a>�*I@O&��D"��Z]"�������x<�F�a�1�b˲�giP	Y��W"�qg�r��N�}�Շ� /y���yg!O�s�1�����d���!l�m_���*�G�Yuuu?�b� ������t���f<�r����3o���}�0* ����ϵ�Ҡ�	�F@����.]:��O�F
�.I�ӧi��*�u��������*�0��`2��k8?;�}S�TB��jՄ������lA#9��q˫���������ͥx1��k.�,�Pz"������5����%�e���2�
�k��z]�\!�I$��h�x}�Y'��>�˅B�{���.(�G�'XR����G!������q�S�Կ8�6tO�p~�0K;�ʺcʔ)3˩��x<�H��[�a� p���C�d����_�Z���������\�N�B�6^�[2�p}o����c�~C��@e��B'Ld�d2y�m�Ҫ� ntO!;/\��e�i���//^�hQc�|���Ϯ��L��1���ޯ�b�zx������v�V�, PY����>�N��ĵ�h��l�7��
��8�"�}FӋ��R�����tC@/�fm�|:�L�`ژ=:
�%�� T�?��������ڶ=O��	 W�QP@������h|��0�k��#�thu��i-��vGG�F��ؓu�+-a��ڤר�kԳ�~�D"�}m;L_ n�����t�;k���FA���s�ҥKkK�����^d��ٯ
�����>e&�`s�Ν^WW���_ ���,�η���R�S��P��O
���m�{����f&��*(������V�%R���x%��o@�9�f�:����_�444�����/zL�L ������o�)�1}m�b��L��( �]����.(
݇�h���,����&��n��+�y ��|����	F�F�mY�%�j &�=}}}�L$�+��̒m˖-�Hww�Y�m�j��������;���:��d&!a�@�,aHc��*d �.�Z�u�B�.ݴ�Z�U���Vk�u���jkբuw+ն
�X���Y0�%,If2yO��E	0�ܹs��������Lf�=�<�<��0@w'����	�ߋ��ζb�a,��?kǒ;찄ڕBDT�������|����B3�|>�i��)�x����E[��l\]]�������t@(��ܼڪ'D�~_"��������Ec�M!څ`0X����|\��
����Ocƌ9���!Q�׏��[kkkO@;�y�����L�"��T�F\p\n��iG�\*�L/�g��DSSS��g��M���_��~��҉v���8Et}s.�FD��u����u�H���ժU�6�7�X4�5�v?!"c�ގ�s�� 0@w������� =�����t{��������ի��hp�����o���jDT�����C���[�P6~
�G19^��h�f���Ս��P�~c��R������;�V='.�G�ɤ��:J�G��]˱�'Zq��G�*DD�����Bp���h,��ت��
mS$y5�o۶혒��AB�� ݽ%	M?y��'lnn�@��g^$����sЦX.D����C�=��K�Q��I�R����eb(�����8����?�I��c�; ������4w���ߋ{tM�)�5�l���7�fc)DD��RII�L�k�p�����N�x<:��P!�By!���Օ��q�p�c��b��>=q��AV�Z�"i�aX������D�h7��ͯ���<BDTwTVV^���x�%��'�}?�ٮ���l�m۶�p����V���~��Z�������Y���r��T*�-]F�v���j(�w��4!"*�Nl߈F�w��b�����Ѷ�+l���m�w_���h��"4`,�\.��ni�^^^~WW�Oq8D��Q�|	���	��|�@YY��8�"�a;��bq�H$����2�໅�HDvz:���q}zq�� 4`��d\P����ˆ����iR<����pݺu�B��@���3�c���0�O&����eRb�ؽ([���/��l��l����h���c��C0=�X��was|������W#��cB���	*�[q�""�%Qw� ��Tl�~F��_�������QޥR��t�7���"�I/�Ybq�����@ ��'��\6�oyG�� �K)����B���5�߅�T��3��S�T,�9�:	յBD���[,�ǟ(d	�NC��+������q�M�.D`~�e��Q���p�PA18'�қ�^��������E���P��o��Q^���z��`08���%�����0�a��l���ݝH$��Cq��=�Y---MB�\;���!""�����\���^q�X,v���(/"�\.˫�B�a�N�pj���zSSS[ еKO�%�݀
��b�G��A���""��N:O��ի�Ņ�����u}t-"�֖��ҿe�@�C\���,� �z�⚉�b�I+�7�&���ҽ�K�(K����s��dpDd��خ�F���щ\J�v��/�&Dd�g���;�y`:�'d�1������V>i<n\̼p�b�����24r�
Q��pY[[��p�+DD�[���8yS�J�_�����yBDVx<���;���	�:����hz��������.��Y�i����(cƌV^^��Z��l��~bw��{��'�_���P��y!������l�^��˫Y�:���g���E	�������sR�������5B��`0X��\�($DD��F��{��F��v�s:����:�"ꯆl��Ώ�n����ӎ�Y�v��Zګ�ǣ�@@��/��ci���b��a.� ���-�C!"��+�.Bc��=� =���ڪ��sMf���%��6��� ����bq��~��q2@_���h4��� ��\l#���kPo~'���ʹ�,����Y���c��r��xd�P(T���$!�1@�:���f�����V>)O���ֈ��a�늊�+V�\�)D9:�m²���х��\^�nݺv�~����)�=��BDيF"��l�L&�îR�rlt���R����a����������_/����c����Q�+���-DD6@}uOYY����WX4����N�x<O��#����М�v�(��i'�4wKt��z�L&���a���3���_@C�U�r��܋��v~E��l��w�sk���uuu'vtt<��	�ɼl4a��!$y� �v� ���`�6����y5X�q���4��JNG���\9��?��B����2M�+�/�Go
���ʕ+7�B�c������w�ѮD����l��P;���ps%�ԗTbga��O\Rr;�;_���g 8U�r�k�WTT<�ã�h(�d�ȑ�J�d˖-���!Dyp�.��%@���ܼA��*�'}��NP��˶s;G(o�Ӯ����V�BG��g�~�J։��M$���n�i�Vyy��8�'	�TTTh�f�VYY)C�e�N�P�bv����A��ҟƏS��ާ��;���`0�7�>&�7�iWj�������'Հ�{b�Sn�v��B�h��O��X}ӈ�Đ!C��siiio�>|�pٺu�l۶��w��畔���!Z��AzMMͱ�^��e�׬Y�(��x��P^1@���%�,���?������|���<grR�/4�>���s8'D}(//����=�Æ��5H׭��[�������By��������ե=�8�h�ٺ�Ҟ4q��A�}N(���.�B�� ���D뭷��98<��oۯǎ{yCCCB�����z�����vk���{|�����:����'�'�,�z�Z�j#��cp�>�"�7�mذᤒ��}��:���T*u&����s�V����k�/�~���"8���hp����gK'����=�^u��S�N��������~� �X�D�$��+�����P�1@�=9O��� X$�1`---=�k��@ 8?��L�������^��u���4Pg�:eipOO����&�W�WUUUVV�8~<B�\m�?e�8���x<G�tړt��H$���'F��;4B���C��n��b?�f|Ѯ�r���E'�[�vC�ֳIoφ�����g�u�U��A]�i��m�����՝�ks~<L�ܥ3�J=���^��(��By� �����[�����F�����.�8����[ZZ�!D��\�I�F
�h����[I{�u��n�d�7X����=&��z��7)�/ʻ�+Wn��},��G�}J��c~,{gO�uQ����(d蔍3F�}ٺu�ڭ|RT������+���(�R�/!8�c�A�;�T���$+�(D���I�O$�����Y����e�.�E<�
�NL&���qB�hݙ��|>���Uق:ecXEE�.���E�4F��z/��)3�)��h�)�4`�1�:���9eeРA���v)++��4XGpЉ@�%ݳ��-�Vg�Q|��B�hnn��ç����Ə�	Qq����d�@�ǣ��B�`�N����!@_�fMK О������qb���B4@8�>��\�R�K��d������8W H��W_��V����D���|��X쫄ܤ��S����mt�V\o�����/Q�����,�n\��H!�0@�l�k�p�g]rM�G4��KːP��a�c�9!eM'��	�lЂ ��T*� ��4(��t�i��7�������}(�q�x(�������t�rR���cO:���d2���e��N�N�B�� ������Y�#���Y�h���Dz)]Jm�� ����Kш�Q4�]�t�k�>AKKKv�ݣ?����\>��<=�;�AB��`081�����,���\]]�;۶m��Tl������'j��E![1@�\�
�.�z�tz�s��-��F�r���[��o������~hٲe+�|���������ehp}��$�����9�ǯb�M!��<8��~�k�{[�l�"�L�R���7n���![1@�\J&��P�����jLii�Nx2A�rd��p:���h��Gy�����׊M�i�7]!Co:x�~-�Ͼ��?�X�̦7��0�9(۾�MoY�����aÆ}O����[��QA�x8�G�|8o +f��������/ITH�PhdYY�S8�_��aȐ!��շ ?�KC&�'�H�W�X���G{�������*�JUc?�3{]NG{Mt��ªD�v��a�V�3�|����C��7n"��9��|��8�
َ:�j�ڵkO��A!2*�!�Dt)�IB��s�=�9б�p��:t��.\��I�h�3x�Q(�@����`�i�>�G�
�)))�3��z�@R��h��%�ȡ��D"�<���<��:�5�,�:A'0A���Q?e�{��sQ�_
��64v��������D��A�`p
�K�l� ��n��-//����K6lؠ�!!r�?��q�@���)B� �r��~���X,���E/*��px��.�V�^����&��y���j\�y\��fu�5�����V}}�B�9G��eee�A�������<����l�s�B�9eB� ����K��.P��(������)D�3�����ǵ!>W�CCÜN���fM�%[}�����h`�*]-�����2jԨ� ���[�L�r��ltH�W�
�:�.���|����� ���;O��z�ip8�����+Vt	��s���op*�:�_	ٮ���d2�KS����]�A���'�;���(�=��c�¶�P�0@��*�x<:�J!�Y ����h�h�|��>�Ùpr� � p�~��y��oѢE�����{_֖f�h���M����C�u}6Jg'^$TP�i �V[[{�U��J�Ap�wv)D@�s+�����l�M������|8_*��� ]�p������-[�Ye�(cI,{2��|�9}>&TP�i Ftvv~������I����6��-����zk�����A����1@/����'***��ᨾ���a�z����v.�F�����nD_!Tp�i@JJJ.�ÿI��K�7�@`�l�`�EV�g�ڵ��r� ��>
�&L����&d+��m]���]=&3�$�J'C<�����u)G�f�4P~4pO��~!���n>���&�FII��B9C��a�B�H$���O�
Ao����Z�޹��krx,{�� ��e� ��d����p�=�`j�Y�H$�B�?��Nw�F��e��K��P__áw��e���{�ޞ��..A�C��X,{9������"��:Y�����@!�P�,4z�����!:^�,�s�6�~�t��^p5�w��>����:8�S�p�^���j��ȑ#{'���qd3_�����+d�d	TBWc� �,3q��A���$!���#F<,�/�كn�,�z�����rɂ���L�K���X,�j6���SVVv��1��%PQ�������h�t�@ �{)DֻG'{�YMM�^�q�������Y�fM����,Y�,��Ïf�;:y���oذ���)�t��{�t	�񃅌� �,��x���	B4@~��fT��Ky�����~�g��vsxA�:ͺ!N��4��s��������4HO&�B�'wD�ѕ�<0=��kBFa�NV:�������e��S0�@��G�O_�fͿ�����f9o�ĉ70#�~�gv*��!s�c���:y����u�V!�X{YYY�7����/�n/!�0@'K���\��,!�@ p*v��<Au�P�!(��f�iӦ�
WR��+�������������{{�u\:�)�
Υ755�e�ت���8/2t�
�����\��r���݃�#D��e�<�~����w�=`�C�D�W��***zǥ�RlLy'�Q�2�#8ײ�s��:Y͓^���)k�Ph|ww�.�6T���x<Μҁa�n�C����H$�D�V�T����3@{Zt��=�B�_h7�:.�{�-!#1@�|�| �>�	*�����F$������<Bc�.�~�5�����B&���l��ظnʔ)�!0:v ϣ/VVV�l�\����5��f�`�Zf�2t�/���}E�v#�m۶m'��j@�e�P����T�B�8O�0aَ=%Ki�����Rl�����-D�B;��(�Z�/�{~����S�|���݌��h֮]�+T*��<��p������*O&��b������B�s-��Y�M{�;;;�(OD"�g�}�A���:���c�N���x<�`�����_���ko��<��h�N�5�ͅ����p�憆���m�/_�eʔ)��Ϊ�D�IF�)۶m�]�����nt�R�K�}p(������0�S>}����'---����DC?�u:��ڼ�+Wr`� q�5�U������\!�i��ez���k�:gy���E.٪���:��Z�h�)�<�T�:�O�4�m������&(��$4`\b�|([u�$�6õ�$v�`�������y�fٺ��P���󮭼���l?f̘ax�B�c�N�v*�����ǇP�,��!�GK<A�
�
��0��P,{U�6:����^'<=?ϯCK��ۛ�cә�BiW�Z�jc�Fp�m���� ����?^����(촗�����lg��]K��˴H�x<����l�rfv�􌊊�ޥ�6l� ��p��sYV���탲�!G`�Nv8�����^r�Y�fy���+--�;�L��}z�`κC���|v�!�(���F�q!�,[�������q8>����iʻNǔw�J�n�fO�^��j<|��#0@'[� �vG
�����wvv����N޴i�NpC�B$Y%4`(�k�V�e��t���	�F�%�sp��2�WS����{'�K��$�2w�nk���>�/���B�� ����`0x
����R8��Ϡ���>��ڠ׉mt�"����p֙ �8��^UU�����-B�I���6	�����>�~���D"r�M��������P�
!�`�N�A�u3*�g9�xL�6-���}���n?���ʔ��ٲ��C*�-۶m���%pm3@w�Qhğ���B�ill\�W�p�]��ȍ5j�������ϱ*f�onnn����@�N8'��0@';����ƞ�Z6u�ԏ��>3�S^�����	l4���p~�Y�n]��U�;��K���7����~|�7����ǎ����>����>�<]�����w���1�`�ItN���I?��/���VZ����q�l�:�[SS�!8����|{�4zg�%*��[����������	!� �sz��'U���ի�ⵏ��~~��+T4���.�����4��v3�v�����hg��n>��s�7	��ZZZ�I�Dz"�����NV�~�zNZC����^�� ��ߝ.�� �F���-���/㳷��3ӦMۻ���_�G=�'���B��\�q¹pkI_)���9������S!\��ޝh@�#d�ɓ'�FA�iM_/++;�4�?ϣi�ڃNT(ڃ��)�-S]]�Ǯ\�qp���@Է˅�4[�O3�@�T��? �{q���TTT܊u|�����6��.��p��Bl~�JsЩoЩFz<M���PAM�:uB*�:�3�LGcn@������%D����!ˠl`z��]���B��90�mev�.^���Uz����CxOwIC��H7�^��9�O�8qP�Aȉ��Ӯ1@��@E��@ ��h4���m4Uu��ɓ��>����O�Y��[�n�݈
liKK��B�A�1�		ΥA�k"��![466������36���|�ѢE��QS�5������9!'iI�R7���6m�&vC����N���egЩP2w�XQ�ٌ3*�l�r�������d!�.��\�;'*4Mo�ʎ	c�=+�u���W
�&�&���'�L������a��#P���m8�[�x��.�ebe|�{�w�+�*--ej{�S���n�F������G!h>��	(�O�?��k��:c;R8��YJ{Ѕ��k�P�����\^�&�)++�;�v�K�i���"P�;a�F�#=	,��H$�h.����Z�F���������dz@�~��U���Y�h���5�,���cʏ�V��^/=�tR��d���h\�jНo��+��f���[���|�a�KO�:u�G_y�]�ijjj��$���	��<�ħ~�ZZZza.����>��x�C��S�i����Q��m۶�AD�r.���L+�T*u<O�I���YZ�|Ҟs.�A�`z{��
9��o�B�_677w�"��nw���R4��{{z\,��������G�8C�8o��kuu.��v�fN�:1a�4����ȷf$�.����$�H�)�n�����ڞ͚5����t5(��T�
�^8c;f[yyyN���g�G�^QQ���㡮�L&���B��g��V����k���e���5kZ��#�ӥ�~�m�P��k̘1������.�{�H�����,̝1@w�����S�J���p���K�v2}������Gy<�����[���Y�eb����xtժU�,U^^�����mԷ��bL��544$���\^`�KO�4i��ؿ�̓Ӂ�����z����BI��8_ϝlA�U���Z���w7䒓���K��bX�ua �+��KH�M��w*�:���4
�a��a�^�M�6	�I4�T�r� ������u�Ї��e����;kj}Vzƚ5k��k~:Α����q�m��.�=����mذ�r|o����Im�a�N��Tf��R��\�9��ĥ�����OԠ�'���S3/tR8"�l�k����������m�.]������8o�K�>cƌK.\��D1h���o
O`���l�Ͼ����D��f��hO��k� d�E�	�Ju?2���N����@���)��35�G��Π���GV�Xa���b��6T���b3���h������p8��l�1b�ћ6m�N����˚�
�A;�Z�x96�P^y<�o�������tb8���ˊNL������^<[�lS��UUU�s����)�0��L�>ɛ_@ӏ4��3���� �+��lك^��Ǎ�MR�Խ��Е��ޯ ]�g�����f����CBy�vֳ�h��\~�ˡ(�g��4K����S�w� ��t=B�R݃eee����CQ��CP��Ù(HOľRf������)D�PYY��P��*F��i�]cc�h�;��u��8���@�d�󴴴���8���7=:�N�(�_�w�������͖����-������]�^���b�qYMM�}�^��<y�h���iM_Ǐ��g�}Ie���ٺu�������r���P�қ�'�E'���ͯ9���T��=8�'�F�:��U(A�p�?"d	|�?������w�=|��0�w���1@w���R��.����������:��AW�ԩS'�R)m���x<���K0�HpR82���'
�A0X�XÑH�A��߀�c��j����X,�(���v�p�w+�m�[r�\���]'�۳Mm�]c��2}��+��4H7%����@ ��-��{�L�<y��������hF�N
Gd0���Q2�
5�]W���P(�"l�����|]�U>�K�.^����3�F����$���8�&���C]�r�ʜ��Mm7n�d&���c��2�
Е���$`������������3f̨زeˡ�S^__����z�05G�&��N�CY�(���� ��w��-�F��	�A{�mСu�i��n��y�foz���������S�;Y�%լ� �e�4CfVwC�ν=ύ���o��kРAG�39��I��R�8c;9�Lo�#�9yO�өt���	��s���~)����ny��2���`�q����l��s�\~a�����J���NG�`��2��AW���:1�!�������/����'O��gq�P��*sKCUo�����Ƒ#G>+�7hlzz8yO��w|����Hd�P^���K���gpx�������I�&�_�l��|���?h'M���������u�|V������w�H\�WS�u�9Y���dd�E���������+
MJ�Ǚ7S�N�h*��J���M\�"�t�=Љ�	�������<��u������m��eKKKu�����"����c������~�P_��D"��:�#v�a�3k��F����̞z�3�]�2y�D"��|��'�5k������~'[���+.�7dt�9Jr�c���{������u�'���G�یm�ͯ�i�y�3���(�g���s��ϰ�؄���r�|���@@�(7=��Lm�t�^lz�m۶ML���*N�:�����wvv���xTV:�|��{��18'�H�LxJ(�j��kJӒOʫ����S�Ly����u'.Y�Ė�����玚����މ�B��\�ǣ��ڿ��8S~ii)S��:�^x���%�������$Y��EP9�N)�4!�����un���DYx���e�P�L�8Q'�#��g�����b�W���~)̐�3�}��DY݄s�H�[��ǟ�͙�y����>�}���PcEj{��;c��2�^z�mݺՔT�����.���==Ay������\ߥ͛7KggNKp�k���ٻ�;���2o�]tFw�����Ѯ3lذg������,>��g�;����(�zw�?�Y�ʹ7���>hK)�Y�|W���`1�f�Z5y�>���c�B����ݔTw����z��5k�����������)��+�A����sR8r\׏���r�����h���Y�parʔ)��^�{ү�p8����S
`����(����|gc�c����.�9�_$N��i�V��38�tڣ��D"���|)�z����#3g���'y���T1p�	�����9��V
���qB��Ʋ��&�W���m��;=Y\A���k4vτ	�F;D3"ϖ�|�ر?��Ə��Gb�Lǝ��� ���SV�b�1ʆ����~����|?W
�L�Gw�����6� ��;�?4�D�ʛ%K��\__ߌÐ�/=+_��|>VCNS�����✻M�wՈ����J.���5	:Vݸ��:����T�5;c�NY�L���M�e˖i�~�^�V�pN
GN�J��� ��8r/4�o���L[�y���)S���j�_z|����	1@,{���nbGG����؊m�[[ZZ����/�yq�F�i5��j,fv� �����A������o��b���#Gr�y��s3�;$��k֬Y,d�Aw�z�߯C��"�7�T�>�a��3i�F�j�ʕ:��b�������I�>"�A�c�4{uuu��?�d�_�������ЋS�]3!�]�L��nȐ!B���ˠ	��r�eS?l�S�����+t*t1[�t��/��6���'N�bŊ�b�x<�>]��R�x��D���$�b�X֍�tj�����b�|��g08�t����<x�13�������#��pR8r:�_�{��í���r�s��IOgw�>m�d�z�FI��)>��E{���zG4ͩ��Y�MLm�v6��ڋQ��Xq�*��b���t�5Jh�4�a���I�5O������]�����|�����"�H������b���t��qzF$Y��o:�����،�Uލ�m۶};�_�������v���N���:���M�Tw&Ӟ�͛7˰a�MvYh��,B���o�}**�z!r�5�#�w(3J�(v��Ĵk#q>�گ�ū������;>�#l~�c<��1˗/_+�JORxG0\�����d1_���׭[מ�/���?�p�FS��~Щ�2��&�������0�r:���N��xtѢEm�:�����-B��މD��fR�~µ�U�#�E��	��llv�h'|���p�Hdv� �����78#��}�K���N'��h�Z�f�~�]��`ZǳkO�	��Y�5�݅������	���;::��q�Tf����"�K�Rn�d29Z��?|�lG
�E"����ԯ��I�4��� =#����|4�?�-�TTT�ڎ�g:��+�0����0������^�����AS݇w�0�~k�6����C��m�;}�@`�NR"D�a��-zzz����d0<1�<&d��^{m}}}�Ө�O���?>iҤ�˖-[-����q������'f����K�e���jhYY�ݲ�&�14V�+���3�������BЋؤTw�iP�Z��Bsn*���v��	&��n�8{�����@���0�� ������F R����i�v�%^��t썛�lO����PhR2��
?�V��ΝxOO���5k�Ncgj;뚾1@���i3e}mMu�{ｋa�L�$o�斖��eѢEY(��Fġ_���?���t�Kmgg���� d�#F<��޾��6����;.@W����]�,�{�?Y��G;�\~!�w_�hj���9���O����n&���b7n��#G:���Vl�kO9>�ǖ-[�!�'@p�c��l�(�������F�������Z�fͿ�,�p�p8�(ϱ��?���XCC�c'�F�+�n:��󝍽���^������kh���>��ؙڞ���o��2&��wuu���:T`>3M���iӦg�>���"!*.�m�1��^��64�g���em5|������+�,�;�`���	&<�H$n�&��+�>����z��#��D�#m�۝}Z��>1@'��E�K�i`l�Y���]z�	�ls�.]���@������ЖX,��:{1@��9�����%d����皚��p8���<�ߵ�-Rh������ߤi������ ��u��k��!��d�ڍ���� �e�}!d�e��BӿUS�u<�w��[��� �J=���Ҁ#��s?��!BT\��Z.��w1�g��sK(z����U�2s�����s��L���ɓ?��ߥH�b���'!��?~K��y�A}nKK��lm�#�V�ZS���_�v� �,���Eױ���K��q��vϹҫ��?�A�����5�x�t��N�2A�����W��e�D"�k��.d�t���C���^4�����y������>��sIm7n����R��ߨ%Ք�
�ك�7�d�̝8SR�;::zoh���Ea���y�����˗o��"8��W���� �~ÄhP�����A�|!�466.���_��Z�_z�ĉ/^�bE�S -�@�5��G{����G2��h[^����%�VtR�j1�-Dj;����R�U{{{o������O�R����O�Y���9��u%A�4===K��6B����x��Xkk�Z!K�dg�pX{Z�g�K�]^^~�l������&
�K&�7K�'����Һu�ڳ��@ p)^��5��H;�t�s2t���MIu�Mu5j�Ui<o`�^�K�.�g!f�Ep�/����x�X�!���)++Ӊ�N�R!�L�{Q��y�A��4�~��y�\~��TK/d�x��T�nif)ǀ��:�I��z�` �ѻ�-�6���>�x���I�3fXyy��.*n�	S�)����h��B�hhh�O8n��d�_���'[�b�f)r8_��������K��ز�%�?h���5t_��6H�Y���Zh��7�.c��`Z���G�4�!C���|���3���ytѢEmb������>"D��_B�����|G��d���|�����U��� }Hyy����'.��А��`08m������<\W��m�<����0��9S��� �e
�ʢ��Φ��	2����A�A!�>���4�.2*���g	Q�c�n�m۶c�#�C%����v�Y"�Jݏ��&��oMswE���DtR�c}>�	���c���+�>'��:1t�B-�F�c��2��7u�˖-[�IeɌG׻���c8�?t�п-\���5�Q�O����� ��6+++�Á���H��!��0]�5���v���d9���ǚ�5h]�����Ů���G=�37G�UVVf=���q&�w���̄�v�=�.S� 93S����@{�7lذ�˖-s�,ѡP�
��\�e*z"��<�![�R������M>��Y:�������Ci"�8�ߊ�Z�j#v�<�m��p|�/d�B����Ch�ރC�&3��� �e
���c��gƔ�T@uo����84>@��V���爁kh���+Wn�t�h � �]WW7�o�Ѐtww���	v�4wW��x|���jii�*�+
U�;ӎ�Qbm������1}bE�2���p0)����wE,�+�{��Ä�%��^�������ɝ��:�R�Y�lنp8�$O��u�2mڴ��ŋ���p.��IK�}|2�ԛ)�b �b5�l�'}c�N�2-�]z�R�]555�����NO��b!r\�F^��8��C`s	ꮿE"�ǄJ��mС��b���&
_��+b Mm�,V���O��vZH��D"!��J�	�BS���7�A|>߇�`�]�\���l�t�H	�wjz0��5B�6|������:.����E|�0@�Jz�_��LMm��c�N���:ݠ;gux?� �L:���F�=���8!D.���� � ��d���2��lԫG�R�:�;�ᰶ�h�K�?y������ �M�~��}M�s�tuV�TzGO�^ۺu������׈���i_!r!�+�l�@��c�BG�^�R�; �&g���b^W'�c���@`0��y8#*--��L���>���QQˌ�1(�]+���~�k�XlN���Â`0x
/}/�E'7���ںV�vڃ�Y	��u�_����ꗆ�������P[Wr�ww&��LH	��N`���]8�"�^s�V5o���˘����Cǣ�RƔ������D���
�f"���x/��p����P.��YL�5�3�ɨW�ʙ��pXW��{�Xߔ)St�����؝!�2u�����>1@w�^��+Ku��	&Lkjjj+��A��_�`�b:���wY���匧�:Y�۟pn���y����m_���i��w�6�1�� ���T�S�i���������P���3��hnn.��p:�1c>QQQ��	BT�8��@<'�|9���]����r�dɒW��޼�un�9f���}s�ʕ�B:)�~('ġW�YΘ��:A{�KuW�=݃��s&��_�v�f��S�~����EBT���Z�����a'�ί!�Y�ǟ�>��q}����k�ȑ�c��5������~�.y����YP�� ��a`�{�cȯ��:1@z��o�=5� �U��K4@o
D7x�$���/N���K�R���;@W���� =
U��ϠN5hРެTr>�.crψ*����i\�����h��b�X,�����f�ީ���,TΓB�GrƦ�G?
{�o9X�t�S�Li����u�z'���ʆ����B�����t1�Sfm��fl���˘���cѓ�do��A�C�S{��,��F�O�|��t+��v\g�S��&G�N����j66[t��㓰�G\m-=W�Ce&\��� �eLox�8��a�UK�������Y��E��Ǐ?����Q1t-N��*�������#��#BYC���n����gsw]��s�h�~W����� ����C-lLKu״<��'u]r��r]�z�[�P��d2��W���%����B�w�Q	��?  ���UBYihhxkʔ)�gw��/}��<vѢE_~�.87���b�L���t2�6��k�?v����&,������l���/�x#6v��#�1�Z�`P��zz��N���ۂ���i+W��$�-Ms�;@��]6�_���S��cvk֩��NŇ��8�᥅Ζ-[L|χ��_;�͘u��K�ݔ���n"���k�7J�R�.�C�گ���O8�N����ݡ,x��y��C��3Ms/� =
U!8�{��tR8I*N�]�I/}�Z������k>��m~]���⽽�B[ǥ��A؃^Xh�'���NF����(�G�-�T__��I�����4iRݲe�VJ�=z����kp>AVZZ�;����\�����.-|4�=�H�iP1^WE"���a���2����}k�n�l�D���xV�s�&� �@�z���-�-ʆ�����M�ӱ�^�P8.�������d1��T�K	3��� ������G7����-hP�E��^1L$YSUU����2}o��tww�*�mBT4�g�WK���nmڴ�����8i�Kk�{���y ��v���jGŒ������0@'�e�^۶��v���w�|�����sb����-x����
��d���D���5��D{4���{�އkkk��Z�j��.�\������!\�_�����Ó���w+ʿs�pŒڞ� �o���@�M{�4�������3\�*�IOdwu0\�K�'�#sŅ

elG15�ȑ>��Օ�4�"�>��Е��M������/�e:��	o����8�NUfVwC'0�B���wx<��(�<�����=��:^�̳F����ڶ���;	��5��Ph��-[����^ol�l~�3f͚u�9s�Z������M� �[@���>1@'G��i�֭b����)4*��ok��盂~~�!Dfa�^`�c�p8H�
�Z���G�ѿ�I��p8� ����njj:���`8����O،Э�M�IJ��o����ʠA����KU����	&�ʫM����{<����?^$D�@c��tmK�Th�U�ǚ�������.ԧT*u���)Dz���;6@��|���á�cz2��{0@'����2w�޺D"�t(�Dss�1!���@ ��߈*(*~h,�%d�GQ�G]�Pmm�TN׷��Ɔp8�?b�K�VWW���N�����F�:*�C<K8V�U��#��L&���|�O��qc�h4��������y(��
Qa��F.�A��o"��u�ɜ4�o�\�����YYY�i�	��Y�;v/O�/�5�٣�.�]�X&cp@������@8�lCCCB��������l�S܍� ������S?���v���>�����ͪi�	����\z�{��Z�Lmw'�ʤo�L�E�A��w��Rd4@�����L������?�s���}�:�](:�����YBT �F��n �W[{8�.��{�W���+�>����N���O��V���~���h#�����qI�����tCl޼9���۶m��jZ�"C��3/�!Sx��k�;3$u�R��󚛛;���~�Q0�)���A7 ʩv!2����jjj^oiiyC�f��zʋS��[6nܸ�^��iֈC�%���c��� ��pb�wp3�oZ�|�����.�F��)5��.�L�Og��s����.|���|�$��n
��ơ��"{��]�v��	�=��tҸUUU����zO"������V��m�v����-�B�k���Rs��8Df�����/����<��SV?��}���۲�^{���gㅠ��09�=�<T���ÿ�H$�K�{��g'
Q�Ņ��=�%�� s�p�����('� �/˗/_�u�3�۔{p��ɓ��ˀ
�B#Q�=���Aܐ�N�� �@J��~�<��_���N\�O2��ս���"��Y�/��b���3�|�w�s�%D�e\�έP=����s������q�E��������� �3���D��d2��A��������1@/�Se��y�	�ǎ+��#�Iu����f0�D"����)ǟ:�
�K�|b�n��==L;$���1�M��F�7	�*++{A��p8�����1zmmm%>s>E�M���k�� � ҽ����z����6��g��1XG�����f:|�����X,v�8������� ~�"�1@7D*��\R�wr�Q7�7�8f��|Z�hѦp8� �3m~�ӦM�w������༫�K{��0o�ܘ�κ�o�c��<Y��g�b����	w�P(]� �uĺ�h �����b�,D�k��t!r��u#H?u�!�����k���]'���|����Lm�az���a�dp��9�]�߂��^�=�;�,����9���F�~�8 �g������<@��tC�t6��A�|}���O�����'��f�(;_��YR� m�h��p��KKK{7�g�%%�Iߓ��@�������?�1m����}>��6���~kx��BN��D"!�m4,��x����ӳ�^��B'���'���� �\�����<ZUUuxkk�q�+Vt���px��/��ɓ'�l~�L������L�ю��o��U)��uS����v��S�fЗ"�����8vě�F�����x��	��0@7{�ɉp�N.++���YN�G�H����3k������셶���āt���æpJ�^T-�=��B�A��ڸ8_{�QP���E,{�y
����1B�Oh`q�!P�l"g�����-]����zM�����h�>k֬oϙ3�ێכ0a�X�:��Q�gh��2[)wN	�m����cѕSݕ���=���{2:z������4޷�����f9����F�s7�ȡ�Y_�r(�����i�����������bƽ�曟����~���Ǐ���~��2V;�܎�Z}sJ���D�pS�K?'�����ƅ��Y����;S0�7��q�e�P#�������(b���R��g�Z�})�t�{^�����׫�Q+�C1Y�Ү0@w!���+�;u�
]z�I��jkk+����|zR6G�D"���<����!��:!ctuu��E�p:Q�`0x0�U�BK�,Y�_�{���:m����x饗����>�6�sbs����Y�i��rv0@����It]I-u�9�9����I�'#H�$�f͚TЇ����GM{w�� �����nݺ�@ ��;IN��;����N_�j�Fq'Ms�����H$>��_�~⚚���M�i���P�6)��8%@�t��0�FCMu��af H��gt��8Dz��U�`�%�Ql^���et��Dq����>���5ẻ��� (��S�����x�3�� =�N:[����-aj�{z8�ON	�كn!7^��8�n�*����}>�1�x<*�)�x�i�;λ�QИc�n��� ���g�~�mRD��f�W^i
�Ë������:nҤI#�-[fɊ��>��|����:::zۤLq�N?��;q��ẻ����;w{���N��~�������ѱX�� zS��x�����	gy��9&;�E�Q�8/�7��T�G�D�5@�
��b���>Q 8U'��a�Ly�K ��H҅��.8��(��z]���|1hjQ2�tb���� �����w�8H:��Z���o��X!Jc�����"�z�{oE����"�T���~&���u6���`�B�~%Exc_�t����렳�oN	���mn�X��x\��N��ٮ����y؝/6�d��fuwh�0�tOA���8��g����w������=�Tlz�_C��u�K�����L���<����x�t���W_���������D����+7�=��� ��g��@��ʒ�gk��i4�t�ˌG��4��c��ΊF���� ����Δwb���S1�����t� �)nk�����y.�������w�9��3@�3��P�ϐ;Ү�^c��� �Tw�J��yүB�~�8Lz6�kQ	��)�8'�Z�̓kt}	g��7��'���imm]+.P^^�A�%w��/�i�Y�uuu�h�܋�g�����t����z�D��	yo�����6l���i/z*���J[�7!��ǯ�y�?$�=�F�A���ŏG�Rgg't�x<��l4Q��zg��盁�ӑ˻����G��)S���������u?�dɒ����u����..�� ��L���/d��ŏ���*++�7���v��A�N��d%%%�!H�S���h��ϤS�u�wN��.=mmm���<Lq�b7m��Q�������i��i�&���{����C�=�m?q17��A���ɸ'�8|ۘ|��СC�{��I�˙��������IyOb�)�r���Y��,Щ�i*���o��R��j��KZ�m��)�	�Q�O��1�c[�I4H�6��:�=��� ��pR6!8Ԃ�lZ��#F��ݨo�ھu��b*�x</���t4}S�{��ѣ'WTT�*.� �8�����@nq�MT?��HkhhHL�2�/h��]�~h������Ɔ�|�����v��7Zggg��-A:�z���\� }jyy���d�b+���u50煽kE�ghϳ.�v|<oZ�n�.�x>*�g��]l��O�c�n �$N����`0�D�"����蚭�i����y_��Nr˕\��A��Qu(&�t��BA�w5/����4P�v�2M��Tm]JM/�=�w���t�"�3��Z�pώF��C��%
�3�L�?~Z�(�:d�n ��N.��9?���=�H�Z�dɋ����q8��>}֬YW̙3�;���������x@�av��t��E���͍.�����M�����&��X�������h4]��LW=�*6L�6P2�\_V�%��4������C֬Y�"E�h�9�W��������=zt�%���ㄲR���==�+�]ȭ����*�Q����8ûJϮ������R��q<U�h��\'d����-�@����*$ڵq^��q�7�����0�(@�.�D����ߊן,����tr���%d���0a�)MMMm�Ph,�����>����� �Ě�8��P�4��B�.M�R��B�����;��466.��+p8Ѯ��T�7��2Ž)����b��Щ��s��;8$�H4��a[&�^���555��{ӧ9'#3�s�n���:�A\���-*�����#;^K�_�6m�}Y�a���]�M��&�˅3��  /�IDAT_'��gF"����ZZZ^Gc����Y`���;��B���r-�1'���9�)E��h]/y��ݵe˖ލ��A�~��b/�.�I�4�]�sz�a(�
ߍ�b7�8��E�7�&�-Ob��7ݑ�=n2ꊷ{xs���"�1�h4z��W^y�)/����x~-76l��^�/Y+�H���ޓ��e����.�̘sꓮ����7�����+WnC��5TT���s��-�F9	{i��b�я��`[$�[��Φny��������)�!ݽ���v�����	�r��{� P?9��G,=���Ǐ��J�~��g
9�/��
e�Z��DR����o!HZ�D"�x����ba,���oܸ��/�8=ݝ�ɮ1@7���`���ly<�z�Y��|A08�هq�,F��4<�[�z�[����|'�����BF4hǠ
�к�p�2�+�n�D<o�"�|������5~�ϧc�7o�,d/MwW�^T� ������s4(�\h����<X�&nlTq�y��@���@ ps,�:��hh@ͯ��{���C'�����3V2�d���F=���x<O���x4])E �N7� ]ۮ�k��慣��vLi@Ł��C��~��ٹ�@�KG���ȑ#]u����1��wt�������=kժU���c�/��|�C#�g8���i:���k(���d4�'�������:~���;���_ݯjp��慗ikO�S:�X����t#v߱�y��|�w���R�.Ŏ�������|���洖��7�����bw�����2*g��,�J�-)a�;�Ԗ��=�:�H�/�N�[�hѦp8�+�����j�����A�A�=���� ����.1@/��I���]M�>dȐ��{1�έ�ss4���E�h�.)hH=��Ȥ��6My��H��¹� �`Lq'ڥ�=��)�444�l�t6��t�on6m�d}N��Û;�� � ��	aw���K]���y��#�D�>��������)��/Ǎ7���L��M���G�p�P�b6v�صmmmڂb7�Ύ���G���[�>���]���q�Ro��d�$�?�Iw>腡W����$�^L���4ʻ�&�ɩ�gF��7�H���[�3�����#P��ߔ�7%�^\�`zC׾�D)�
��:g��~-�.�Z�paG}}��%%%g��q�+�iӦ�V���tb1Hw&�6C���9����|� ��)%�kEA�9[#!��b�9RDғ�\���7�6���
{�m�Ϝ=���k�:Ѯ}#D�fq��l�}�Liw.��� �~G`"6һ�:��.æ�<)CflMǭ�m8Λ�9����+V�z*1��3��Կ�m�P^�:f�n8���i_!���	��w�:o˰aÞmooכqcv�w�tX�3bJ�s���-�k���@���A�NI����cg�6��Jl�~��z)���p��1�F�**�kjj>����$E&��	�\U��O/:$dA�tUu��!�dXd�Ȱ��0#�D�����8e��������HDǀ04饖�N!		����y��{2E����u��.��y��[�tuݺ���=�w��I��9s�|����L���eD�P����x������ �|,�H"��3�-[��?��h~վ�`���D����l��F����>cĸ��~��k͹��X.�{!���N��1�������[�}��S��pǅ��pEн��Bb�0��$�*�L���<���y�7oVJ{���Hg$��Fu?��_�*R��ߜ-�sO��c��1�n�]�n��&����������K����f���F�Bmm�����r���	1f&��z����t��#���g���̦M����L(�m���uo���o�k�I�s�
�y�/444�MSS�i�Lf�	(�:L[|$����|���u�%����^�B�T<7��={�!��'`?}����(c&�H���tE�]�/�Ĺoh���}*�]�N�����	�d2������|c�֭���-��5�h�2�"H(�]�q1B�<?Gx��9s挺�:���г
�H���t�o��@��_i��@h+5�����h4z(�NU�@��ں	������T<W_��c�;�X��r���4����(�"D1���u���.Λ�������Өj�Hg���j��[
�GRt���ȹ�9��K��Z@n{�״D"ј�f�@�l�#FEt�w!���c�7���=��`�j�߹Mn+ZkD(�6��LwP�~芠�����@0�� ��?��R��&$��������u���b��2ڧü�����U��D"��*%Ĩ�0�=���R?�9��b��p�	��,�O�e�>�x?�\�^�zA�"�A���G455���d7!����9�����t#����l6+��q���߈F��eb;Я/��r��R)�Wl��Z�g�b4���dB��N;�4(i�3�S-�>�zA�"�A8�05�<����y,���k׮� �d2o��CZss�\8s'cP:�e�	9���Jq�8,���Y0�!��Ox6.�0_f|��Y���8�͏��P[[;(�1�l{m	�G����}�+�&]�0~芠�;*�"q
N���7p�τC�	)���������x�`�u��6ل�3f�n�Ƨ�5�B����N�����XSa~V]]'��[����Gͷ�"�_����pMz%E�R���>�:�m�����o��>���0蜍�8N��I�����_��޾Մg_�gh��|��q���	M��+V���f��k�/I��w�l%�����N46!������}Q�x'�?�SI�>�zA��^�l�׳�r}�"��}OVW�=g-^y $�C	g�.�f�'�q8Ύ/��I*�z��h�x|�ϓ(�q<�E��C�"���|7�eR�G�W4 �dB�hQ�H/L�#�b8��pT��� �Y�p����~�zO��x-�]�<��aq�X,�o[�n�lݺu��h+�d���h����:)�,.�h���s� �.��2���~�����hfB�Hk�ǊDza�Hg��Z��4���;��*�fS�L1^�Ѷ=�U�>����s�x�\��ǌ�Fgg��8�SMM��p��8����4A�	��z��(��#�Ar�෌Op*����FQ���g�&�t8V�O�4I��
#�^�q�#��FLO�3�^@�\� Ӻ�"�����s�����Y��+ȳp�r"����⛨�P]��^����5�G@�؉��7!�b��m���R�u��l6k���uQ�{�@������d4� �S��a�5}�����T����b!?^��⬽>������CF����ZZZb�<����$��T���O�}'�.�
���1�^����n|D,��Õ7�n�껄��SP�-��ͽ�%҇�t��#�^%�����f�8��n�~v^���X5f�$�cbE:��#�7��x<�kp~WWW�#���ʈ��D"� ����WN�5\`��m��O�s�-�L�Aa���d2Y�½n�1�k�o��eB}%���#!�^�t^7E��NF��8"�h4���58�Q����s���򾦒H���������;,a!�� ��x<�(�J݈{V��(8Յ�Q���9ډ��xW���g@����(r�Ƙr9ƖV�3���v��x�_4!���y%&
%��_�]���E��8�cq,���(�=k��p>$켸�۽��ya8��/����ȟs�`�R&���>���䫙L��F�G�F�'�^Z��x"�?m�U<�]#|Akk�&�Q,���G�b���c�*�3�u�����}ߍ`��(w�|$�Q��5�q4�פK��	t���7GQ�5�]
��,��M�Gȣ���Z<��$��]�"rc������E)p"��Z�s�����m���'zLk�Q&�2���o�R��1>�)�#42!��Q󑰑t���P������H���J<煱i�c��c��a^�x�=8B��t:}��z��p"�Ki��.r��s����>X�?It�Bq�o$Ѕ_����d26>dΜ9S{{{��s���BS��=�X��`�D���q#�]U�#�B��@H��q��֦ocW��h4�w�S��KFM~5x�?577���k�)��П!��#����P�?�>�t:���!Lg�w�כ*g:U�jG�G¦��x�aAJMwW��0�!����ya�y�G���e`�VA�9�<D�b��P_oĸ���|ڢٳg'po}��I�+6C��@E����Z^���QWf2��Oinn�q�����x/�Q"��t���X�N���i1(�^	t�煱p7:#v��]錨��_L��<�:�%�8�aQ�^�7�p]�pM���?	�pBq(��#�w#�ǰ�ߘ���S ̧C�]��?¼�Rˈ���þϮI��H�}8�5�״R?S���bD�"腑@%c�~��7�y>�m�k�s�՝�1����/H&��e�+�R��R�Nq�}�)2Ǫ�J�����|��r�����4`^�>�wۥY��c��4���nB�W��#a}9�E��NO��?�x�;H1�6>?ݽ�H���(	>�!/^6*n���;�I�&)�>ćq?>!���󻺺:�p�uF��:v�v��0ŧ�+��/��.� ��܅���40>�������	vk`�	9I����%�ON~�u�:~4����)Ǔ;�H���7V�+�}d�9	E���G@�_����}g�1�2�����l�ꌮjƐ
@t�~�G)l����u�d����M-�7��3!��>�_������K�ƶ�1E:��Ɉb����U	������ѱ���th��tۡ��I�E�H�8CW���h}z�hoo���Z^*�Q8?�����	t��f����Eކ�������4>&�HL����&������#��E(l��<�U��H:}N^cl��n�[���Ϳ%l誉q!q^[�O�ފ�����ۛ��.�F�W��{Ȉ��]*<�p��!�:�EG���1�+��G�Y��<C}hJ��J���M�H�իWo4>f���<?��5�L�[gN���{~���D��t���r��~N�e+�>>t�D��!�89�v5R�6��c__�	;�^����X,�$���u\?���ن�m�3f���"��0_G������5hF���ӿ�N&�����~�MMM'����1!�F�k=\����cЪ�"�g�A)"��F��G]����jE���K�\{a��G�Yz.�?��f/Q!�ʲn�:��>����/�.��s�n�d2?�r�h4zd,�>�&��}��X�뵫�g��n儾-���,����+�>vt�B
;�b�GK����s;�ɓ'+����~>	��X8Pw��\��ӳ�!vD��\���\.�]��& 477������Ia��Z�Rm�^������|F[8N"}l�*��bŹ��}�$6��냑]D�>�h:��0����o��q��B���pn��`�w���^5`���	|���<潙�
aך�qǇj�t�u��?��־�a{�._�0�!e�t�r/o%�&�h�Gv�v�tEӷ1���pk6���:B�	tQ
o�����~�*��<��y�q
`��*�??�!��+E�#�|��
t�/�k�ugA$�CJ�Ź���#ӟhv挿���4�M�q@��p��f'��m| �]���ߟ:u꿭\�2���	�G�Q<,y3���3�L �W�9s���1�^��b�5	
O[P�R�WI�_��n�`��Y	�����]s^�`�{(�&b�3��.��/�x�}-����lֈm�֍7n<B��t:}���P�(�.��Y��C�. & 455�qr)��s��2��B�V���~&?ݽ�Џ���H����z��0�XsN�Gq^l�4��7��E�&�Ѕ�"��Y��a���D�ѫ!ԯ���c\�d�0#�.v�{����c&���	���b̼�SM�Q�|��Gd����U����+st��0������x�jQ3�w	��Z+�>�=a�!�/���צR�%�"�`\��ֆ����n�m?����{�	��3���׌���%r����	�Jߪh�$��	)#���*��Q$��@������+D���hzA>�k��E�X쇸nmmmU��\?�{�-4�!�ั>�M�7��ecc���1��H�����(�H�V�&���G=��$Ι�^�CW�}/����%��<�M�!Ͱ1�^�����������{0�]=�l�=�%�L�dDSSS��b��g�t����@9E�Xwer�=Ey��R�h�演�܅B(��j���8�hm����n�5�B�V��7B�o0B
�yF���`���	�V��>�b���	yU�|5w^K�RnG��c����	ٝ�Dy�@9nD�)�X�ܰs�`�t�����ϋص��^P�<2p\����l6�0��Ǜ{zz�!���Z�֠���; �[M�@�������0�ZF5/�%ym�6q�#T*�|�ʠ'/ĸ!�	l��{UjoI�~a�&��S��2���H$��X,� ��k3��*#D�P%��C��}�ݍ����b�
on�R��͇���}��8Ux8[}\Q�����o���R�J��{uw��!�R8�ت�+�x��q,ح������X����4�_�}M*��o#D0�@&98��R�C����ں�����Gzzz�w"�1�}�mnô��Z���["��<'U�M5�XÊzHq+���O|O�:�BP�W23�/(�^܏j-�/u*�׬:eW�pܿE�;�?�A�t?���	 ---S0^}���w�FCQ���H�Of��7��b�H�����@/w1[E����lꎁcx����hk,���k׮�l�����n��4��G�/=�J��}&���l�<4Y�m�#�j�}M:�Hgv#(�2u�������[�@%Q���rt>R�H
�Wzc��/�����������w!�C ��A�)��$�������M���r|օ�����$;��r�Tb�X��T�NM�������*SY�q��R:��y����r fR(�^��f���N�I_j��8�t�Mܳ���l�W��'_
�4�L>?��H�D��d|�q����j�x�D:#��n��O��7��G]3������h��\��� ���hߊ�w��߅��Vk{���8����t:��P̖:�����p�1*��{~/¬�^
6���~�x�k�_�*�W	t������8[W�5�#���P�Wrɠ�hz��5l1��!�����5�L�4Bx���@���_�-������utt�����6���W`Ǚ��N��m���/ʈu�"��w���{�qGY����(��5���	t�P[[�ُ���7����$�݅��,T�j����3:�y�ϡ}�T*���hze� ��e
q�_F��
�?�����cM$�g@���۞F�	E����"��4ub�*&V�S�ӯ��4���m0$�=ķ��yr��ҩ�nuZ���;c�ʟ%q l1�[,*�A�d2��Q]$�݅�{��W�����p�B���-�(g�\~k(j�O蛾��;�g"��4�Q]��ŷ�(b�z�Jm��k�F�bg�Ey�u�4i�`$]�g���7�}�F����~��ӳ�Qa ��*4�	��D�_���>�jeX��P��45�?6�ޯ�cA]��3fl^�f��#��WJ���2m�ڃT���p߮M�)�^*�Q�H$�x<~?����R�?!*Ɣ���k��҆g��m�ym��ڒ�dgX����y��Mظq�\�3q�>m䣎F�U����G�r�rD���(+V���b����S_aJ���Îާ��v���h��L�{���x��!�����s�O�F�M�)(�;;;ی(�x<>��4��eg�N�����>�[�lQpc��i���h5C�1�Aѕ_|�m�11�Z
v+0���hzY����}}}���8���/�6+��5n�E�Δ�*Nrq��3�~���jW����6	n�6��4G��3b�Чa�DQ��b#��
�j���Xe|*�9�͵2�D���w�2�n+�K�{M�H�>���4���pm7@�?��槙L�i5�W����7�Pm���w7Ƃ.�Ʊ����3R�h3�u���vF����8���Z26�%'����]�.�>\�U&`�s���N�3|n���vH�ޅ�x��W4�,L�}	�����h�b��C����!J�U
B�K�)�k��߷���i'q�'O��Y�r���T\��Y�f���E���Nv1�d5֗U$}8x$�E�����W�4�Vƍ�=Ye�|��s��{E�+Bl!�υ�z�{a�i��/藙~@�߆���^����Ox�^^��}#�ӦM[+��(ʛ�����h4z^����Z��b#����`�p�{�	t�mWL@���آH�z�b2����:C�ȹ���aצk�)+\��-��e��h�T*p�(+���k�)��R�Tsk]N��[�_C��ioo�`�/�wZQ�qG�����p5�_^�o�t�mtpٕ	�"�N����u}�� `�q �L/�;�[�㿣�Q��bg5���#�һ���@�X\�����?�����bз>������D6m��8���ƿ[{Kb;x0R����}�)�Q�O��� 6;T������&�H�{q���_h�`;7���P�CGĦ�A�\ؕ��W�z	���Yggg`2{�{$��;q�ӈP��Ҳ�֭[�D����B�"��e5#��&=�~�2@$нo�@	�Jbg�%���+�+5�#��W48�WA��b��9������3h�!Dhhll�T__�i��M��M1����jf�	1�H���m�֔�vT���fC�Q0P��8��xq4]�ǟD��N;����ի7!D�H$����1h�D�±������+�O*u;b��Z� "��1���+��U]E q\��r��W�]� ���^���i�������#��%x���<�E�is��8�����lÐ��ߘ���c����b��y�cB�S��M������l�_�oq�_�r��SA��*D�hll�=����X��O��FTE�E)�Q��׸�	tR[[{n:	�1"q.M�,rl!��l<�#����^�L&Y�;�%�H4����g�)�G�/�kk%�����-��^�H�wuu=k�z����r,{�1*��D�t�S��鲟`M.�A�����x^�uttt!DYq�&ߟ���18�8�h�gP�\�'zlḀ�$�������%�G�M3��F��}kj�����@��}+�>������FQ2�{C���ah	?b���ނ�r(��Èr���PЧ-1F=�G������وaH��*����1���W#��np�u
�e���N��o!Ĩ0B�gg_4����C�G�ύ����J@����/��Y�J�V� #��Q����a�ͅF��s1vm:g����^꾎�����U���r|��f2�UF���J��x|�Cpzx4=��ny?7»���0�X%D%�O�{�"=H�Y��	8R9���	���#Q!1t���J�t_C��-����;�����7ΗC�<�ז�R����	A�Dcoo�Gp�������WV���B�E�(���	� ��?`��)�pL�F�,#7�<��`צs@R4=L�8�<M��C��<�+��
��?uww�B;g��!��͛�q�F֝�8��As���]��>F���6�W� ��}���iB�])-L��k�E��	v�)N�D�ѷ)�)���
�T*���c�>e%��p����@��̓m�i�?����P��[1���'�G�'�1ϥ��_�j���`���E&�P�O��,Q<�x�ص���K�]`��;?�:&Bo��<^{����_�y�_nmmՌ��---Sz{{�C�s�#�)��1C[L8�p�kW��bo9�})�r,��ؿ�\�.�����K�����{oQCC�)fh��P!q.܀�����"4L����H��>غuk�=�SV�?{����d2�ʀ<+1N�ϟY�n�^ds!B����r���<u�^��~j�O!���]���Ϙ� ��0���/��y�	���-��Z�j8�����̬�F� ܹ��U�ƪ���+3g�l[�b��s�{���#�HK]]�^�W>�{e��}Vo#��B�oe��KM��@�	�d�����BI��B��s!��F�{{{M�L�}�c��+k֬�po�)�~[����~�⽭��+��t������nN�����n�9ƥ�L6+�%ą��`ܽ���g�	�>����l����� �"��p�Vz��t1
,��!Ƕ	2��h4��ށ�6�v�6x���X�z�F#<��9sf�����f�Z:,�6~Lk�w9�I�!D�@��t:�؄	t�������7�fh���AqΪ�BT
�I�&F�Q�H���ս��l�ۼ� �7�^JC�u��	��9�M
��7�p�D"ѐ��f�9�����L3T���,�Fy���.���;��~!��j�>#�L>�~n�M��8Ղvm����E&C �b�>����6D<�Y������k�p������h����{c�ĉ��g�{��ٻ�Z| �^����#�����x���"|׼�k�B�
�|�R�-�>dʔ)�nܸ�`4?j���E�Q4]T	v|QǶmE��%'�x:Qy����6��F���p����m����{�����-�=�|���l#�;��d�χ`�'F�>�x���˃˱��4�g��)8��y����2ǩx��Sx4C����F�m_{�h���B��S��S&�H����+Wr��	h.�5�C��g�[��q�h9�W~�(M��J{e�ٮI~�=ɏسm�?�!2ҽ��L ��E2F�}�熿�V���o�}^�1�o���B!�	Ɔ2�̷L��@�)�T*G�(��������:iL-�)���I�b��{
F,��.B�#�BT�e'N<c �;�H��������q�����F�rEr����B!���X__Bkkk����@�9�d�O�'Bh=f��2
!�B!�_x-���ֶ�	�  ���X,�)4)ҧ!�B!��>+����M�R���>�7���x�����_��=_�B!�«�����s�1��؆z�H&�+��!�l��8��!�B!��x��4�9�z�hoo�3g�G{{{���F!�B!��U�6�N_�j텐@ �W��XSSsr4]����&!�B!���\.wj&�YnDA$�����Y7����h>���F!�B!*��$gB��iĨH��d2����q�H$r	N/3��!�B!*C�����8D�$�C@OO�555�WWWw����B!�B��/�)t�?��iE͋@=Dd2�U555�@���ӫОm�B!��=���r�@{�و��@Nj���K ���	�}�B!�B�h���W���g�7�!����!<HC�����q�#�B!�c���Q��J�^0�d$�C�#��͚5k����S�f
���!�B!F�9�=}}}�����5�5$��6���^�aQMM��MMM��xΏ��5B!�B����Lc�ΩT�Ո� �.��D��I$����G�u������M4B!�B� ��U��A,���]Q��eG]�����s� jfΜ�D"{A�Ӛ��T��G�ў�b�B!�^#�}#|�Mho�q3�o@���r���g�A��7�*H���q*�w:�#�B!��d$ЅB!�B �.�B!�Bx��7w���-�d    IEND�B`�PK
     $s�[��C�I  I  /   images/627fe4d2-0152-4b97-938d-4b9176d7a483.png�PNG

   IHDR   d   S   i��A   	pHYs  A  Ak!T�   tEXtSoftware www.inkscape.org��<  �IDATx���U�u��0<��y#�W|E�b�M�5V��6�������Sc�hMl�1I�G���51jbk5IU���F06A"UE�	�0�83�c�a�������s�=�{��~]߷�{�9���^{=����7`��ɦ��ǿT+8Qp���
{w򅱬��1���z�B��O?$8=����8��}����8<�}�1A��'�s�ۥ��r����C���O��ÇM�~��._�
��54���u~www�D�
t����wK 8�Np�`�`���"�>����0�mۛ�~�3v�	�_���r�u��R��3\�g&�@]]������_9��Ѓf!=j|I�E�u��	6K��%��� 8Dp��$�Y��
��#86���F�7hР�8y'΁�	絋��'�U������uMxQ�Cͤ���ꊈ4��^&���1v���C[��@�[p��s�fm �s��y���f������Q;!�rK`\ ���͡C���&�ǂ�'k�ȭi���y���}������g"
� b����|Bp�I�?f�l-8��C�S���b��竂���/c�}�������L�7��O�3����\�`~����N�jC��+��rD��$��f�w�Q�gq��H�~k7v�R���XL�so0V� �]�q��e�o��]"ߗ
�zX	��~0�&}� �q��'�5�S�52+AJ
�`���r`~'E	hY�d��'�%����K��p!�"���D�(��?%�Y�q>#���%�	����-HDc��S�uttDc�Qv���� ���@2�<��Cs0$
���*��4n�\�P����N�/����
n�5c�!S� !�pH}���6?%���|�Up�_X��0�>1�eT�;�H��~�=dȐh��L@�3�>�`���zfWða�v�{�ƍ�˭Ok�1��36g� T;�T�4�*�E�{�7+��J���I?�I�����	��P�R��*���ݣG��b^-?뛛�omii�$�8/�3�˂�͏$.��#��0�,�	�A�@����1��O��q 1mY�bOVE<��t�҆�����,!�b�U���ۯ*c��D�@�Ϗ)S��-[��k��Mu���Qx��#��F��!��\Ey�T%��BL��|�c`�|�-�lr��?'��`S�=q�����8S���/�D�rW
�,�wq�)�,P�X��3���X/�{3�A��1.4�X}B�,Vtm۶M�Yp��%t�.�r"R-(��_�Q~�+x\X^��<P��`��:{`mt�n�{���}F� -��3�}�TF�Ǔn̛7���է�P7jԨ�{������v�?q0|�y�*�!��|�`��=\�x�9�����C)f0��0I��X ?�/,X������4�]xekk��q^����	FO�
A�4�� �#� �ϭ��"�������3g�M�6�nz�f��Y�S����2nܸ!��A�뽂��b�e�p���-�8DT���4�'YEWE�E�#0��&oV����� ��9�FP��E�������f":��y��k@Q��B,B|��	��o֊�F9��]$U�*���lM����O�� ��ޒRn{���Ks>|�� %Q���o�䎎�C2����P����a�cC�K�^�UAQE,�G�����8P-��a��w��%�MNb<.3|�����4����|�'�\&�xF��V�>*�*�����ͥ�^�+
��x������5/��r���2p�0�	�qG�2{�V*��	&���/��M4�ս�bM	w|9�
��]�W��`�/�ҠAtQ�a�k{<�%�@TUCo��"��]�n�{�tV�E,(O�M����E�"!J�z�!,(�����2T���@���I�,�K
����MG�	��̾��ZU�����<y���s�obz�9��2]@��Sf��?��}�m߾�O�/���Z"��j���Cc�"�M��IVWn�0�@l0VnF�=��E���Y�_"��&a�4'\&��W���{�d o�s�|��Y��_��kiiQ�L?N��FV �&V3�׋IAH�J����������H/"�;Y�F13��<���2�mӦMC���"�f�PF����i��7���755�?Q��h'�z�޿���5�d��l�^}����I�&�k�@8B^�7�����X�a!s��':�h���뎝;w*q�ٻf�?� z�5� [��o7v�J�J���_�=����4��x�c�E�Z*�#�r����666�'��Ῐ�7����`�}2�|3�:�g��S� �6���g)a12+a�?2v-39O蜥^�~UpP����o׆�5 �I�f���} �����}���YwY@	��TWI}ɵ32V5��D�"��s�<?!$@�Θ`�L:�b�]�
!��P��X�gJH�~)&�_�㵒L�
�hӀ4 ,�>�4�n^������[u�@�_�%��,j��9�L�:��͛7�Q6����e��@���u���* i�������U��"!� �K�ڵ�T 
��M�6��-�2��.�p	6:��mG�9GO0vB�O*�� *C��]xX�p�8l���w�c�-�e���r�D��1�|f��*��f�	
W]ƿ���������zIN�GB�y��+���lv�X��&�yR������$3�*��s?ق�Gj���M��a,�l;׸��N��!T6�X+���ٕ�^�QD
��B.�����^��!$����;�i!��g���A������L�X�%+����E�(�=�P�̒�r�X�&�B�u�$�����Դ_���ls샆�p�Dd|b�D1��������OV���9��e���ث�Ʀp��
ΪnY`�M`b�56-	O���'��� A����J�"	�Q-B��!q)DY#ˍe���fo�����I��!��W8C��VWlJT�t��y������-��
��Xfv'$B�c������u�<"qr�=���[$�r�b2�rc��z���"�M���2y�VT�9��6lX���w�G��39 JL3f�Y�zu���YZ]Ie�z��s��5���2�{SA;����BC�i����on�ԩSu	7�ayCB���Ŧ �HWID�rVqf}�A�ys�M^����S���	10]��1�F���PF��ɚ	Y���M-G�V$�j��B�e�Tͼ�{V%�� B�g8d;��4����J"�qH8(Z�цH�5G�� W������<�C��è�<;$�#H��ˍ=���IKͱ�]�:��fAG�śBd������@D���At��'v�9��~���o���Y��_0v� �.�"��W�c��Gc��Z�`�w��!��,��+�� ';˅,B8�M1�).)����f_ɇ����g�!i���K��'	 �r�o�W���dEh�D� Ib�ƾ�c	�{*�8��������z\�����i7��3?cB�`��=����I@�P̕����$e�j�%��"Z�LG�,.S���+zJ�b�F�Sɣ�Fp@1�m.F��9J�am1��r��$9`a@�����⸩���z^��֮]۫`@�\���lm^@��s���M�ِE�[ӀX�g�+T� g��������c�ql�z�?��=�q�6`�)�ω�`��z�^�\�5�ё��Ϧ�%����EB62�l�o�z�8����n�EI������VnWR/���*�������ȭwĈ��N��UQ�ó����*�JJ��Y͌�L����E9bx��:2��,"�p�}��� ±y�L��o��� �X��E��PS9�TM��ⴂE	5ֻٰ�.�R�ܪ�r�#����p.����~z����:t�۷o%��XeX1i&9��F�'nӏ;��	�ۄ�?[I��ِlV:.�`Q���XXQ��q�)�DIN<�%-71<?dȐ�tvv;R����V��B!���0駶8�a��O����y\�	v
<��p%�C{4_�L�Ę;wn�\FQ#F�@��r[Ȇ|�7�#577�ٳgG�ۺu���A�e�g�X������\�2~�x�6�Z)�9�\c�_�(��L��L�� ����u�dV���;�q�t�4���K����E��q�~�)�&�Q���!�3�Mr�����w�!)w�1��fp��?	@R::r����>��� b���e����(Z�9g�+���,�P�F��q��utJ��8�m���vD�s!�ľ�^*�C�Y�'Z�.ܒ9�FS�@�Q	!7A�%Rcu�礡rއ� f>J�"��H��y XE*ǲ����y�G�<�_�7�\c<x��H��F�]?hР�ك��I�
�V��0�Yed�K�"��t�*�@t�e��G��'��=R��]r�V���+����l�C�� v��p�"�\l��U������Q�w7:nY���K(�3^X��&8�w��{R��)XR�]"�Q>Sk���o ��Y�����d=�"~�w�H���/w655�����Fyk�u���!�*�`�$(���<sD��$Q�,i"xL��+��2T���J	�?K/-�1��	��lժU*�XGG�ÊA�����-_4V���`�RVO�. �"�a�g<)��G���{!
l}���M/R�3�B@�UI��u���� K�;` ����9;�0�~L��K� �〔����}��n����5����!r�r������Y͌#
�������ߩ����J��(�/1BQU�KJI*rgk��yԨ�!]]}䎞���<Y��5v��PI��`;3��2���pPduA���2����E8�pv�=GV�e��ұ�*͓�r#J�����ڶ��/��/j��o +F'N�Â��ޒ���t�ia�� 9�!�� )����刣=@y�Z��=��v3�>�_*3�N�eVF�hA5|�BHƜ1N�a�EoE8��g�k83Ɣ�7���[]��_�>X���o{^`v�t���]I�>�Cp`��Nu�ݙ��4���	�Ń߰{�nD��~%pF�7�a̱�鐾Lk����+����~B�|Ѓ�P�QP����]�CX3��y�$��ve���YQ�:�Y&P�~A��1>���K�3@��Uro�|_V�����!�Dx��%����d����55�B�ڤwM%3��B��*��]��v:��ń���th��)� 'e9�&��{D�%��,�*�G� 7�����zC�I_�]*�Dw�9|��Ƭ�x���Ms��Ɖ��W/����4
1Ȓ��݄(�<ĩB��;d9����b���d�x�4�����m۶�<s�̗:::NOz=�B���LT"�h2�<�?��pa���p���`89�>wn�K�"�-q�!�sF������b�8��C�Nj;v�g�3N�ed���a�{GD�bq�a�{��:��}R���#}J<�(y:����Mc�B���:b��$	;�#C�Pw����j��A�gI�G��&�,�mH�ަ�B
E7���I�
�����I(%X��g$��i��i@p�/�!�p�W�=���1���u�&�����m�__`9A��)�:�����jڪ���C�ꦯ~J{�E&O]de����=�S���eM�3{�}M����Ʀ���nu�(#�&����� ! i?��ܻ�y$���#t���ߥ��qqi'(�e���{�[�|��;�3G_&pyJ�ǩk�����U�Y����u ����+4
]�Hð��`q
{F9�]��}�ɞ�"�(L\�
����?g%�9�¯�K�T�Ǝ��w�� l}�t�H)���l��kG�v,i"��G؃��w8��>���$LF�~��#Jc7���r�.A�ϥ/݌���PPV���KAB=�_�%�+T����Z�n�,�rѓ���1�6�Db��2��GXRE$�e��Z��:�5��:Y�_�K�����}�Gd�b�"�������,�P٪��M Xn�C�9~A�<J���z^:���ۢ	��~�_ �p�,4eN��3�}��}ǔer��C�<A��GD��x!z�Nk��HE`��3o�8�4�M ���A��_��k�=d�8"%sB�[pT��?O�@g ��o�3���.8�b�W    IEND�B`�PK
     $s�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     $s�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     $s�[y�E�wf  wf  /   images/6a97e33c-aa93-4e7b-a2bd-349ce97096b8.png�PNG

   IHDR   �  F   p���   gAMA  ���a   	pHYs  �  ��o�d  fIDATx���$Gu �Yտ��;��_��h@B^K6Z/,��5�kV�فY;���]�y��v�5�#��Y����#�3�1����ŀ�Ќf4�;����wNf���Y��u��͖�{�;�]]]u*������4M�.���»��w_y��u׽���s��������x�Ew���}���p���ַ��iz=|��݇���n j�ZI�Z��j�^Ǎ+/�:�����B;M���ןh_�|yV�i��s�#G��776k������4M��2M��w:x�6�-�;�n�^�uV�^m4f�V�U۷�����Z9t�P��g��;v,�|�觉�{���Z��j��v{f�����=�	�9�g����gT&y��?�����ŋ�k6�1�,LZ3�������0�})%Nf
��q�$��s⤟����l��R��2�	�ŕ��Oәn��DR6R){�^���5�q΅ߧ@02IE�_����~%I������Z�����S���N��7;;�N �.�ܢ��u�LT���ʝ�c-�{�6���\G�/^Z�i4�ϝ;7S�Vڽ^���v{@45$V�7�q(�D
~i/������+W���z��7�o\�|y/~^[^��l�;{�
x&���5.�@�)�]�S��
ު�ʁ6����w�Fc�Ա'����|�O��O
=�A���_��߸��V�y�ٳ�^���z`e�j��

�֫�w�u��5�i���w`��p��$�o&J�I��4�Tb��^�Սp��}T�<���p~/����P�Gq7�Q�6��Q5����40�~��4[����LOQW���� 7�� u���$< 6�!a$q	�q
�q� ���@Ը����:��o`� ᩇ�i%�['���U:�"`\Ҵ��_K��"A�&��Ե�H��Z��k�{�����0V�X(ݙ��gN�^k4g_�җ�טi|ҥ}�C�#�8ѽ�-oy�3g����v������0 {�+$*�J�Z	j%�q�#���`<�=8p0��S�<|_U���f ��	�Qǡ�!9�� �F �P���J���x�00��&a��yUZG*��`z��� ~��W�k��/��7D�pC��1I��(�
$� ��E"�W���J�d)��h�g��U"���и�\�<�++pFgcc�0��0�=���������޽{/�|��馛���w����M;Bt��{�O��<��-���Hp���`�" 0$3�b5� V��c���CM,���Us�=��z��t�?�'X]�@U��(��jH��`F��_�H	/u_M�2����F���ϧ�K�ϕ.t���;~�����{�׌=>]K�{�� �T��$IWVV�<uann�Ү��Ξ={������뮻����o��o���F���/��˿��/�H� �&@�$ = �X��T��%���@�s����5Ԩ��s0So';�c�9� �a��)�ǿf�,�Y�h�M���$5}C,���mRM��3�jbx��S�vΏ�3րs���7=��Ր��F=�z���w��y0�?���7����=�z��^��WW�>�g��'क#��~������6��w�}�;}��̀�IPTo����%Џf��P���p�JF`��p�@���5ǉh�H M($�M��(�+�i�稱��Ĺ���{-�������^�:i��El�Ζ�z��O�_j��
�0�k�_�� ?=ϝ�K�w���M��0�:�z�%�O�Y��i\e{����n����/�gQ�Dtw�u�O��t���捰"^ v`nn� � U���J�]60��K��lv�&���4���!�U� �Ԉ7}�t��4AH�:x.
�D���Zl��s�QDƮ�����=�9F:ft?)�n%��b�+.���х���O}F5��d�ÁJ5�sunmm�`�Ӿe~Ϟ+����`$ѽ�o�Y����u=���p9Z���P
��Pv�9D�K����
�EJG���>:�TH��.Q�{�	����T��Fzri���پn��YxO~��=@u �lŹ���j��ΘSW���I�"J/���*T��鈍��ƹ���[��D�����S�N�n�o�b�n$)לȊ'�%8:	��:��ʯ���)�4�Lf���	�}o���Q���G�����5}cDWe ��[R_�@��?ķ�.���q���	/��.�uUb�I����}�Itp�6�f3���	�����⌠w$��L�$1�]���ƥ�^>�p@�ޭ��;�!�h;Y�X_��zoti��g��!�j]�����b0�耫��������_��6�΋U.��hM�^�1&�.(�D���c'z�I���?Q0���ɧ'�W�����T��K�_Wd�&R���DlFF �`h�[MY]�G�?����t�����H�'���E>�!�&��@n�"=N/dr�h�DWI%I,��,Y�V��e�z�R��[��H��Pm��+�\������*��<�&�����?1@i�g9�����I{��E\z�s"tH�
 �6�
��퀚�v�k#�*�([��D733�Î@�v :DV�>��~�=(Y�����}"3n�W���Iٟl�/��B*��D��R���1̀��&��8I�j��;3,���`VMm+�ItgϞm�Z�
�1�0��e\�[�yg�u� a6���f�U_��t�\���sj��<|w���%����D�JB#H{�Z 5�J#e��3mvڵ�׮T�'�՝��?{��uʈW�L�Hp�M����b	����z�vGY��6A'1�(� �P��L�.�����|v����Xe�M��(z{��Z�}�ێ�H�K�/QDח�z�[�+bqv�t�a�@m�H1¨v��(
��5�n�n����0rˋ�T�����s��b��3O����X���1i�u��ư��u��Q#��D<�ƵJ')m��$: 4L��R�����V�e?`Z�����|i�����[�2���Ax\� 'S�+�y��F���V,XZv�Q#�!̜� �K[���Օ�����t 
}����Y�Pd��@��E��i$�onkg���D*���8����I_bD�
��H�g�QH1N��S�^ܽ�����hF��R 8=[@}���Q)=(#��СCկ}�k�ڍ٫�ȹ�Ӑ� r6�?;�n)�Ȅ�IDƣ��*��������}�O���4�Z���PMڪ��'�H�H����bd�V��Fm���F݅�_��ׁܫ�1�7�j?�z�l��6W������\/7ƞ�T"�ɞK�-�{y�{��ó��+��K��viӸL����t�$V��48�U\$o�o(�ǝ\F�FG}'�p�Z��A|θ��0�M�*:o�b�`Q8�@t=��f�^^]�E�ٲ�It�Ν��j�>^����Պ3>6�a≉�
�2�Ȃ6�;��/r��7�=B�I���aQ�r7�C7L�'��nRM�\�������j+LaNM�&Cpk\��'V��
R����2��|�ħ3G|g���q@"��0\o+�M���+�\?/��q��r���LsؖQ��,�#�ncc3K�X�J�y�v3q�|/D��Q ���T2�����5D��Р�N�g\+��Dq�6Lo�a��M�*PGHC��0N�QD�U���B #Mf�J��I<����z9���)l�(#���v��$#��F<�a�Oy�=c�H��YD�E��9�o˒�L^]��O2$[�뙯1�(���veq/�ĉ���v�nEc���m(�C�7���%1�y�s�!���x���#����b������#Lj��(�t}���L�8��"��8�$���9���ZБ����� �L�sa>k�-#8��1'(o˻&	�Ļm�cz'8������j�����<ݢ�d��O��{�[:ӤLDS���:��H��ԉ"�c��)Z���ȄO5��9��A�S���&Tv�m�!��ᰥ��N j�P21p;�ME"׌z��R�1>�����t���t��%
���TۋY��6�Ќj�`8r1Sȟ�CR";���~�[��#>�۩�)2 �N��1*im�����۾�W#CA
#�K���D�*�lh�N{�Ww�،���aR!� WR��������D�\A�{�1 #�A�v�7rtڹ.��+ZQ�ж���x�J���� e^o�j*�!.g	��l�p��g�`�C�gj�U��S���o��(�R�"��+EP�#n3Ђ6�'�F.�\Wf.S�U]]]�!����m�Ca���%�!"!s���2֬�*��Ǉ��Əb�ONJ�vXN��P��&H�ɡ�i��6~:���xFX�b�Z�u>��%���ە.CIt`<`aN]'x#mHD,C81b�>[s~Ce�D��%f'����鬈��]ũ5*���b���dVD�c��U̭J�.�9�9�t�?$>�^���mM���백$��\|I���`H�ɵ���Tf�҈X�J8R���@}t���W)�=�d�$���uӰ���u
.=f�}r��p�m	�YڪA4:ʠ�������tIj#�ȘƗ�y�ҥ&v�ƃ��J��	 Sn;K3�4U�Wd��j�G�Lٓ�w�Y�)��:j��`|HX�v��8�����,��x5w,'��b�䱦���E�2�~f�ũ��?�Q�U\5bė�C�Q\�Z�(�1���Ȍɝ����?5�PtF:�WC�^I���`M���o����M^L�h�������{�OW�2��>MH��ٜ��en1�g$�����������&V�������3C�/�A�aRO	��,9��X"<�Y�d�K�ѳ�v-�w���u��гkkk�^���Ux#��`|��N\�}�^��Hq�v��hO�V��g���Y�~G)��`$����mCl�$��ѳ�-�gY��p �_��
�T"г� �}��^¿�͍��%q���$�k�IW׷�*%�>Df-���v���^��)�|��*�� ��iG�c��_4��Ū3\��(�B�Q)��v���ȉ�U���}�� ���O�;x�`��O|;��Z�,Ҫ$a`�+������j���pSZuB�d\qόXŀ{�,pv��m�&��X�M�7�~,qS_L*�mG���B��5�Wl�l61uE�K2d��)\ǰ��hc��&ĥ��WT��D���BW��5#Ӱe��%5Fr�!"������S�����?�!lL'��j��:�������A�g����%�E��!Rk@`/$8�	*�;�V9���5w�F[��t�P�n�C!Ks���U�&+�қ��o]�|_��X7�J|��ۅ�)A��.�Eō�r�(OM���HU>7�*�-)ɺE
�r�?�^������.������)�o|v�I|����t0�N1���h��u��o�@������~�Τ`�.�m��Ս�X#r�<�r��C]�,,	e��1met��~ZӖ�mc�S����e(8,^=y$��Pg�h^�Kx�)0�6%j��.��_� T�F�4(K�����`@(Z뙟��8��͋x���Km����OG�Ex�G&�]�+�8�}L�n� ��~0�
�TI�oYdZ���D���VI���lun�'K�l�Փ�x�djBX��F?�!�\ ���d��F e��_l�$[ȭ�`�>�y��������z���؂;�Q��V�M\���RZ�����%z��y�1�W��
�=�r�2 �1Q�ִ�f72�¨i��j�{*�t�Na ���tm��={s�fI4���v������l9�G�RS�&��@n*vE� ���r�m����Bt=�jY���P�Zej$�>�];V&�� ��gb�/�|�\-����s��݅Щ��0���&�t��.�i���z����
���x4��+gd�}�4C/#��������Ms4��v�*�t.��IgwA�>��D��Wz��iu��iY�E8DF���\��J$�1H���1��%�� ����m<#)��yqY���ӵ1āш-�K��+�����Xo���U-j1�G̐�R� �V��c�Tz�$P2Z��8v�e{�b3�'2C!5�*�> Q\�������/?�чG�6��?^_^^�ln6g�T��Vgc�gx����J$����wMa�$���p�D�'Y���&6c��	������la������;#&ӌ�ȋ�����{m��.�2�0��.^���u{1 ,us�����	�����'*�	�l�R
t
�~��!)�.5���)���m�7�F�G1�"�7r�r�H�e�<�K��{�����?r�'G]�L���nw��Ɯ��D�Iu��=D��y�j�T��o�D����}�4:�Ό��|�����~����3e�0�^�U"���|��^(���ոT��ȓ67[=��P�[�waJ�$�'x��}��q*�&ոjS�����l	���9fӟ���4p��H��)����[�FX�7�ֿ
t�v�n���!�Z�^�ln*�o����>��|+\�D��-"U9���0�7w���fk��w/�Y����S�٨������ghI�d'$(��z)�=��VW�v�(�#ޘq�nuf�^�b^ ��`�=|�]=e�R����yO�Jt�u���*A�~�����D�ͥ)k��԰z����j���4f�^�_�R
W�#�D!%WC~�W�i�%n)�>b��;D�+Mp��h��#9�F�E�c\��(����(vi)_])lZ�J���OAZp̃���3g�͓�>��pv}��2��9��]��C���de�q��_��r=����EtJ-JgZ�V���设 ��Nb���$�Bj�J�u %��D�b��8/U�U��`R\N=I�E�� ?����
N	"+҉L{65�[�4q�-\}���q7�N��)�D��N��Ctڭ�,vⴹm�|a$O������D�-��Δ:r��9X�.V���z�(���Az�&�0<�^ƅ2��*0���Z}<�Dk��1Q�I�&2�
hJp9�:Fj�~Sjyύ���@).�7α"��h<i��D_^�朮l����3�&������\��ã��*�.�l�����1�y��6��xLUq��1��N*cb$�$�qo_}����+x\�u;��n9H���L�Q�m�V�Tw!+l�?WmԺe�S�FB&�u�/�IO��r[9��b?Q��1����h��L�K��{5xM�WpH���p0J�iN���I�!�0v��˨�no�;�Ra#���ի3�t�f�H��BjOl����>&��7�h(՗�pW)l��,��<q?�H�K	μ�N�z<�R�wwC�F� [$V��+R%�@�s���st��J����5ja�X��fH�b ��梓7���2#,Kx���Y�+8 P>���E�E�oX�7,�5�_*3�:�nw<�ncc�(��Nw6�{r
"�b�3�����6�Ė�^��Y���^�;	�II�tU׆E66��*]�=�Y ��A hR�hJ�%Q�9܆�R�y[�P��,^E�����Lt�=#>�AJ���v'���ƶ�5�Y�[p�3�7��J�f" ���j-QfD�E�^�q�(�,��Q��I��
�!�&<��@pY��SA^ `/��������ER��������ܮ�J�SN�	��/�)\�.��j	(�V����e��y�t�..�)6�CJa�Am%�/��9��=�Y�+8dIt��./Y+�,(�7�k�$Xp��'�w���ŋ��(q��$|�N� =��d�bh&�������\*
�}�n"��N��3�X6p=*�Ѫ�t�b@l�� �g"���Q137;N�j�ڸW �G�N�����fz�@��w��F�IJ�6e�Op!�����T�8D00I�)Y���j�ۨU����H���Ϋ�J\o<���h���j��t�T�����D�b@].���CPP:Ͳ�7��-�]+uh���K�<NH3�r����VvJ9�J%�XZ�6�I�Q'Y��N�N�	p�H����������{��kuݾ*I�lvv�E$k�j>g ف�cx����G|����T�9ʜ��xo���=�Fa�H��Z-�0�薖�jgϞU5�����
a�^��S��D��j���:AH�T���q��-�r;,��\׳����4�M�hid�NG��:��F%Ե�o�ϔb<�,�.��g��fv	����m���2Gcv�ъS�n�?c N#�;u��[��e�!���H�O�&䎢�&)���{q�A�A-+:�v�R(��p{U��t�jHM�(��	Ք�)%Ԓ"�¨DZn�|�7�����dy.�\X�,��9�qF�P~:�0vK�Qo�+�}o}u�~o<a0�n@s]�dx�ݲ"
�5�~�i�%T��;�2�x�=hٍ�؎�H$@��\o_Ҫ��Ff6���U�F��Z�@G$�<F�e<t�A��MiK*� ��i�$�2��)��JA�DJÁ?ꆩjs�͔����4�5�q����G���*��Ԍ����_���?�;���e�{X֪@�Y�JԁYO���O?��֞����
�3��xvV�il��l�d(�-��O2=Ќ���6�1g� G8�j���Y��q��F&�IY�Ҵ�%|¥%��b��ʧ�ɏe4S����2~�����3�����uWwzo���e��(B{̂+~h�cR״.M�o�,%�d�7&n!
.U�(0r��V�F�!箭�ۂC�����:���9�$��^w�|=^#2�R�$�ӣn�O���t:q�^oa'5ED�z@���	�j��1i�^j;u�'����ݮ��7�̩r�	N7 ʾ/��	n�h��QY�qH�;����r��k�������y��q8�>��@p	s��+ �I���e_B��W��=������R��ˮf��&��?5[P2<�P��F��b����5��uٱ���Ոl�PHT����Q��@4U�=Uп���cQF����M`͋�6SvV�L2� ��H�J2��"x���P�l�����lQ�&c��>4�}(�bi�^{;\���h�_9�����-�D,]+1M}9���m��^~*~.e�8C�Z��h	l�Z�2۴Qv�gx�� e�a�0z^�ʮ��Z2,2��Y�b�W�څP��7q���Z�Y1-i�����(��C@��ɠH��e2�|=��d\a���yt����T�������3qK�'h�F�Z%�a�գ�3���ܕ�HSɉ*5{`ۓEf�\��Z@x���[đ��v�;�6���t�Ό%�f����	eD��sS����P�v��μ(��k�ہ�רZ<��D%{5�Ð�F«�З�Ŵ@
�Т�zfХ��M���O��t�m����d�k��\B�
O�#mD��������Hl�4�O3&-��֣	�^��T�5a�
æ(���n��h4z�v[��|�P�ˍ ��~�F�Pb��x����a��8A�n����)$.�a"U8�=i�{IFt��ۓ�ad�!��RȾ��M�5L؃ �+��ҭع��N�e6���Y�`�O�Y��ki�ط���Ua��1L������ԎX�j���z�d���ԐH%��P��t8�u�xٌ���*���"Dp�<SJϓq�QnW��$�G0�����2n�Y����u^��W��ӟ��g���L�I��l��J�\/��Lս[�8�El^7s�"��g�pQ{5�7"Fi���9�c�&'����c�(I��641e^I�����Ws��N�E�|�[u�ѝ臙hTR�0
Te���`�D�"�ޟ��?'�!Q�+��T I;�MI�cuE3dtխ	;g�L:��S �/%�K�#MZ��پ"n�B|����G	pd�CjL�K��xZS��2��<=,�$m���L@�/1��N��*���\�>���S���Ώ�菾�/��/>>lx�]euu���M��]��vl��I�x9#��5�h��R�R�'J�twKM¡]��R��HjZ�����������Rl![��,<ÇC$��đ��D⓴8�b�>'$�)���X�q,��%E�׹�`ۉy�-2&�Sb�I0�i��Y�l�Gn�T��k�_2�q�T��2�ӕ��U���Ա�2P��b�䬛"�pH����Nol�ݝ�?�`�d������p�N���o��&|�U̳I���&��,~�}�tMIO��i�从z�H��;���P8�J�U��)�f�
�2�N���1֏��]��[��ӕ�1�z��i�7�ӫ+��OdF��S-�`VVVD��U�+�jcB'�	��ƹ�4Ħ��f���u��������'�D�L_�����<��2M��s������)�D��JZp�`S�bh1��򢊽��f�J�e���	45yvH�rq��Ez7	�Kj�J�u��D��O����%�b�')��2Du>W$Z���(�r�#677u��Z��*�4y��D�%	#so��&�b��������1
��Fy�ӡ��\��U��hg��-e��b�(+<"-sk;�$����j���~R�Ȼ�&Mr�1��{�k�j��8:���>;��C\\UI�4x���HQ�ȤD��D�b��*�v�vYh�0���"�AQ�jobe����>�[ �)Q�5T�R�L~��'�����b�Y�q@H	�Z�E�d�7�%���ЋF�Yf��vb�/*��M�$ʈS=�yeY$�����g-Sn 9 3�.b��3D�%��;�)�*m��v:m���0q�9�4-y�s�$�\1&y�W�V���#��ʕ+	�rL�T<�C���HZ�)�k]���D����|:��j�3�V�+B[[[3i뚋����Hq>�����I�N��O/
���ˈ
�.�7���.�!��3Nx�6���l��7
��[t��"��e��v"��84�(W6�Wh�D�qϞ�����+�ȅ�ǎ��*������M_��z�jgj=
��O�}�\"�T��l^;�ۻwo���^�x[���Қ��������;�<�ضI�Á�ՠ���Z�. �S�V�PY�T����v;� f"�%B�%�i�2{%VQ����l#7)��+��UX:�f\>���\�\8B�[���,u8��!s}ې_�F��x+\e�h�"���5N�u���Aq78���ӈ��m�T9��l�6�G�]m��&�V����u�	� �m@n�n����AWr���USyԳ�-ݪJ^�t(ÐP���|[H�c�,/���u�V�N+T�j�Fxs�vA�Hyb(�f:����5 (�E��̬)�4�6b�nj�'US�9��=��6�e.�t �<3��U)�M��
)��6Lϥ��Ԍ]*��uK��*d+0�?#P�`$�z-�KM����}���I(M�S�� �A��j�l-Q�0	���ڍ�W��alv��j�>�Hd�ZE=|$c3h��В��c�ڔMP�i��p�pC�2�	��J�� �D����M���s\��*Um3�&о!*�Pk0�U_�VS}����9H�FQSO�4���Ca"��F� 8Gv�?`�+E}	,Q�z7�F��p���`�^�waA��ݫ2��/�3�a�6,�I���7�e+g�;l���5gL}jI����2=��9EMLгb�ȁ`b���U�R���f���z�ffg��B�eT�Ѡ��I� "���uq��e�����S�EK�va7��d�YK̊U�+>}�;��r��)�jE���g~^m��&>/��'�A�<t�������L&��K�WD�^�|�o��O�V"4��!,������%K�0��c�h��7� :$�~G����������<���ܜX][��X��������<��z ��-�h0�Ȕ2@�<8Ǳ����k��F��9|��YXA) �\'Hlhz�CQT�cLΖ��4���ǎ/zы���\�ˤkes]���r�Y�����OZ<��Êh��-�,��rj��x\N��RPc�	����������[���^3�^�{� �+@d3������bfnF��ܯ�x��y�"��?�G񝧞�9BO���Rgl��ׯ6��W�/��[i3��h]���v%�����������Kb��>5���=��A��ϋ�{�Ңӝ�o�|�K�S�NE�<�?�Ӻ������1�'���:�P\%i�����O���]�~f�97;�&��e�X���^
�%�-Y�P��!���"ʻ�[��mo'O����:�(^Q��&��g���aϞ=�����յ���Dr��3t�<�2��¶0��l�|`O=�B��'#�5@\�*q�����aa��='z�ސ���������e���CM(��4��/���ĭ�����c�]��\�*'�*��W�:)�g��a���d$kpϝ�Av�y����:�I��jm��k���  <L�=�n}�*��^P+ R�J ��ʃj�⾌>$�..�>r���v�;Ɉ���m������c��MxƆ���1��O�`�� �6���a��.���~㚉nqqtS���_��3(F·,MeL�3a2���q|E�'�D�©�����@pJ�/_���E��ƺ�l�3�E����y ��n��x�o^ٳ0���hq���ݕ�4V�Ц0�N�Op��FFn��U���Bk�|�%�0��F���,� ���b�=���W6��&��N[KQ���P��;]��Y����֕���G>������
c��+WbIz��'P�I�(\
ʯl�XQc&0�-�������o����u\/W��J &����"�P"��C�H`��Ꜩԁ�a����,Bu�����}��h�2?�ʄ�Jand�Y�7fZ�K���>y�7���g�������O<t���;�|�ɇ�6a$с��8P�������&P��x�l��a��9����*n�� ��.�x.Mz�������}-+G�(�ʅR3���5P�7W���b6H��~����׾�1Pb�����#�F�~���`DvA�m�ml �]�<��S�?~�-7���G�L�Ay����ۤ����V
��3 ���F�+��sl2_��^���c�?�Gb����w�Z��v��Z=q$���������%�����/~ɋ�:���	_����Za$ѽ�=���� ������}���%� eD��\[]S�"�����~W5��;����|��n��[!8�ǎ=��X��Z�0�v&VP\�u\�pq�'�" 8x�S��=����ܬDC.�MN��i���#�۝�^��Rű����}��/}��t
�]��(���b�=J5gt@uX�7��IO� ���i��%���"h�(��%����V�76�L���<y�����d�x���R�;��8]��� h�+�1��ow��p���o��w�|�O��nG�q�w���,X�>y�߬����ן|�ܹs�ߣ��P*�M��@��p��r��v �� ��=U�G����A
�s �%X�_��{�V�^]Q��k�^0�C)�>�"\�t�R�J�q Z���,b��̊�U�D�P^�{Ao<77����k��E�I�����B0�j@��u�7۠�%&ԤB`&+�
�Aqx�:X����Tt�pKp��&Y�;�x2�b9��YA��Q�{~��bz��:H�lo�1��zAu+K/W��XȎ�@̧�J���ݻ
��f�� �5բ����/��x�����t�z�ω�%	`�C<�	0M�����$CG�b�K_u�c!$�{T�Հ��9�(���8��G�otu�jPu�CP�N�Rt�E/�+e�p�r�JP8Z��BP�P)<��QkjH}�[YYY?r�H�q��V���E������?2�m� (�%̿@5�����! �i����_�9˸ °�A�D^�DQ�m�G�X��s���'��\��W���`r�n�����)-������z�X8p�9���˹��ܰU�Hddm�&���3"`�0����$]����':0��>%�8�|!���@�N6��0�� ��t����TQ�GpԵ�s�䄐�7|��~����\&�bB��Y��O�&�?�=�'^/\�Pj��qA�R��$W�	�������N�O�r��0�9�0�vBڐ�OO+Y\$�HW����Ç�� p%&��Μ�7��'F`����#���x:�t0@���U�w���╾o�+I��t�4I��↪ FWH��u�ݾ�Er��jQM�7�0:��#hP��K@:'HP�C����)�A	�:���랔�
t��J�UNu>��'F��D����鈽���M,���O�Xɉ�Į/���*�k�q#���,'B��ЮG)*)�G�iNG�����s �^��,K>�c)�N�8ԃ�Y��c��	E�?�s�159�s��� +�8�9s�y�M7�I@p��n��>�6�E�IC�t�k����s�z5lx	���YÜ�KKK��I�0 Jl����J��RU�q /�ز���Dl��!�?�hN��n�����N'���c!8�� (�J�o���D�t�,G&�,m��"�x���,@�����D�����p:�K2��w�Z[�ݧc�F#�dg�HG�EW0��;d�;�����I�<ڃ���t�O�7�|��':$�6)r�p��DtewX��*7$��H�'x��';�]w]0<�~m<?���L��w����88LB���\�t)�N���/t:�a7n�E!X\\:��8r���!$g;�n)&��JW*��`�fӕ����/��� p���)�:������W#���!�$���l�������&��Qv������\�r%��+`EG�g�W���A=��g��W��  Q��+�"���`�9�K$
x�+V�s NT9r䯞z�!'�I�=ǟV�D���>����a)�ӑ��@NW�=�$�X� :]a��N�����Z[[�	��U�$���p^�4 ��y���8Μ9�v�mb0	N�ď�!8���U��ؓ���)W�|-R@�+�+���aQ�q�7-�T]�|"��U�*���N�:<�,�f�!"|��h"�g���	������FK����s��BAp��<5?��'N>|xF��vS7b���?�}�v�Ԑ�E�,F��N�$��ŋ��zBS.�A���O<��$2]{ւ��#�JE/��|� A����		E���x��Q���3���-���w��F�@p��lk%t�i]�s��ť�V6%�b�S�Np]�t=�`Ο�0<��t�B��`�O���9�b.�8 �BBäӽ���B)
/]]�z�Ҿ%
 ��j��7�}M��к.���^�TL &�=�*�fe�"`r��"i�#�Z��5l_	���XJ�B��"B��Ν{�����}����!p���@xO���x���C������>Z����a���ʼ��HW2
��z�Q������������o�P(\���n�����ѣG_	8���?��3���{�wK]@��O�~m���!X����|˟������\��X����y�-������/}�K������?�������Ba8`���)F#N�<��c}�;��A8��n��;�����߾r�=d������y�3}?;;������>������-7~0o����W���!?�
�ї,@��?v�X�yX�Cw�#�o��8�w���
������gy����|���8�����{�k^�#b�0Q�&�v�s俿�%.�$�d�[M�o�D�x/��+�� nw���)J�2��2�<=�C������a� �(�0m�g*(�Gp�)��l��0��;�}�K_z�[`��0�;�yu/�=��!�xV��9{��~�8~�[��/0��� "���2Lj$��Fၨ�#���x�sh��Y���a�I]4�a�~�/��/���~��>:.<����\�.�;BU�'�xҩ��8������{��: �|>��q�ŏF�4,�A4�v�R��ȫ��1Bt �P{!��ߠ�>��ǁ 8ȝ��k�x�=���:�w�0\�j0N|�}�hl�<.�8�<��u#�(j�_	ȅR�+7H�`ǉ�'���_�Cƨ{�DV�=��D��~��u�C�6�����_Dw>i��ʹy�&jkP�<K��|��gŘ p�������l���&�1S���y �'�Kjǉ��>�����݅q[\��oxY"���={vlet&g�(p�*nW9�ű	3	a6�4;V��ς�Dns���g������/jz._]��Z���8����QC@}-=J[B�+�ޓ�?� ���Ǐ�H ��R~�$mX����V�6��l��u���^[F����ĉ�B'���0������7;Nt ��pEvX�W`��<���|��w�c,xNX�[1�-'��&l�j���Ia��	����T+._�<��p��'��k;��_(����F��n�ZVm��D��)�}�IA�ٮ��KE\������6�|px,�{���,��:�;?��x��W���!z?Y�8�sG��+�@���&����h������"�J�Z������u4�{���':����'c�;6ҵ]�,�8���R��?Elf�ཋ~�_�3��I| ���s�;�,Wt֋@��L�A��%���zk��>�Ĺ!C��JS{�q��@�~�Dl��G�pN76.���R{��z�0D At���%o�{�%�b·
777O��8VNǛ�����5�		M��D��kaR-\�rylxb��L��29��yА�`ǉN�N���7���]����h�`�r&���!NR�Y]kU�V�w�aii�ظ�ù��cʏ�g�~O=����� :g�pe�Hx����"Cbmmm�^��t���;a~��r�r�8jo�G@�X����?��܏����N�0��ϡ�D�
΁OxR���N0�@�D�?h|�r���a�����Y���$Fտ��J�F�8/�V�V7�|�جl l'
�Gp|W��p�Eb!ئ�!��a�(&�9<(8���̻�#�%;n�m�w���XM)��.1�H��*Eq��"/^Zc�4u�1<�ϳ_|?'����ؾdqqlh���}V�����g�w�G,�S��p-��){�G���+�D�ddEW.�cD���^ �y�ѱqd��Q)pqP�w�o�_������ :V�V��<��׽�u;����
�v�0�;Ǹ�E]�W5<xp�^t����&5�G4-�Ř�?�*j7nRА��*\&�2'�s����|�wP���_ĶZ���`w��ߔ�٭�r��wqBX^^kk�Җ�J/ŭ8��.��Ǌ���u��U\_0p��~��������1��,b�X�%�q㬠��?{=�*KKKA��':99��_����A���K����]B�͍,1R��Ձ~)67�:�!�Kf����B��M��X��`�j��?^�6�q��@��X�E�"�b ��M�#��}����;J�X���SN^�!
��Pj�PD���Z��¾���?��?~B�n��T`,���	�ʟ=W�7�k9��{�'�8p�-����	gt)�L�!�+�O�����?���!�66�DJ?S�$�n0������>�J�&YسX����_?��~�k��k!<�z��(��7����5��~�����ǖ�G~D�4�8�q����H� (J�A��W���=��3֒9����݀y���'pZ
�1�du�������_�՜E�]�ۿ���� ��:�+B��<�������?��#�<�|代�YN�!�ߨ�Ф�{p9|�c_��W �{ϸq�s�,�/�1�Nc�%��~���:���+_������w�Xl�]{~^,��b��@���������~�3���"�8с��`��nuu�Mt��!�k>�8@���СC�[����/zыvdE����g�yS��z��в=i��P������0ן̇~�o�~�����3���!�뮻�7O�>=��>V(��R�3w�#<�裿��|�O��v�A����k�Z��_� ��BE�h>�Ey_������i� �U���`R�}I�(����x�N�|�+y��'������27܎nw���_;u�Tt���,Zg����oS�����^��׾�DhBt�A�'��:�y ��`���kH|�A8�C�sO�y�#?�������ȑ#�{��ǻ ���ؔ�����LO_|!\�|�s_��?�����Z��o|7��A������L@�}��M1!V�+�~x�����z'L�[A9�A|$.�%=�o���٧�j���n���K� �����"�T��/j�u�ܹ�w��]
W�'O������t;�6�Y��%�x���Ή'���g�b��sQ,`Y"��8�@�A{�¢X�Ɓ$�lΜ��x��᜵�� �V��
�2E��e�� �3���7�Ӊj�ħ�ފ�\�X�D��r�2[@hҮ=�8�3�&'��B�s�X��! 1{o�ߩ���VVV&�NW�D�,�Yt�� |em�
DW����đp䠍�r�m?���P�E,S؇�݁>z�ҥ��{�Hp��G! �%����P��^o���Rb�Zc��k��8�����ν��N��ޫWx��4X�6�柹�M�v�Y__/���Ap|C:���`� JP5�ä���D��H�dC�U`��6���!%) ΔI����A����_����xE:��\&Bt��6�	��Ժ�|vE�spN�]� GglxM)q�����]�����Aɱ>��:]�&̺��ŋF����'m��� ��bsCč��S�On�����hs^�UKp�����'�$`"D�ӹ/�~�G����.��b�ķi2o��Lf�F4�o��%�+�|:��`L��K�$�""�{Y��9;;Tl�Q\��M$6 ���bP+pq$ Oe�9�>���׿ޟ��7R��D��'��U��}���dx#â6\W�^���:�������o�}Rg2DW�Ex���
�BoS���'����,��Z����KQ(4�>� ��t�We�%8�~�!J���ѣGCo�f�~Zč�]�'p;�ҝâ��(
o�&Bt@PvB�"$ ���Ow��ŉ�
���
�=�)(GN�v���}W����lN��T�K1����	Vfh\�J@�0Պ's�F��S�Μ93�RH<	�x��E�(�<�c�&Bt���LH9�M�.���;q��m%?��p��ؠ�����%EbP�g�W )G�C�u?��Z�=��/&�]�)�'q�Z4F,D�e�Њr��� �a"D����`Zo����@�L&e�p�#'�����(�Lxv	��n���qlnnN̒���@Y���;����o߾�D�.��� ����+++c�3�$����`��B�O<\c>]I�16p3@D��ʜ��x��NW���}�U�G�5�����O;�Ŝ9�QRP�%Rp ���+&㕖��t<�G(::���u ��;^��͓8���COf�I"�:I�"���skP	��&
�ٵ~FYW�\	�W�Yw��u�vNAc���-i,�AIA]�שׂ���K�Ug-'��h�s�B�"|�'��>�"',Ln�*+�)��X��Q�:FN8`j��L����}%C���>=�+�Wr�W<݊G(8����LG�S6τ�WK0*�m��ä�Ι>84��b9������`���@���ɥ�&.�b����UV<!��|���Ͼ�d�8]�:�``��Q@�Au�,��?_�t	��π{P��oŉ@��_��L`qL���C7��e���A��)X��ZK��w��Ю�
�-ֳ.S��6':PW�+"!X\���G������U�a����r����G��v�r:�0���_	g_ �l���y�5|�X�XZZ
��ǹ�r
��H|\�\\\9�cĴO8-�<���'��t�p�h�֑�c�9O?�!�XE�/�	�	@�?���(�3U���0)NgW'r�7��zx�ܹ�:ul" w	o�S�hB�y�r:�(ܯ������w	��tV��r�;"!�+�Lx�A�^]O��>;\���N��iB�L�Ϥ�p ��@�k��I�L�H�b�KQD��_��ל�^�G����A���q��!��C���SW�#XG$�8rG�Tx~!l &-��x**�#����9����r�����<>�����L|��_dM �7��!�=�3�A�ĕ��t�`,֏��xNW�+L����v���*�+(��# �����p
����s"<s�����OG"n@�F����k��A��PD���o���K^�`8��{~18N"Z��/qCG��~�����?�p<�4�r���s�+j5mb&�"���o�����7$�z�Mh�������������'�%uL�Ҍ�d��Y�T�&!�Ud�������`ŉE�R�H_"X�����;�����"<���_�3��
��t� X.B}A�RD_9q�DP�+��J��4/!Pp��}= ��6qv�1��S�	����L�����D��Gz�UПy&�=�=7=@�q�6w����!���Eۨ��0u�8a��N�y^~{U���̠�YГ�/����� n�!u:��6��p�@���IE$���Ć��/9,��:]��r:$r5�@��6rd���
���s?�s/�{ޓ��u'��t����xܧ+�	&ʮNTni�H�}q�r�7ݦ)��5=�;���'q;v�������RDp~>,���&�eRg�-�`}Kr�9�O�n�q��p􉎷j���s��QW�^���O��]��P <s�^s�@��|<8�犅���a�^?�?��� �/���QK3��&	Ep`�=�?s˕� _}�'t���p�9�
�d��哹�����9O�������% g�5���GQ�&X�S�OgW����B�#!����i� �<z2������[�PdH`9�`Ra0�}\���r������5,
/�1�O:]pp�&Ա�tNߐ �e�8]��pz��9i��+��^����3�R���YB:�So����M�����
��o^����J����ڂ��\
4��/�W�{��z�����xE�ߑ�7$��秋�Z�V�zދ_�VfЬ�i��lq����<�9���y��w���O}*�9��|1��ؠL�sDT��%��9�ЩM~��G�U �*ܽj& �av��! �55���w�����@�K���������t��P�%!�l\_�[س�y�+_y�g>���ڙQ�"BQK39m���R��� > ����Ƙ;���J~�+|73)�C�41>�Ec
:�t%q������-��.C0��588�ӕ��%��3r���������;��;�	 Jć80q8?U,�vR&{�q:�.�W�^C����:q�6RH��s���M�����^E��0�.�&/��UH���8�RŐ�ד"�9� ��y����C�P�L0\�⟑�Qckރ� �H�6�&��%�0�s�}�BwW�uC*J��c�؂+�!4�����|:�Cp���t ��'�:��~gϞ����*֊�tN�0�����������=� ��=�p�DY�{�K��6��E�}��B��N�� �\ ���{-$�!��\��P ��JW����<�E	��!�k�!�ؠ%����R�+W�t��ַ������ J��m�q<�Va�Zu�z��#ItQ&nL��� ��!���E.袕3g�LL_�8�����Nn��I�8�}$h�8���<��3AS�`�
k$Hg"+��W,
��l\A���ĉꩧ^������V��ɓ'���	�*��3i`|��6���"g��p� ��Y��~��'��E��Ԕ�f���A�&�2�{������H�Z��~%_0��� 5 �or��a�~=����}���|�"$L*��Z��:Mߙy��ׇ޵/7s��
����KG�������!�.z��D��{�`R��S<�(�� t���+,�O���������*��Y�D� ����/1����wI��I�2qf��s�S�E��k���+�c� �~��뮻���7�����?��!e��ߓ��1]�a�=�T?��Ҿ}�����g�gr�^zE����f#$�!�N� ����|	|N���8]a0�#(:��IP��n����t�666�柹���.��%�b���O��+����;D��`��"rd�&5�����t���r[oR�(��&6� ���}��ŋ��Si���^=0�!N������ח�k��#�0��&�1I����|�W�^Z9b����9��� �)��mo{�����`��26�C�҂�8	7��N�s��F�[ZE��	B�t����?�"�\5���s�i�$8���k­�ɍ �(h�IU��U�M|���z�>�w��{�� G��IAE��� b��I��v?�����o�0��Q�����~/j��!�_	t��|���4�D��������[����4�E�G����`�.�қ8�>}:����]�1�
x'΂������Ͼ�w�w?!���E�U\�E:'��^a�}��g�m2|�С�m@�{��8O�.�?�ِ��1k��)�CE9>�]�p�w�-��I�d��i� ���M_�\��ƃ=H���رc�9s�f�����r��fo��_�{��{��ƊJ�K�F�4���Γ(���غ���%�:ȼ�b���?�y�h�p����g '*��W�|!8p`�R���+{�+�R?lS�׃��>�%�%��Z��9 ��/��/����~��E8p�2�c���"��,�|t���! D��/�wˇ���ꗿ��\��V(6�!��#޼K�W��֭��*&ot��-U�~U�
��t���]ɵ� ��A%��/}i��zk�������ѣG�K���+/�#'�om�ٳ'�_	���s$)���$l���N�裏����<�[�X���ŋ��� r���z� �s�� �"��4,
9q B��{��DH ���t����^ח7�t�t�t���x알	L���O���z{��?�p�H�Z��7����{4X�")��ө?������t~�&Z��M�0���]�%!7*�,+:~�xЌ���ć��sd�yS�yI�~?��z;M� ���ͣ�=������A��ۢp"4L���i�ԹL�gF���0���������?s�0��80v����"���4�q~:�t�2��8���3����u����Ξ=�f��(�f94����fPU�'qb
oU�P{N7]��:������G�Nb�yg�
R�s��l6����
�E@���'�_K�d��`�}�J��c�=&1H�I��&����w�A9�ߍ�! ��ɦkkkSW��p:�8Tvi"qbq����M�ڲ
���;(e�a�]�z�'C"��]�yy$�+�&�WY��t%q
OlQ.�2ġ^�O��ى�S�IQ��}j�e/{٫>��υ�[}�g�P8�Z�a&����y` MWa�����0�b�	5|�����&���$0�!^vp0�u*'�������LW���c��PmoF 
zp\S��:q5޹ɜ�95����������Px½��ɚ~,�h�5 ©+�qdU�� k�Á�z�&;i�(˄���>����^�
�yjSQJ���U�(<��B�Q�i+3��L)BD��k��_}�mB��1�F���m+E�o߾�����-.
��`?���R�0X�Q���	����7&���E��>d��� ��^}��W���`"�;�����"�(\��H?v<ty_.��HQ�빹���2�~%�L�8�o�h4Bw�D(�X�#a��s�t��G�T�\"���Z���9]:��e�BA��&8���L^�G�B�9�@��ɓ��%�8��y|L����tE$ �$m���ו`�/A�銀z%m��E��u�]g�]4J�F��Q��DSĕ���m�B¤�`UX�N����OB�sVߢ�h�7ԟN�8���t:����:�xӥ����8���IE	P|����Q�Xx~�&BA��8u�TP�����K��1,���¤*��ϊ ���s`%��}!8ܕWZ�����Z�
�t"$ ^�¸.7���1�.CBx���q��\��>WB��:��\�\~�t��#�<Zt9b�;�U����t�A���\��O"��(�<��[�`XT�FP�_*�ۄ�n
ǃ�	&U#�8O��*���zH���A���t܇XԵi���P������&��7��z���?Lf��B�iC>ǫT+�(A�/-5�D�g~aa!��x�J^G�w���L����T_WZ^^�9��v(��3�}O?(�Z�^���c��f״P|n��.N�Q�W�q8r�Hp\}=���%��� ����M&yq�q<]I�H��@Y&>\�|9�_	p�e8s\��{m�Z+��i�I?q�;���ʞ���~�Y?oWZ����N��ӕ|��pl����aCvҝG�n<s؇��q���Q������DZo8��]�޴`2���?$��NG�9���q��E�9�	��L|��&�2s�SL瀑 ��:��Gxx��]QǄ�Km^�:��B�S�x7�I�I���h2�}���ٹ��[�E@H��ƥy�&��������+��ߗ�Zr������=1�~yyYqb]��r�íN�:�9�g<1�Ju'�>!Յ��駟�~��|��<+6/�@:Wxqe�Tp�|�I�v��[HQ0�|n;v,�#�i�Nָ (UݯZ[ZZ��bk�����<���2��L����Gb�_�Z��|��������0~���":d� �aR�~��kΐ�m������t�#�t��ᢂp����o�9(��};�g�1��q߿�=��ˡaR���})��D�?��H�<5�[�� �Á"]A��y�+����w�T�+��S�i�A
2]'џ��I�[_�����:Q���`�g����9�y�t��&3�3�*��I$�!1�����Q"2�.�ߛp�O=�TPN�}��gʣ#\��H �5��s��$e��W$:�V�D7�]EA�Fč���6Y�a�����k^ПȻ&�۷o�:q�9�s��k?�t����@P��Le��U�c%З��	8X��:&o��;���t&��@֏��<+�~{��$c��Do>�A����AU��@��ǭ d7��׉(���<yrKzO�
+��w�}߱�߽���!����W�s����x<+�6��t�.��Bp�%�]�D��a��v!8��.�]�ۅ�Kt�v�n��.��Bp�%�]�D��a��v!8��.�]�ۅ�Kt�v�n��.��Bp�%�]�D��a��v!8��.�]�ۅ�Kt�v�n��.��Bp��cr�6�|    IEND�B`�PK
     $s�[Ɛ�~<  <  /   images/e65d6d59-bd1f-4659-a32c-fe6c1b0070ef.png�PNG

   IHDR   d   �   9ty   gAMA  ���a   	pHYs  �  ��o�d  ;�IDATx��}�%eu��W�s_�m�Iw��A�h�DQ$����(1q2�,��k\fMLt�8c�%Y�NV�BL�ɬ���D�@F$0*J$#����@74�o��9U���{W�S��sOrf��p��S�����~�W�	oy�[��Ԕy�gL�&I�y�����yӹ�>��陙�V��6� M�hll��w�n�^�M:K�l��1�Ld���R�,u;�Yc'�ƢN�㌍�5S����G�v+i��)~��vb��P_/������	C�G���&��hzʹq��ܱ9K�jE62ݤ�辈^'R��բ[���Z��OiL���xk���!���R���q�Y��&&��q���╯�{��Agbbt�I�޺u+�en��U��@��G?jN;�4��/�fh������/��/�����'�V���^���U�<���W=:�>M�݇E�"YB�G�s.B��ƿ$���.�]�8ZI,(-��"Z3ס����h �$BX�-&�o_\\��<�q�o(�]����A ĤI�&"�0��!d��Cm�����Iw��vi��̷[��b\B���ݿwowjr��Vk���v~��_���^�v��{6mJ>�,���0��Ч_�ݻv����{D���>�z���O�������-s���cǎ�E����7����W��u�~m���G��J;w�&I�e����6]�ۢ��2��{�������xl��y���"dƦ�{��GT�ۏ�zJc�B������a�8�Z�f��D�?�ir������8j��O���Ng�(f�;v�|��̈́��3�3���ٳ�>?��7������p��]r��~�ۮ�A��G�e�_`~�?ty�\w�u�+_����6sss�駟6��s�y�;�y�s�=��r��]�.��׾v��%tϺ4u�$!�# ��F�ς�D�,��,/�_$޵)/����-D����'� �b>��ฑ���o�ǀ$��o���w�Aӊb��n���B-!褣G��E�<��Ni~b�޽Gv<�c�կ���N�}tz͚}t�Cc�����;�

��k�m��f�O�;�ü�5�y�ƍϿ��.�]~&Mp=�@�l���'he�ؕ�0~Ie��{�K�/�(�9P�a�<�/�Q�t�eMD�?�潆>B������s���蟰�R���Gp��f�'�ј�,,,���;�ҙ(�2I��8p��N�kɹ���o�f�j��|��_��ċ߿}��7.��)�N�����we�\�3����"2���Y���!iߚi�p��MN�tgz��g�J�1Y����寁 �;w�S� �<�N�͘Yoh4������ݩ������w�;�y�r��@k������z�9�s��U�=Da�b�+^�e��He�]�2ȜK�,�k��О�vA1���q�l����gl+6����O?k�|�ʮ�� $,�;�k���!o�(�5~�M�}J�gSMU����-�A��m�0�h@�^.�Կ�@�-ߎb�hb�6n�zvX�\�����\�=����{�ڼP�NR?����Jrْ_{!�zPp��3�0�抠})65x���G�9:��[ݣ�+�- ��0�
[�G4#�y�Q�=�	�����*��VL��g^\A~?'�r��&\c%
��mt�{�.M���?m���W�[@Y����>'\:��'5[�&�]LM�&^�۸ȋsHMƮ,K�VfY�%����3�No0�����jwoK�L��%.�і����]l��Wi�*>WT�W�OL�kWaJlC�A�[���Z�ds�UV�E�-˫��e�/T�R��"�o,�f�k�hv���:���
0Ɩ1�P�ڄX��@(
�ͭ�*���B��U��@:SE��A,&m��+�V�6+v��"̴�, 㹵�v����pYS�	�|βrVeL�@��I����ԥ�[�����^j�����?��ˎ�����+�5�m�� Z�t@�Q�G�"2H`%��+��}�)�&0�*Uw9{��v�u�k@L��jMl+!d,%]�3ݣsQwq���J��;+*o�p0�@�L^�2o- ��{9(�lj�=��UV��5��V��}i�(-�n�!G�D�6cG��AZ=�B�a������W����gU6PL�걘���f��a��Yʋ�)͚:�'�R�/4��-�k��a��R=�BD��=�1�J���@��d�W�ګm�aΙ"B^;��J��]ڟ5�E,����!Pu�E� �*qNMZ+�j?�0���m�n�:Ѱ�ؙ^����c,0��[�+iYZ%��ڨ�� Q7~u�O�u�ϽW���l�n�
	l�S��s'ܪ7��/ڰl��үY�$M���b[�Zd����~�W
u�|$�����Vk?������z�blFMi݈hd�J��姙��f��ꛐ��ԗ�|�ߣ߷	�c��Y@|Q���I'FbDx�U�Fc�a���A�:D���F�n=u�c�U|7��<e�iŭ,ě�����1m�|UP@!"\l�"�k��u9vF>aQI[������	���L���ѹBm+t�ڗ=��U
u+��&�- ����q7*A!��������Iа�<���E�M�*s8��e�w�+��<�a�M�����|�B�%n�ɱ�_]�p��W�lnh#�(N�hi�2D�)l���A@�.
�2%�1`y-311��ۅ�hc�h��k
kS�h���|l�	8d��lC��+m��a����oD!�0�$Z�k1�Sz�;%�<�0����%� �����$6�영wX�Lycd/QA.�ܞ�����ZmgT+Ңa�^�5�M��k`�XXXhD!"CH-�r�P���a 2|�eAT�����&^��J��l�!��}��.��gKT0���ex_���ʣ��[����QÁ(D���v��^�����O�<!."�������<��:�c5הG7��PMl��A�r7jZf�{�rX"d�PI��!�N��XS�������1LX�Ԯ��rw;T�ISh����j����Q闦
�������R;����6~�����!��4��nK_h׻�M��4�a���>�@U��?����$l�+iY=w�����&Ě%OQ�YW����>�����D�
(#%������n �.Bjk꓊i�s�z�$3�;<�/��:���_�LQ:��Mr�g2�"�Z��rz����b�Fky�,v�`��}�T�f��:19�{��$����a�'hYq�%6��芈ql��L��>�L���V�:j�������1s���]��B�>d�:t�{~s����8V���1�S�=9��99�C������8�˧o�'�ĺ�)����[cx�}���R�BN9���a�77w�dB�W�#Q������`<�<&��"yfoQ�;ś�fT�ϔR�S��1~��'��q~�FYz*�!8F�&�1��)���Bz
�"X�M�J�{ģ��Ě �s��D��_@�X�l���2dF�6K���U��M?�3?������ʿ-����jE��	�X@�T%�y�D�ƭ�J,K�l@���|`������@LpR�B1�~U^V�;���8ޑv�"��4�y�����B��_д)��zuA=�b�)�(M`E����E��9`C��OD׌$s:9Ū�k�`�u+��T�@����NA���P%�\Z0|�X��9?ž����}�#D-��ߕ���G�+h���#����\����t>$ؙ���G�e�W�2��=��yH
�32���ld$��byTIU}Db昤�Z��$MW��n�����bk��Q��B�D��A^o~V$�}v�����+�?U%Q<�׻̺�w�����XL�)ҥ_I��/�}@��^���h��������>��"����!�!�G~�A�5��[�c��'�F�: .w�s \G�dFbh���v��;E���
$4��%i�(Dvwf	��[����ِj�۩��� ��h 6H\p#��*�i��I�s3��dG���L47���B� ,-.F��*ͩD��r7Y���[6t�d��i�T�eF )`�	+3~�fz>���"8(
Ð��ցÇc��4�0��.:�lI%�~�i`��}4�*R���_��e�]~j����
H�aA���i8>��o���wH"��oZ��.�
��c�#��,�4n�H�>�-��� ��
>��N{�ˊ
���Ei��_V�Ϭ�!��!��Y1^7�G�J����Ĉ�4�BN>�d���N:��Փ_�O����X��`]Yv[����Y��
`+>��9���S��W}t<��P�5F�r{�u��d��T8���6������g 6�;T#E���NX���FT�W܈��F�\�\Da�ß���*����q��V��x�w�U.|�QN_A'4����|�~�T�H�"���2�2K�U�!���l��u�ȇ!���'p��!$�g�kO��.um�Y��%�P�K���J��p[\ZG�#��-к,dU��i곴���Z����2��pu���,M�rj����	����:|X��J���a��	�n[���m�~J���H�]��(n�G��VUghpp���y�r�B�[#�-�Y�?��:�	*>}k�Թ��;�%|�w�u���f�I�̰)
��q&*��?���*''�rCP_K�<�ٙ����u�Ԯ�e<x�Sȑ#G��3�F�W����E̬$��5X��D�8�,��Sri�5�g�X����*'`�#�!�����XV���u!�J��N�+~R)ԅ2�Jz��U�%>��X'#�?�P}��	+X�3�ڧev��5���ij�7Q?HU�0?���Sް&�H Ň�SG�q��8�[@��G�ʓJ{��LI *�F����+%�.eK�ɍJ7
��͜� ��eE|�J_d<M6�3�dN���Z����a�w���B�Į�t%��aOO�\�'�,�8iN��<֫�^3�\��5��"哇�,Dh"DhlɔY�:d,YD�p�����C�Ŝ��V��1K���,
!���w�*'+�BԶH&2wt�S��[�J���gFV��=�Q��{+,K������b��;I������W�vJ�S�0��E+�DB$�W�x��������rHu3+ջ��Ÿ$K���ȩU+h�jh��2H�OIYӇo���G�ۆ��V��qj�X���+�33�s�}�!�e�$h��פ+iY�$֤��WlK�򆤸���W�G�R7�����p?'��r/ϲw+�'zoj�hR��!g�,2?�m
�"®]֢��T-h?WJ����N!���- j.�T���㳬E��;�����IF� $?+q^R�.�
5&�E2?� 2�.�Wz�y�ȇ\?q<�a6�g���o<��N��?�S��ύ���~C��Φ��3F�v�~�zo�\z�)�E�!�����v/v�ݓ���6	׹zW��"[e;�t��%�M�"տ2D��3݀m��/��[��|y%��#]V��l~��fR(>��+�:/CKF'�wr��i%�����5�f�X1W���@�I�g��P�LY%�>��$fqq>t@���[Ǚ(.�X�_�x�0$����c~dL�����ٖ��,��ޕ�1{����3'qѻ�Xpg�/����˂BB�Z�#圧�_36o�H�u��WΟI[����"B����_���/�+��y	��
A�-y"��A�瓦�<� T��ש?�����W��~S�h��LcR��s�0#�&b.1�ieK��Σ	.%cUE԰	�4#�pX�J��81��B���B��c�x�I�Mćes$��j�F�k����Y!J��'W嫗xv�X���.۴S��Ƒ��E<�ԇ*�i9ȧ�?E���ʻZ	ٙ�g2U8����}f!3_*[�t�SK7��$Iy�"�֌2n^t�XU�6���m�?�Ņ��t&>~c��'_q����n��uY(*=���֤&�;���D�G��&D�=B� �Β߽�7k!�޳)G��4�z�	�I�&Ԛ�슍O�L��?���_1�Hi���;��"�HW@B&�x(a�k�F
���΢�t�Y\��EP��[%�2ݱQ�@�y��<�q��!�����M˳��E��<5���Oݎ����쉴�K�c��Q� {eɓ���pl��r�qʩ�����(�j�2�#�h��� �ܴq��q�������|�)^��=�˙��е��SS����O7�6m6�7o6�֭�Sjtzz��<���_�"��	^�ڄ.��b��;#��ʌA����"�_� @v��f�4³A���m[����5^x!z��?�;��gbr��u��1���_��ݚ �L'J�,��� �,�y�{�E�\LH�;s�Ƶi�F/���-䭷��>�G�H8HDQ�<��F����ȪK%M�}���u"��3Gf�Y�6m���6�qRW1�#G�.�yǝ�k֜d�" �B*s�-���6	5��ӫ[(6=9ٝw��������~�lܸ��0��>|8B�)6d�å�Qӄ�(��y�{�����n�=Fj�Q�B��׬?�LՍ���s���G�z�m�O%D6�� ��v�/'�8N������I�q�;9>љO�;B@�7]���[��{�؜gKxȌ/t�^�q�y�U�Y����/�������8<��qD6/�h
^u�����x��[1q���x��������f�1H��:�'��b���y��_׭��3O�^NSX�6jŇ���4����	u��-3mZ�=03fK���z�frl�F�4��k��E~�D���D���n�M�M����~��}��ѣ~��d��!���a���z��+�|�'���w|u�X@�gIն۾�Pgaa)I:����5�u��8�̳ӹ�s�o��o~�G�������O>�Y�����_��;>&�
�i��:I��iÆ��W��woڼ���u˟q@Mυ��q8��ye�y�z��!�n��?i>�ٛ��=�m�;>���,,�W�k��f��z훮������o}�\a.%�2g�&C�up�iR߹U������ҁ�n���M�L|Y�]�YR'�y�+��+f���뉔qϑC�C�y�z�`��؜����[�n��m��!�9�Q�"�}�xָk�n��;������o�4x����Z�}�kM����/��$����9r��9g�xT|P���&hkAnE^�hO�3֞ᵲ��~�9��s������d7�Z1��X��?>?����f����7_����裏�R�mo�ȳT$�����ɾxΘ�|��ꋐ?��?���?3��{��^C;�77���s^�H���Z�{~���e�_n>���ج�E�6�#��]c1 ���hҠ�V;�\XZ��ۿ~���g߁U��}�v����v�O�ƢZe�ܾ���� �_��_6u�L]��y��|�3���ױؙ�<����N��,�NLN�a`�fm0TgH�^����X v�r,7�L��'���j�����~^�kp8�)n��K��Ƶ�2�ڭ``dt���.������4(R�`�����ͳ�w���?B�E��@C�x�/�ѥ1%�C"��3��E�Y6O�k�>���B*
�{f�iA+�y��lѓ�Tǖm��D� ?� �SI:�.�Z��>�d+�Wqg�q�IH�qb���.b�|�=��� ��įF�b"�m�84�Z&6�B�	ffYR��y�k_����:ݡ-<�3�`ȟ�%���ҚF����t}�"'h������fY ��h0c%B��P h;P�%s�E�h�����g��P���"�e��NR*��!��؏_$��ty!cYa�02Iv�N�=u��hv u_�A��!�����0Ќj@J���A��� k}@=Y)3c9`�ѥ6,��sd�$B���J�s��E���&��{R�-�a���F���p�B�F�/l��K�h> 6\A!�X�z�$m	r�������D\�%%�2�=:���j#d�ڵ̑C���?C��ZyJ���7oN8�G"���z_��yU�����*6�}�9���}��b����Y��߳}�9b�v��u�o+Zm����B�cTRF�/ ��K������|=Ů,>�*L �!#H�%C��9M�q�?���s��g�u~EAM�"d����G�5M@m�������֬�|굊aa��B ����cMU�N��vpo�v��g.�+trOЈ���v��Ѓ�;h�=��,�N�Q��C�����m+���W��r�JM���);������^�B�.��C8/	�]N���w���*QcP`��J��8�g�PV�1��j#��#�����		�n]���9��ygT��?R��|����3�����'Ôd � ɦM�|�T�˂�o*Jej��A�u�ֶm�|@�ښ��w�6��K��GM�n�:t_²$�#��U~3@S�C�I�t��!ȓ�ǎ�u�^ �bZ�E A���h'���,7�F��h�P�� a���	��P �l�̎���aH;��������/�|��xGv�}�z�"�7ܐ|�C6�������y�?/P(���V{�}����n�m��f���:Sj#�c0E���UZ4���G�:��ڱc�9��sW��?��?�=�����RT��G��e��r˥��z��׽�u�2ڞz�)�k�.󒗼	/KGh~�u�\��Hy�n߾}w��]���=��Sk�j!�;�&��K@��rn����i:!�n˫^��w�|���>x�+.5_�җ̵�^;P_<���F��b"����vI�����/�����7=��E��:'h�@-�6b{o"�F�}jǜ1/ ��j˖-��C��7����y��W׋��C��n֓F�6"��0������B���i�_{�e��f�M��k������i��N�����>D�c�p-����~5Q�EW\q\(7�y��G~�GV��o��H�� Q��P{�ċ-��(���;��?r����O��ij@m�E;�4�ߦ�mց���n�����7��ڳ����{�UW]����Gc�i7���WiA.�w���ޣ �^��d��W�w�y7�u�]+΅��o��۷���{�_/� � ��E�q
m�ɺZ����	ki���m�$����+�kH��OT��J��1�]���Bȸ"��z�|�g�'���o\O�^�/���ώ��]Mm�Dr�5[�1q�%�����A-�������4��J�O�'���� �?���&j����٨x�O�L�OG�Ք���O<�#ĵ�jr��{�����Y���D��y�֯[?��ZΈ��p�4d�Q�rAH��h�����v�Z�YO��D���ӄk :#�	BRx���߿��e������ZmJ�� zs����3/"�2�� D��5R�F�	�%��wv9@��fhq����L�8�u"O)�'�w9��X�����;Us����^p��E�-o*���V�#��m��Ha2�d�������
{H��7����;�G���ƣ�Ϻp�1$6KvQYΥոۓ�m�]��s�k�rʖ��z��<N��9��TV�7��=����BxwdBA�+Ѱ��	y����c�	U�H�A3,�]ع8D�{5&�0����M򧕶H޵I+�LK�n/��|K����hZO<֔P�}� I8��S���G��;���B�Z8�J���?{B��"'���c���c#�1��5:P�e�><��EE��2H�T�H ���TDƃ"D���5��E��#1�1֪������D^�߅�Y鷜L!�œ�6�ic���~�y�[�j����a$��-g���0y�\���ڐ��S;c_/Wb�����8�Kd#���On�B.�|�y��Z�ñ�Hb,�GV����}�С3�:�ʒ�Bm��?���ה��H6$�{v%no�� ��S��'��_}xu,􅒬�kNZs�9g��j�x�d(���h���2�|Œg�,|W���a>��P/|�e�!��,M��J�Y�G4ˇ$�4�<��y����9&����c߻��~����4������	G�J���N�#�D�ޭ̞⡠.˲2�b�_�ѻLP��y�̬[���*�t<��B;j��	Ǐ-�N8�=>>��q���������(��UY�g?0-�)������u�ܹs��+��?��O���e��}(��� �N&C���t�w�
a������<{��
�:IQᘁ��(hff��~��~����WdYh������}�B'I�F�j<��������{�5y���n����]�nBX��p��W��X{��{��]"��A)��ϐṛ�Qm�����&#2 ����}�{�?������=�Ȋ}]r�w$������ٚ%	�3�1�|ٽ{�}7�|�o~�c�����}��aah�`1���2	�ߥ�_����'Z ��N�o�zʖS~���O_���裏�ڛ�1�n�H�ڙ��s`�E
����!��3O�{�-�|ta�3?��B�Ⱦ}�@��P��.}��9�L�:��~�w������2.������004B0�={� B�;��-�G�"��+	����c��Ϯ{b��E_������<��K��f��St�d9"'}��z����=���h���_�����{l���G}|s�y�����y��
���~�9����!�e˖Z� ��8�(�}���F�Ee�ȪDk�%N� ��/X�@i��9������L����W\q���p�Ї̧>����A̟��������0_Ѱԫ=�3̍7�h^�򗛺04B� O?�tQ�� 'V<]��X�CH�)>ع��LP{%���[���=�A��y��Oኝ%��C*)�pH�.��bw���sT��@ĊGaM_#���ج*��y9ؖ,�h@�!�V莩�'���ֲ�{�@#��L�H�+.T��zwh�p�G�椔y��$�U9<W;'dڛ��m��"܀��)O�M@Sg0�d��7�9�؈���8�(۵z��c8@D���Er�|֮ m0��k$)�'�:*��D�@�sD�s���F���0�}ᱦ�N�;+"��A#��~
y*�*�B��A�T5E0��>:Պ��l;*�*C~�^�T��Y��8[��a�����g���4_\l�z[�eAck%-�ك�2��f ��:)9,C��,�	�!�+��_�:��B� �H�;��Tg�a׭[W�p �ICA�l^R���l�Ӈwt\�.4β4H�8 �o��@�]"�AA�E���ڵˮ�P��t8WS(Q���B#�j� -d��1!$J��|$vmT�L]F�C��m۶�:�"��P}�L��\���:E
44Ʋt>���(
�`l�h
�Q��}u9����:QE��5��%	eF\��4Ͱ�`:e��$���h8�^K�*6 �����_u��u�3i-K�$rQ
X✊d86͜l�U���������e����q����k�F���}Q�9��ؚ�F�R�8��9���hDC�T�kRNrw�uhʣŲp46�@�}y|G�?�w���TE9�bJ�dW1؊*��2��e.��ւ ���+�O�_�x}ѯ�St=C�	h�p@_�Ž0	��J\�V���cۢ]�@C_�V-����&~$��.�\%�8�t���~���a�)$�9��*� r����3B�*]0By��iyҟ�l�&�1
�?Q=:o�T�\'\�*D����Q>�k%�Uwj��	r���@�ŸFK�5Y!L'G���r���:�^� ���Q�E쫖��c/�# D�A!#ǲ�r���T<�:ÃE��a�����h�N\'L-vrj�ԡF?f.�Yf�hW�[�X�~G���wPf����g]��lظ�V�X1eqt�m��j����b}M���5���f\'i����,>�N�Q�W��,�N|�Wϲ��=x�`l7�p�GqV�]S�
m.+5N��h�g��F"Ņ:�*����Q�zb�9Ίf�.V�����;�<�v��a�
e�s�vb�"!0r�����wV� �l�$<8Yx�X����*�P�^�l�Ey�9��lAu��x��P��J����E-A�1	9v+�l���X� ����\V�C�p�-����_И���A�U�VEә���u�¬,��K�<$�p��J�5]hEE�{k* U��X�Q[�W,��j�3�{Fee���@Fr"RC�A#͚D^�,F ���ǌ�P�Iq�X�Y�Z.Qqg������J>�L_0��h�O�1 �a���$�x ������յ�M(���d�P��H^�W<_�B�E6w!�� �Q$�����¶$�@�n�(���R	�%�#�C!��d���P`9�^�D��$9$�����)jb)`Uۿd�*k�"+�O<{�+_����۷���NJ?��+l4���BM@�jo!�Y���������Z��
�Q�Ca�2�4QH�`�j�S��HºM@#��f&l�WV���C�Â�YL]'u��C����$��r}(�ܒ�:r�M!���Oh���Ak?�H�(W+#]��d1
��xM�ãl''&�����X�L��%�&Z��c1$*�4���;Eb!:��Y���(-*K��1� $��[��ƭ�,+3F!/�R�v�@�����!����d�_�r��.P
J:ɱ�a����ζDC��be��	|td*[+�2
E�6�d:��@ �+|�1�1�a��4��$��
HA3����;#�('�z�L�!�n�b�E�-�rbb�u-�D��Ј�l���s��ִh,R�!�w�&1��^ˀǢ�ǆg��i*�6�Ȏ;6�ݰ ͑�\&�E��u�S7!
i���4�:��b��z�B�8Bo��ٱ���?uB	е��ݑ�����ϓ0?CB�B��ȹ�Yf��ڶ>��)���GNPqe��kP�!�����TQp��sU�:Иګ�D�����"�4�P?����w�7���wNG��k��_�e��t�둰�&�ɼ�B��v�����P��.:.��~��݉��]�v��C,E��>���6r���`��,?�sr���z�c9\+H����7���0LOO'��H�=MTl���:d��#n��Գ�"l196Gy�@İ�	"�T�?�a�G�-\���P<<&7rY'�����U� x�r�E�����S��d��"�����R�=���"נ�׉�kh��ve9����ϫ���F��h%� �ZGЪqfrQر>�b��{�T6�'�Z
^X���������jwZ�6@4:I9�{>D�Y>],2D�E���:F���j���kZ����t�+[W�����N?�������C�TB�mk���`��(��O�&��IB��z�>�e-�T�z{��E;4C���N4DL�)O-N��9�y@���H�g*kB��".�T!p��޽mg�Ag�K��|���u4�����٘��I�Ȩt�4�ۛI\4@-g����xV==�u��if3���d��\M����H(�)E����Ն�B��M;�N��� `d�=z����E����;�ա����iO�1T�:e<44)��QGx��} �Lq�RĚ�F�d��H�I�Ixf��"M@�'� ��K
	Pa��p�9���y� �*X�ZP�V�hY�����5Rv����M��`��D�jaY����֭�G����
%�4'7rǢy��V����-RT7�U�p�"���Y	�S)L��U��哭G�.C�����Cu)��(�U�!��Q���SO=X��Bf*�KVv�X�F*H�Z�,��YOM�	?n
���Bi Ȫ;vt�D�:m�[Q����=�H���6M��r²td���M��]���,,�:j�r�ds�z\�(X��9��;��@����ES�+���0J���Nv��yJ�G��C�f b(i�M@��� \ĥ��ۺh��( Y$x{��&*�`*�I�^DN�TL�8��'��klں�]v� �
�u�od�4d����i��h�T{���*$+Eg���/�j��ȣ�D��R�*1d٫�ÒȨ
M���U��y/-��uu�/T�সe`+��+X�M�6ن�;�b�"�$�"B]��64��N;t�L1���k��e7��^�ʁ0[7���K�ֲp$�NxQ�IHyڍ7�&X���U]n?��>P"��sQ�!�G(��ݮ(}�d����k��-�1|>id�kY�A�ʼ(��~W'F!�y�)P�J�<R���Oʴ,yR�|������e�!@H�a"�ƨ�)'Qh�E���v)�7RB]�l��Le�

��ք��x�N���Nl��ګ
$B��"髬�ۑs.jo/@�d�.�$}IF�,�$��'1 ���a#�TV\<�7�2G�BJ>�,^��W|��U��B�c�{+s$��Z�B�����O�*� �l?xp)n��6H�r1 tN�X��l����AV*��n=̫;��ȑeUs���C��AR#^^>��aYB�N����ԡO'j~�X���5B��!(�_;bȆa*�3@W� �p$�ԮJ���N� g�����Յ&-��>�)���
��(�!�i:z'��!�.���z�h���x�+����:�f�ԕ�(z�f.
h�!���1���sN\'�+���4���<�,Ͻ��������F*�p`ϧmH�eqnݞ��PEk�=�R�d��;:�6�,��,��mD������/s�+�&PvB;��PV+ǫ�j+'�Xv�F2�N[�y�����$���"<F�=[�B�:�K�O�҂81��ix�^�6��EO�\2�FeҌQ�$��4��>NWb��\ �/�����=,p;���OcW�����_�<�=��]G嶠<|�^?��eC��g36j���"I)#��k"b(ڔD#����j7�i��VK��A6�������� � ���+�@�L��@��c���ѫ'`�p!#'2bp!#'2bp!#'2bp!#'2bp!#'2bp!#'2bp!#�}�zW%`    IEND�B`�PK 
     $s�[����E �E                  cirkitFile.jsonPK 
     $s�[                        �E jsons/PK 
     $s�[����H  �H               F jsons/user_defined.jsonPK 
     $s�[                        ڎ images/PK 
     $s�[�R�W�  W�  /             �� images/e30496d1-6e1c-40fa-a66f-2add70ecdc94.pngPK 
     $s�[$7h�!  �!  /             �9 images/a7fde0f7-2836-4f0c-aad0-66dcccec46ff.pngPK 
     $s�[��n GV GV /             �[ images/5a738b76-89aa-4728-b8e5-f09c859dbb14.pngPK 
     $s�[����C   C   /             u� images/ba153158-cccd-4fb1-9320-38bebad1b7f9.pngPK 
     $s�[Y�u�= �= /             � images/fd2cb464-8539-444d-bb0b-3750bec3ea07.pngPK 
     $s�[�z��gW  gW  /             
 images/3024baee-4b71-48cf-83e2-7da05d24f50a.pngPK 
     $s�[�ة� � /             �h images/8f771a2d-db90-4bfd-8b3e-8d66edcda07a.pngPK 
     $s�[��/F��  ��  /             �� images/0c7fd013-2f4e-47d0-a46e-2d19cc1fd6f6.pngPK 
     $s�[���� � /             �r images/bf314729-9196-4b76-b154-4ab11fec66f9.pngPK 
     $s�[Q��0�U  �U  /             �� images/a88da2ca-7e0d-495e-a5bf-cdc1eeca5e78.pngPK 
     $s�[�����  �  /             �� images/879f6d20-9391-47d7-8a0d-9140b0e14aa9.pngPK 
     $s�[�^�}    /             S� images/c5725ab6-c6f4-4984-98e2-b9c0e10adf5a.pngPK 
     $s�[y&��:  �:  /             �� images/4a8a1475-7a47-485c-913d-9939fe0b1f0f.pngPK 
     $s�[�Sd�%  �%  /             �� images/3357ace3-f4e2-44e5-8366-d3a4568261a9.pngPK 
     $s�[9&��ސ ސ /             � images/b01488b3-8551-4b4c-b09f-2812c4acc168.pngPK 
     $s�[d��   �   /             � images/d3b73945-fe79-451b-b309-b64aab767520.pngPK 
     $s�[��RL  RL  /             �� images/f093df24-6efd-4d47-a863-17c5645b3aaa.pngPK 
     $s�[2)h�V
  V
  /             � images/72f663bc-d85e-4d27-9085-2f4219a623d3.pngPK 
     $s�[
�8b  8b  /             9 images/a7e3301e-fb46-458d-916f-a05c0bde95f4.pngPK 
     $s�['�Y��  �  /             �t images/4bf63cb1-3675-4452-8ab6-1403298522d5.pngPK 
     $s�[Vm�80 80 /             �x images/9ce856c6-be81-4769-87b3-53be9928d02a.pngPK 
     $s�[��C�I  I  /             V� images/627fe4d2-0152-4b97-938d-4b9176d7a483.pngPK 
     $s�[�c��f  �f  /             �� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     $s�[��EM  M  /             * images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK 
     $s�[y�E�wf  wf  /             �= images/6a97e33c-aa93-4e7b-a2bd-349ce97096b8.pngPK 
     $s�[Ɛ�~<  <  /             x� images/e65d6d59-bd1f-4659-a32c-fe6c1b0070ef.pngPK      ]
  ��   