PK
     o_�[Z���0b  0b     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_0":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_1":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_2":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_3":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_4":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_5":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_6":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_7":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_8":["pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_0"],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_9":["pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_1"],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_10":["pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_2"],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_11":["pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_3"],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_12":["pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_5"],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_13":["pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_6"],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_14":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_15":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_16":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_17":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_18":["pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_7"],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_19":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_20":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_21":["pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_4"],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_22":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_23":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_24":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_25":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_26":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_27":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_28":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_29":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_30":[],"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_31":[],"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_0":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_8"],"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_1":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_9"],"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_2":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_10"],"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_3":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_11"],"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_4":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_21"],"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_5":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_12"],"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_6":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_13"],"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_7":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_18"]},"pin_to_color":{"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_0":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_1":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_2":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_3":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_4":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_5":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_6":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_7":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_8":"#00c7fc","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_9":"#9E008E","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_10":"#0E4CA1","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_11":"#FFE502","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_12":"#ff8647","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_13":"#77bb41","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_14":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_15":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_16":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_17":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_18":"#e32400","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_19":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_20":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_21":"#005F39","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_22":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_23":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_24":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_25":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_26":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_27":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_28":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_29":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_30":"#000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_31":"#000000","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_0":"#00c7fc","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_1":"#9E008E","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_2":"#0E4CA1","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_3":"#FFE502","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_4":"#005F39","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_5":"#ff8647","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_6":"#77bb41","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_7":"#e32400"},"pin_to_state":{"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_0":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_1":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_2":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_3":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_4":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_5":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_6":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_7":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_8":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_9":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_10":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_11":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_12":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_13":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_14":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_15":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_16":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_17":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_18":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_19":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_20":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_21":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_22":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_23":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_24":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_25":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_26":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_27":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_28":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_29":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_30":"neutral","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_31":"neutral","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_0":"neutral","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_1":"neutral","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_2":"neutral","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_3":"neutral","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_4":"neutral","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_5":"neutral","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_6":"neutral","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_7":"neutral"},"next_color_idx":8,"wires_placed_in_order":[["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_8","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_0"],["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_9","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_1"],["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_10","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_2"],["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_11","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_3"],["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_21","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_4"],["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_12","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_5"],["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_13","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_6"],["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_18","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_7"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_8","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_0"]]],[[],[["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_9","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_1"]]],[[],[["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_10","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_2"]]],[[],[["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_11","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_3"]]],[[],[["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_21","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_4"]]],[[],[["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_12","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_5"]]],[[],[["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_13","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_6"]]],[[],[["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_18","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_7"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_0":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_1":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_2":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_3":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_4":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_5":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_6":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_7":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_8":"0000000000000000","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_9":"0000000000000001","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_10":"0000000000000002","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_11":"0000000000000003","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_12":"0000000000000005","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_13":"0000000000000006","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_14":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_15":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_16":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_17":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_18":"0000000000000007","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_19":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_20":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_21":"0000000000000004","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_22":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_23":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_24":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_25":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_26":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_27":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_28":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_29":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_30":"_","pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_31":"_","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_0":"0000000000000000","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_1":"0000000000000001","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_2":"0000000000000002","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_3":"0000000000000003","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_4":"0000000000000004","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_5":"0000000000000005","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_6":"0000000000000006","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_7":"0000000000000007"},"component_id_to_pins":{"3e8f3730-0a34-4180-bbe6-26ef6579f9cc":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"92d25e78-3dd4-4c51-a639-7d3b45229763":["0","1","2","3","4","5","6","7"],"e0fb8dc1-0c99-4975-9f66-ec6cb925550a":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_8","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_0"],"0000000000000001":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_9","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_1"],"0000000000000002":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_10","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_2"],"0000000000000003":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_11","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_3"],"0000000000000004":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_21","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_4"],"0000000000000005":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_12","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_5"],"0000000000000006":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_13","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_6"],"0000000000000007":["pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_18","pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_7"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7"},"all_breadboard_info_list":["cd97cb21-4bc4-45ac-9ff9-5eab3251e3e0_17_2_False_655_340_up"],"breadboard_info_list":[],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[1176.25,432.5],"typeId":"23db5403-7550-740c-a02b-8b3755757442","componentVersion":1,"instanceId":"3e8f3730-0a34-4180-bbe6-26ef6579f9cc","orientation":"up","circleData":[[1157.5,575],[1172.5,575],[1187.5,575],[1202.5,575],[1217.5,575],[1232.5,575],[1247.5,575],[1262.5,575],[1292.5,575],[1307.5,575],[1322.5,575],[1337.5,575],[1352.5,575],[1367.5,575],[1103.5,290],[1118.5,290],[1133.5,290],[1148.5,290],[1163.5,290],[1178.5,290],[1193.5,290],[1208.5,290],[1223.5,290],[1238.5,290],[1262.5,290],[1277.5,290],[1292.5,290],[1307.5,290],[1322.5,290],[1337.5,290],[1352.5,290],[1367.5,290]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"db44127c-0abc-4a16-a9e4-8c8b90de2dab\",\"explorerHtmlId\":\"d0aa30eb-e06c-41f2-bb61-1cf6ff30febd\",\"nameHtmlId\":\"9003496d-cb51-4255-844b-61003da77163\",\"nameInputHtmlId\":\"dc8b2013-6f50-451e-bdf4-b51be526a925\",\"explorerChildHtmlId\":\"a8a687ab-5e10-4f91-8eaa-1c099947f137\",\"explorerCarrotOpenHtmlId\":\"cccd7f49-8ed7-4e7e-aa56-792cfb9e03e8\",\"explorerCarrotClosedHtmlId\":\"149f2432-66ca-445c-aa9e-4182d8e33496\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"8c466249-d84d-4671-b907-1997e2891945\",\"explorerHtmlId\":\"323f230a-1faa-4490-ae94-2465bef782ac\",\"nameHtmlId\":\"8e8d751c-fd5e-4ea8-b699-f37466e2f89f\",\"nameInputHtmlId\":\"12fb3675-ff4e-48dd-832d-1cce4135ac92\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"78b5a5a6-432a-4ab3-9460-cb9a20f66e76\",\"explorerHtmlId\":\"27b9225c-7312-4f16-b407-c174e73bfa8a\",\"nameHtmlId\":\"5026ca79-3035-4380-b20b-fa3b147f773d\",\"nameInputHtmlId\":\"1d47f92c-87be-47f9-8e3e-19e65b778388\",\"code\":\"\"},0,","codeLabelPosition":[1176.25,275],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1621.672258,295.18009100000006],"typeId":"4898f56e-60f9-4315-8c2e-83ff52744e63","componentVersion":1,"instanceId":"92d25e78-3dd4-4c51-a639-7d3b45229763","orientation":"up","circleData":[[1577.5,515],[1589.021389,515.1630365000001],[1601.4649255,515.1630365000001],[1614.1045,514.9239635],[1626.7010365,515.5090730000001],[1638.4094635000001,515.5090730000001],[1650.5069635,515.6160365000001],[1662.5697220000002,515.5428290000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"4×4 Keypad:\n  - Row 1 → A0\n  - Row 2 → A1\n  - Row 3 → A2\n  - Row 4 → A3\n  - Column 1 → Pin 10\n  - Column 2 → A4\n  - Column 3 → A5\n  - Column 4 → Pin 13","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1056.6005859375,156],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"e0fb8dc1-0c99-4975-9f66-ec6cb925550a","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"57.27872","left":"945.00000","width":"815.72483","height":"542.72128","x":"945.00000","y":"57.27872"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#00c7fc\",\"startPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_8\",\"endPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_0\",\"rawStartPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_8\",\"rawEndPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1292.5000000000_575.0000000000\\\",\\\"1292.5000000000_680.0000000000\\\",\\\"1577.5000000000_680.0000000000\\\",\\\"1577.5000000000_515.0000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_9\",\"endPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_1\",\"rawStartPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_9\",\"rawEndPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1307.5000000000_575.0000000000\\\",\\\"1307.5000000000_665.0000000000\\\",\\\"1589.0213890000_665.0000000000\\\",\\\"1589.0213890000_515.1630365000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_10\",\"endPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_2\",\"rawStartPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_10\",\"rawEndPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1322.5000000000_575.0000000000\\\",\\\"1322.5000000000_650.0000000000\\\",\\\"1601.4649255000_650.0000000000\\\",\\\"1601.4649255000_515.1630365000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_11\",\"endPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_3\",\"rawStartPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_11\",\"rawEndPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1337.5000000000_575.0000000000\\\",\\\"1337.5000000000_635.0000000000\\\",\\\"1614.1045000000_635.0000000000\\\",\\\"1614.1045000000_514.9239635000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_21\",\"endPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_4\",\"rawStartPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_21\",\"rawEndPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1208.5000000000_290.0000000000\\\",\\\"1208.5000000000_57.5000000000\\\",\\\"1757.5000000000_57.5000000000\\\",\\\"1757.5000000000_545.0000000000\\\",\\\"1626.7010365000_545.0000000000\\\",\\\"1626.7010365000_515.5090730000\\\"]}\"}","{\"color\":\"#ff8647\",\"startPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_12\",\"endPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_5\",\"rawStartPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_12\",\"rawEndPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1352.5000000000_575.0000000000\\\",\\\"1352.5000000000_620.0000000000\\\",\\\"1638.4094635000_620.0000000000\\\",\\\"1638.4094635000_515.5090730000\\\"]}\"}","{\"color\":\"#77bb41\",\"startPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_13\",\"endPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_6\",\"rawStartPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_13\",\"rawEndPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1367.5000000000_575.0000000000\\\",\\\"1367.5000000000_605.0000000000\\\",\\\"1650.5069635000_605.0000000000\\\",\\\"1650.5069635000_515.6160365000\\\"]}\"}","{\"color\":\"#e32400\",\"startPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_18\",\"endPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_7\",\"rawStartPinId\":\"pin-type-component_3e8f3730-0a34-4180-bbe6-26ef6579f9cc_18\",\"rawEndPinId\":\"pin-type-component_92d25e78-3dd4-4c51-a639-7d3b45229763_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1163.5000000000_290.0000000000\\\",\\\"1163.5000000000_35.0000000000\\\",\\\"1780.0000000000_35.0000000000\\\",\\\"1780.0000000000_560.0000000000\\\",\\\"1662.5697220000_560.0000000000\\\",\\\"1662.5697220000_515.5428290000\\\"]}\"}"],"projectDescription":""}PK
     o_�[               jsons/PK
     o_�[rfƣ�  �     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino UNO","category":["Microcontroller"],"userDefined":false,"id":"23db5403-7550-740c-a02b-8b3755757442","subtypeDescription":"","subtypePic":"0b351edc-7875-4477-b820-546ce15be531.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"4x4 Keypad","category":["User Defined"],"id":"4898f56e-60f9-4315-8c2e-83ff52744e63","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"bf314729-9196-4b76-b154-4ab11fec66f9.png","iconPic":"a88da2ca-7e0d-495e-a5bf-cdc1eeca5e78.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"17.20701","numDisplayRows":"30.38685","pins":[{"uniquePinIdString":"0","positionMil":"565.86878,53.87644","isAnchorPin":true,"label":"R0"},{"uniquePinIdString":"1","positionMil":"642.67804,52.78953","isAnchorPin":false,"label":"R1"},{"uniquePinIdString":"2","positionMil":"725.63495,52.78953","isAnchorPin":false,"label":"R2"},{"uniquePinIdString":"3","positionMil":"809.89878,54.38335","isAnchorPin":false,"label":"R3"},{"uniquePinIdString":"4","positionMil":"893.87569,50.48262","isAnchorPin":false,"label":"C0"},{"uniquePinIdString":"5","positionMil":"971.93187,50.48262","isAnchorPin":false,"label":"C1"},{"uniquePinIdString":"6","positionMil":"1052.58187,49.76953","isAnchorPin":false,"label":"C2"},{"uniquePinIdString":"7","positionMil":"1133.00026,50.25758","isAnchorPin":false,"label":"C3"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     o_�[               images/PK
     o_�[P��/ǽ  ǽ  /   images/0b351edc-7875-4477-b820-546ce15be531.png�PNG

   IHDR  u  v   ��:   sBIT|d�    IDATx���}tSwz/��$۲0���Mblc0fB��3���@��0�b�!d�qN�bν'�tAgڣ�rf��i��Ճ���M�8�Ms�z��� N�`L�~��-�/��ClE�e[/{k���Y+kY��O��g?���S��ҡ�D�P�C���{HDDDDD�;����_��{�R�=�p����V)v9""""��Ή�:�t(I�R�)xZ�Q��5�cR�GBנP�@��x�1�cR��+o6I���t�|�&�I ����W��ǙM~��<>/(�^h�J""""
O����=�p���`T��F��:ix./M�8�IV�0<<,�0������ ~�}�M�Kb�J�/^:���Q��)��ӣ ]��+���!�L-[�,(q��~cP�Qx��+u>HT�*�GT�K�N�F#�0�����BN�T���@{��c�NQ9*���!�S�=�p�n�DDDDD��abg�{�aR祄W��="""""�G('v�~I�v|b��
[�M�6ן)�B�;JX�&"""�^�N�dRDO�f੅�`�b���y��A�����DF=T*~��"�bb�������_��g}� �L|v;>��f�@�|y`��6��~�PN�JU�Pث�B�GIDDD^B1��^Jx�PI�g9������~�1��y��\oo/���@�Z����80w��Y���G'Q�f
���c��	��0����'�C
���䎈��h�P�:�aLv��0�Ə��8��/�ҡ:m�Ҡ ^��٨���w��cqyX˸�˸�Ըb����q7��
B�b�J��X���Z���qu\e����MRʕP��{`<�}���R�a��A�<�,]�q��G��s"�������m>=?*v�~I��v\���H�����_�W�J�@�g�DDDDA
]1���1!����(F~�r;"""���N���);`W�*���	F~�r���`�#"""

�r�f��0e�tk�f����봯��f �S&&�ݮC�RA�R1.�2.�W,6����O�P ֋�y�q7��I��f��b�`xx `�Za��  � ��������"��<x��:�����e�?�S `||f�FGGKllRSS��!�2.�2��q�b��1:j���H��R*��?���\�e\�<n8`RG����`�Zq���ޅ��?�6�������9Z-���/��#�uB�)�o�<`�P�B�|ǟ_W*�P��D h��q�?>�v�Wg�˸�˸���B��J�9s�tA*\����xu1ʸ�˸��L���������z��c;Vcn������ݻ���|���>�����ݻHNLD�R	����	L���X`������͎/&&�y��]�����BZf&������(�k�Z���?}(��"<����8f}��6��1���F�oV�[���pa�P(`���q�q%�+�@.H]/D�q7�qCYd���fý{���ڊ�`�Ղ�y�H���%&c�}p���� ��#QJE,���0������F���`Q����b����ܩ����)lF��� 7&����q�q7Xq������˸��	���&A[k+�:��א9/��x���`��8J qJ%�J$ƨ`�����������'�=�RRR�z���.�Z��ƕ6c�MPR8.�ZZZ�~�ʕ�D�0c\�e\ƕ�J����;ר�fɒ<Q.D�q72ӟ�|U��Ʉ/._��cu��j��Q����qc
̍�A�J��]��f5z�菡/-EFF�#�"v4�=W#�x�I�ꛦ@�`
�����&�)�e\�e\�X,V�_���~�q7��"��d��_��G���I0wv`��W�1
t11xT���}�O���B{{��1"�ݎ�oa0�K4������:��d�o��a�ڄ�9��&��$�� �T���x�_���＃��nIbE"��� �&�D����(�0��r###�M}=p���`W�A(M�*H���D�u4��?��ݻ��$""""�DLꢘ�f���1|�7��SWWP�����k���gQ6��t��W��!Q4aR��Z[��#;I�� 't�X�ɱ1�{���ٳA������(0��R###�ZW�m"�;�2�r:j��qq���Z���m� !�r�a2�MY"��������(����B�sc����e��F��vxW~�kV눈���|��.
Y,�7��|�C==r�c�����~�vÜV(V��ЫE&uQ���Z�#���N��,N�D�݆�S��J�
�J���@DDD�b�@4��ݥؖ�,�Y��5O�C��`���54`�ܹ�Z���
�����s����{H�'��9?>T��A'Ʊ��ӽ~nll�!�q�qe������u			�˸�BqC�� �L����z����_H�X,�tu ���m0�X��!t~�%��^QJn
@7��C�^�N� @�MY!�q��Ұx�b�~gxxV��7H�q�qŌ+�����;V���Ì˸�+s�P��Q���/��T���/�P<�Q*�Q����,�PB��.N"%��@������D�/!!j��q�q7hqŒ��������{j�:�J�2.�7T1��2��혫���phn���cm]��~'�PB�B�����=��WU(��K/��^�1.�2.����Q����˸�x�P��Qftp�PȾ��LT
��^ht�Uj��h����^:��P(���u�J����.�			���^Mkf\�e\��5�X
E��!)�f*)�2.�70��2C�3�'�J���.���(xZεu��!�*]LLFGG���+�x�v;�2.�2�$qŢT*#���q�\1��211*����ƬT
�G��P���P��/^n
fܹ�*W /r�͆��Q��ĸ�˸���v�,�g\�e���5uDaJ�b&�F�t()X1���P�Jc�����E�ؘ�(�*Y��B��J���nΏ�ؔ�6G!""""q1�#
sBb7�Ǉ$��oʙ����(ېh��j4rcF���,��B�@A�Mِ��������])�x�P�æ(~�����w2�����:�<�������a1.�2.�J�A�<|�rیω���q7��"^9{)��C%1P�	��K��?��Ǽn����+z�իG��~��|y��	Q�-���	Ld/Ď��I����%9n����Ʉ�f~��@���ʡ
�BiP EQD3���,�+uQF����/>Gl|<F����G�v;�͐{aK���1P�Ѿ��'v،C�Û/x���ĩT�
����Qx`Re2�z|u�#h�ڐL���vL���Z�B=�O+�|Z�w쯼��ݎ(lm6�\����

{�(Q(P L�%"""����.�:�ڝ^<��>�R?O��&��		S�#Y����;�?P�v;,6;�=���P�i�Oʩݑ�8N��Z�>��  �ͷq����#"""�hƤ.����M��ۛ^=�؎՘+�ǳ`u�?�-�B�Z7f�#5�		r�h���4��� �Ä �m\���.�2��,��`�Z�����Iu46m�5�������CDD���A�{�i�3����*�P܌���۠��?�{(DS�4jԾ��-��.@��2��I5�v�PV���t�ㅙ�0���/+�'""���J]R'$ ��߃��fHU�6�s�h�j��B4E�~1����� ��q ���#;E���AY�竺=ې�Q��ݏQw���gBbW�gJ�����$�()�%i�����ꛤQ���#�����U4��`	�����I]�Z�y3>�������H�6F�6<U�W�y����6��Q�� P�w�3�[�� �a�ԕ�03�oECKǔ�7u����h����X��3Wd%��$�U��P���V�0[��kB��IΧ$�Ez$͉��B3�zM0�;Ө��ك�O���G�؁�Y}�rпk9�:6?�f4�t�� �9% Z:`�o�}��1���P����(�#'U��7�a8�i�n(5T� �T������R�π�]����Iա��է/OIn�vJ���Caf:*��(�L��A��I]�R'$������e$��b�����2a��j�!q�rV�$�؍ӈ��t�Q�|��4�q��}�^??ntK��J[`�1��[U;a�o��TI�03M�=��.�"�@W�F� �]��8V,q\��t�$/��b�����9�Iա�j�󮼐 U�_���-h�Daf:��lsܬ��.I�FyAJ�fKrq�� ��B3J�`ܽ	m�&�w�|��+�B�!$��bT�_����]��$�%yYh�ډE;O�d���1�p�ؚ<��_��B�]Q���B���)�����s~�m�&g���HҨQ��.˿CR�(ңzG)�zMh���o���AR%�rbR����p��e��Q��`�b�� ,6�J��/�"�����'��^�Ռ��x�I|��Ը��� ��+nt�>���:���˜�i��P�w����[��:��iҜx���L�<�ԫ��:	��s�*]����b�P߈���h�쁡����0�����fA����8Ū�+U�IS���ls\ؾ��(q�V���0l~ʭr"er'�o%�G0`�¸{�:{�>��ӗ/m~J��M8\+w�k~�><-J�$�U�W�����g����U��r$�6!�5�7:���F��)��5l~����`��*�^�S��*�����2�Z���|�#�%��(�����?�	]����ڂ�ؙ'&`��P��͎�+����^%vb��&�3�s����Gб�ȹ��5����h=�t�^��4���gO�	�J��=DI^�ǋ�����VSg���\����k�����f���:{P��%JL)�XP��Ǩh�pT�&�-h��ASg���sRu��v�y��1����vK��-I�vN��:��B3�o�qU�v�#BE�����b)��r;?��\q|��r{�����Ϸ���oEݞm0��$i����9��k
ڍ:�����^�O��o-��(�NH��?z	��7�@F��:����Yl6Xl6<��z}PbF#�+�l��TqgJ�H��wocw�_���6�fck*��=f��4���#p�J'֜T�E}��V���rR�n���z��
����sKĎ+�f/4;�r����V �zMn�[CKrR�S�����dm[E��9�q��b^��A��M0���V-��b��n������3��{1�}0[Q��ǎX{�IV}5�7b`Ă��U(������0[��TeMҨk7E�Ć&u�y�����������I_��yX���{�R��g���J��%vR����I��	�_b�K?F~َ��|���:bO���iHr�<����6���]mA��RwoBCK�V��X��<����C��R��e�����ݛд�nu�;J��ԕ�WjBr��Q�di�#����B3��ls�w���>V�_�;'ޙX�y�?0b�m�p�w0[a�Ќ�T�֯���j�5���0��PV�ܣS*7�a(+F�ي�3W��h)/�s~O�|�B\C� n�;oX	�_��I����Q	��N&�$�I�:*ۓ�/���(_����Hä� 8���j���~�0��+I�q��	&�
<��V�$$ub%���+�kb���5���Q/A�`�xu�t�l5ቶiH�;J���O�i��tęr���	�/��W����3WP^���-�><-�U��T �)�U�v$)��-q0�7��܀�*��.W-�u|�;���*li"�6�7����/4;�f��%VBYx��VT}x�ys	�d7w��\AҜx�t�����K�r�|��g�8���,�ñ�I���ZQ��<�B(܌��j'>����r \$�z�$�3��wl�j̍~�mƥ�%l-7��h���=Q�����0n�#&�Q���	�����{�3u%�=v�44#��[̔�(�FG���#K��ێ�1K��v/X���&i�h{mϔ��+�d��<%u{�9�	�֯Dݵ[nI�q�&$͉w�o�".�m���ׄ�w?F���:���H�`�-�3���>(���C��{��J�4'^�q�$'U7�1�	[P��3j��A����_�
	^�>/�r/l{!��TF,S���3.0��Y�~%��e=�� |�#4u��|6���,�+u�F���5�{��܌k�|Z�s���N�d�f�æV���ǲ?�C�Nn�>���1Y�&<�J��S\MW�4�����d`�"ZBmӐ�F0u{�9���0��n�6g�W9)Z�,�FI^�dӢB�1n����dO8Z:B�
�{������ӽ.�_�lǏ��P����*ؘԑGz=2~�:���q���	�qq�%%�n�atx��a�'<_H��혰�a�c:[|<����d�ȅ�{�T�gm�-���<�8����g�8�)��t��>ga�]�$_DDN����/����S��e�����`�b��4�S������9|s�"�{�C��F������v�Y,Ǹ��ݎ���1O��%6bޢEr�I�R����bb�������_��g}�߿/P+��C51Ԙ�΃�l���-�Y���ʊ�����$R�]7[�Nh�`Jw8��G�4$O�w0M6\�1���(Zp�exj�#���{cc�]|����LR������ہ�۝�u7O�뜺hQH�7�]˳�����s������ΰL�����q�g��{}&��[�M�x	ӳ�O��ݙ�����~��;�q=6�u]�S^���M������R�]7ݴ�$�ڹg��Y�S��q�X��|%U����g��d��w#�N�F~Fηv-f��'��z)��ԑ�ع2��$�Ŝ9j|��9ѹ�g��3l6qo8���0G��Wmw<�������fO��!n�(/ȃa�S���"6��tp�:�.@s�}��|+�!/?#�+� ���j/ݐ<f��'��z)���E����P�Th���x��=��B9?]U����F��U��u�~q��2�&���q��Ձ��w]!6/_��Wc߱��� q]ﾇ���b�'p���o�-y�q��E<��2<�jYT�'�ߋ�[ס��)��kr3 &�U�}]�3�P�w;��q3>��ɋ8x�d㐋R����j��s�O����R�".���_$�E%yYh���l�!eB8����$��q���|k'v�s��B�B��lE͹&�w� ���ηv:�h8O\���Z�G�6����gp���{�9g�'o:aL���:"�($T�=ڂ��J���|�ś�w�I|k���E�yM�7?#mJU�sּQ+I���ϭZ6��-���Lꈈ�����FU�WN��^�y�h�ϸ�$u{� ���,Gv�Źp�s�^
��q-�I4}/jvn��XVr�dSm���2}�պH��ʤ��H&����=�$�;0b	�F�MXrRuAm�ϸ���������}?**�b�êJ���-�[�,jΓh�^�۸��y���Bo�-z����A��8�uݴ�9��m�7��7T0�#�r�� !�}Ͼ�ix0<����q A��i2{�Ed\Wf�Ǥj��DW��+�����\�578��uT#��L���;�F��V-CG�P�.z��<����i��dRMì9ׄ-�\�.��A�h�V� &uDQ����T*��
T*�����װXş��so��I��TJ�`�"\��+H1�]����T	N �����T�����ͷe	y���,xU�h;O���z�v9���0+?8���2��ȩ��F�I]��Y>���Gg��y�wa�\uF]������סP��P�����4�Q��~�l�	���i��$g>z�� ��>���mbv�j�������Nː+n�JҨQ��9�:�TA�F��Mn�ih�@��Ge!�3��q��ͬ���nv�:�:(��z�D��n��d��|\����4�H�v)`RDm�Ch���;��G֜�ٟH>��l�|g@�a����<����<���;���6H Q    IDAT,$͉��}2I����-�v�LҨQ�g�c��ӗ�~f�oD[� rR�Ά*rOդ�s�l6/_��Ϡ��e5�=$����{hl������k{���W�'�v�8y���?�_ock��鏮-��w���Ps�	�cZ��#�:""��`ܽɹI���R��}Թ��� ��O!'U'�vEz����	����J�f�di6�:����N���e�;�1��j>B�>����?(y�h;O�����|4�~t���h����D��:""S��0[QQ�w$y~����(ң��G��K�f��f��0n���t���)z��F�EU$�on�4�h;O���F���PŤ��H���>}�Y6��۳%yY�>sE�΅I���n�lE��+n���"I�F�F͆)�N�bתe0����|#���������o��cDD<L�\\\�^4	�%8���&$Jm.SO�d�03]�ꜧ1L69��9&t��N�:[|?���X�F�,����jl""
&u!*F��J5}�>�(�ʐH�
EP^/Q��>}Y��j*���>�$/K�M�#���N$��ߢ��-ؼ|1��fmz����i��1Q�aR���P��������oJg6��9o|�	��A$�6��@ݵ[�*]��������T�_��<T�����&׺�a��ŲĖ�)ɇI]����\�+}��K]}���F��0�o�Z�aE��^�O_���%yY0^hv&�9)ZG�ˇ���y3�=���  K��L��A�(�tDD�I]���i�_���AsHT���j�JT�_9�c��FѧdV�����AT�a(+v�Y[�	��Fne �5���JN��An� ��\���D�]�����:"� 0[=�U�����-��ڂ�T�s���^��Id��f%��?�ڿ���IQDbRGD$���#^=/'U��i;ö����k�4F��i�(�]�����O��HCVr"���s]E�.���řIQ*/�C��%�f%\���3�  �]�"�u/l�MD��03Ezf�;g�q�zM����K��E��<wo���-0�7�M�2�ބ��[R}��w�֯DE�9��o�s�ٱF��n���S��L&��i{m��}�\5u�x]� 
G����d.'U��^���p�]�Q��w�àe{�9���^���Y{�#��uO@�Q56E'9���"=�w�:f��N9~I^e�(/ȋ��I&u��̕)�f�ø{��lC�ύS�����^�=�۳9)ZN|���P��U;QR}d�4.o�9��۟�^ۃ�^SD~�&�Z���qpL�du.���V�;�	n}�6���֮�%u}����)YbQ��+��(�;�a�a+���,��ن��+#�bǤ.J4u����T�(u|��8�K�P����O�]l
���v::�M��}�$/�Q�+�C�F�'͉w��Ä.��^���K7�.6E9��$�������M�=H�p�Pä.��8Od��<M�l��Aҟ����#�"I5��ls�l9}u�n9+ܳMY&""
Ur%Wf+�Vf��xS4I�v4 ���L�HN� ���p��Q�++FN�M�=0^hs�DQ������>IDDaN���x�U�W"'E����M�f^����K�ύ4L�DyA*����������﹖��VT��1eŨ(� �w����-�>}��<��M��.f딵tD�"��FE��y��Q
CY1�Qؓ+�2�7b`����Փ��-0��4"�8`R��֯D���S��D��QJSg��>�$�U����Q;�U�Q���)���g��0^hFaf:J�]e�VʊQw���QX�3��>s�g� 'U��usĂ�Ξo�"i���1��@��/sRu0�ބ$�zʖ�0[�1�><�ܾ�zG);V�������H�Ҡ�H���+��ك�w?���DD6�M����t�������$��?���+80��p���?,Gݞm+iު۳����LV���l��w?"ѳ�O��ݙυ{��ۯ�7w7Hꮶ��j��
^^����t&uDDv�K�b]3&i�0��03U��x̊"��Y$΂aR烵smXk��ܤ���VǨ#�N[�ɱ��mU�n�;۰{��!̝fBRRt��Q᫶;~�����f�˸20[�w:���7��]1f�U��B�_V�m�%$|Ez4�t����y��I��~�j��Z�q�Q�R���������!��KN��U�(EN����MҨ���P��Q��N����*F���>���	���䬘U���hܷ��ݛ`��r$q�W:�Y�E"&u^���~�slԺD�q����Ά&��#���%�F���Z���	8���T��圮�%��2s�����7w{�S(����|#w�L��4�;�W�zM(�(Z:D�j��yA�T�(��Qw�I���''P�~<ܲ�[�N	d��: """
?rW�\��������C��l&uDDDDDDޒ�b�:�L�V�(u&���� �oq���*fR��Q���h��A�ύ0^hƀي�w?v.Aj�ډ�"�dc�+uDQ���Hиw|�^���C�0.�$�3a C}�ǥ?���)��;J1`�F�>u��E��{C�J9���:(X�	s������&G�l�lE��Gg�� L��ԭ�X�#�R�{�`��ݮ��9K-D�o;��H���df+�O_�r�iܽ	%K��4+/�CE�%yY��ꮶ����.Ԯ�_�~�[�jO\�XW�(����(�c��U;a�oDCK�v:��=����F4u��j�JT���������nݼ���
�I����ԡ;'U���?���᪢H��<Y����b&��+��BҜx��MҨ��Q�/�0�#�R�rL�;U���h���PyA��BN�n�}d�d�P��h��m��9m#����^���i��䡩�Ǒ$�T�0�����6>O���7��{
�M�=HҨQ򰃢�di6�V��e�%u���h�5����L��MN��W,���q�¾�Ez��&��\���i�#T�f��૜T��>��(���sw��E��K��/����dUw�����H�r%(�LwV�\-�B���U���0-�P��hn�R��P��&A4��9�:�䡡�f���"�����)�7&'����4կ� o��#�g����-��܎���&7s�sv=��1�����%i��
�l���&W�;J���s��p͞��>���
�4�H�ހ�:""""��]mA�槜2O*��h�왶�2y/Z	chh�pTU&W�Z��2�q�a���,�v&�B�Vw�e��?�ꐓ�CÉOݎ��ҁ�<f�;�ϭ>s�y��wor����Kv��{�C (�<�j[�p�\�[ ϯz��O��b��Z'���t�i�m�&��ن�=�7$�OnL�"Шz4#�݇e"&V���sS��>�jb,�q������3c��$/u�nI:�
&L��vE�Y��Φ�H��؅����4n��U�
3��p��m�eCKJ�]�Uw��m
f��%�W�������2%U�|1��q8x�"���]O.��Gq��.��e�}��g�CG�Z��x>Ea�\[ߠ�1�.�L���+&uD��e�x��$���ĳ�p;� ��w^�,���EX���Ci�j\""�ʹ�+�C�^O����zf�_�ufBu��f;�֯DyA^@S���{la_�~%�֯t{��j�]�Ȧ�geM�
UɆ�gϵ7YCK��rVq��®���Qs�	 P{�j/����L�]W���;�]���'��|�Y�Z�b�W	��B�䛁W���	���(b}���˪N���A��;/��  ���������5.���K|��t�,y��r6Ez���9s�ʖ7rRuHҨ=&��L��Օ�e�-E����}����n��L7ƺ�-0l~
���0[��2��j��
�d�[;q�uj���}'�㍀`��}m��<�s��E2&uDL�krB����`$vL�HJ9)Zgh�!L1�JI^rRu�H�Mi,�4'~��,ꮶ�03I��4N�6�9���칾�%���.���S �����E8���:��ΔXI��1�#")��9�|�0M�x�ٱmA�S!gC[�	�~����f��$5m������kKա���?{��s����j�w�pt��$����*iN���n�ȑ�y����1a��H�����r !!a,!!!V��^zD?2fW���#���?|D�1�;����7��N�fK褊�Mb%EbǄ���TQ�G���0^h������C}#��7�:3�9m1'U��Ι��~_LO׈E��:��K@M;����w���vT��������E�>e�	d���������P(Rl6[�7�x�b���h4���[
 q
;  �_(�a�4h4J ��Ð���x��i�YG:Ψz�\V����N���n闟�������ݛ���g�J��B�W	S��+h�t44��9���2eSs_�����U.��l��p�d��:]zJRZ:`(+�j�_ݵ[���t
3�e�|���G�
�X[z�+�O���6��^�����INN����Wm�
7�Lꈈ�䒤Q��/+P��Ѩ���E��N�JK�3���,��r%"""��!l�0ymI��������������I:Ez��):peE��{
�f&tQ��:"""""�0�JQ��N�";Y+�0�����z�=�"l�s&uDDQ,?#�{�C'�P�������>�j>���.f��#J�|�0Fu:�l�)���f��A�j_������>cn]��#���hX�#�pm��A[�i����T�sASg�c�Ym�+��(/�s�Z����f��n���z0`����e��'i�0��mJ[w��������&��z�8+uDDU���c߱�rCTLꈢ��x5�t���/��S���0��03�~�|�𸡾�ou>nܽ	�ݛP�QO�e�o��
��Iա��� ��=� 8:�5u� 'U��M��a9J��` ��F�������Z��#"���5uD�rRu��Q���� ��\AҜxT�_��k�����U0^h���U��1�2�Q�~�W퓫�\AyA��P��i��03U�FSg ���C}#��l��A��7���A��ADDD~bRGe�֯D�F��ӗ=�|��I5�4j�z^�Zx��>�o�5�03��騻ڂ$����:�4'ާcE#&uDQ�$/f+Z:<�|�l������-(��Bݞmh��P�,'U���Y��03 �������LꈢLҜx�X|���<����F)��b���&)3%h���z�I��xEz������IDDD��Ѭ�VG�w?vLߜ��Y�~�Ǧ(��bʊ����T�3�ބ�Tݔ�~DDDD��:�(30b	h�����Q^��槜�T\;UΖ�yb(+FyA�����?"""�h'߮�D$��k���Q��77YyA�s����+1�7?r�ss;��/4;��4;�qwoB����x�c�}��hfLꈢL���0[QU����'o.4T)/���|��I��v��S�����?@��l�TaBGDDD�#N�$�2f+�><���{�6��SeŨZ�-Ω�M�=�>sŹ����9Ͳj�JT���EN�ι�x��G9咢Nv���Zd�$�m �67�c�\�e2[q��>���k_A�F���4�g̃N����A|��=9��u��:�(Tw�%�&GW���xSg��'��h�5�� m��q>����H��RYQ�G�F�8��8\�Y���~�(�g��L�ks3�� ����_��`ڟ5�v�\k'�o�z�=��*�F�|���f"+9q��)���i�2��8w��[�"�=��������BZF���'��t�,š�Өa��#��_]����4Ծ�Yɉhl�¾cgq��ޔ�w��d�bד˰c������w���[��6>o�k¾cg �6���uO  j/}�|�u���~��'/N;v�F��[��U���?�'/8��؂����®w��z�=d�hQ��)�O�Z�)X��~#b�J��V�|���������O�?��R�@���_��ɏ��DRQ��Ԕ(��3r !!�k�N�P���~�t7�r�(�}�5j�,r{lB��X�bUP)��o�u|jK+���bhb|O[>~���H��u�(��Κ��k�2���V�w�ηvJCj��\�-�\l^�X��w������5Ed�L���[׹%X�V-Á��ܞ����q����P�q�����p�'/�%э�](�����E�s���7p��E\��
�c<y��oLy|�����}�+�q{|��  ��������_!?c�Ǳ��c���n�����7��s��9��"��o���-n�TG���δ�����
���a��_���]n1�q�o~�L<;�����Y�7G��e���/)f��X�#""�'����p{,sI.�sf��x-!6�w����o&�P�%�ZŐ�6>ϭZ6�z�t5*�b�'$KxYɉxqm!^\[����8|x���ӨQ�s��=��������Q:n�L>W�s`Mn��&;y�X�1m�|k��Ǘdz��c ���X� ��؅�ɳ�G�5��Sn���k���@JB<�-��X,w^*�O��ޫ(Ê�#��>&uDD��AF|U� ������^��B��~��I�t��q��8��i���9�$�8f�d�}�<~v�o,
�ؕ0��d�����p������xs딤�d��d�N���*�k�s���8�ډA˨������?5q9���qJ�[���}�㞎8�E��V�c��}oʴda<��p�鷍�]n�����Z&�6�}J��쭎)cl�?�-��)�g'k����޹�N�tR")��lْ�P(*�@\\�)>>>I����}� �-�r�HU�W�_��?�el���}�G�M�&���%A�Pa|�
�Ō����A��>� �`��c�{�F�W���f�~�v<S����Á:F�?xl!��q�����_�!p$��/�������O��{�!��dMn&�� u�
:���B�~��wܞ�x���"I�ƪ��`�2��?:�������7���Y�����͆�w7���|k6<��F���.�?E��.}������څ�N�gh���X�$�[����;�L����:ׄ�'/:�ҝ�:}׻ﻍ���˨�|�ۿ�8�K���;�S����|�|kηv��>��-:�����_��?���������9�������}/t=C#h�@Y�b(
��@�q���.����Y�P(�34�m_�F�5�*�����q��&H)Z���t�����?����#.��Q��:�dU�W�PV��fﮞH�\gw{,1)���n�����I�Z@��a^�b�'L��;_��2�r�G��	SߤZ&���F�S�5w��HC���g̓%�7��%����۸zʚ2!i���63!�6g����MY;(�ף��5uDDRF'�KY�R��Xb����p��-$ν���ˠP�_��K~F��n�m��/6/_��?y�GN����D$�.��Wv��MGX��ӨQ{�\��ų���n��4�pg2[�$k�SovonŮ'���U� ޻�?+7'""�R�e#!1s��	 �զaђ����t\�R1���8�Ņ~b#�]O.ùW���N����{e�ٹa�'� ;E���
��N �G'u^�Cv���݀��Dh�����B���x�e��[皘 ������>���.��5���m�s���L�$
+uDD䗌��ߊo:�����FO����ڧ���V-s�W�dS����n�͋k����uʪ��[��(��ȹ���}�κ}>�nj��]�ۏPhb�����6���`6[1<t�c#r'(�=��3���O^�8],P�k�^EY�&t�����r��v�R��HCv��c2y<D����<u����'��X�#"��d-�.���u�:t����=$�H��]���e�}��kr8��J񼷗?��q�߻e�?�uk��!�{d2[q�ս5���,L�B�-�    IDAT�Q#?c�3�DM���P_�]Ҫ�������{���P޿|��9�2��^���������?CaSw6�!10�#""�`||f`�L`��M����3f(�\[(j�r���o��ý������5��آ_�2�d�J��N�.�׻��K7P����_�b�G��y�ٹ��9�f�k�2�=՞[�Ǜo#��oI��Wy�*�����\���Jvq�ܺ��s"0�#""�%$$  t:Gu�61�ί?C�|xL�l���mA����8 B���A�^���.}�S�⪣�_���/߀6>{�=�]��T�4��iԨ��.�vR�G��|{������qp�:Iײy�0�g��N�$���4����I�F������jo¼�Q�5)��a���m `��)F�)ڀ�E����ɋ�iWb����ɋ8x�"^\[��W�=�0�Į�bK�	����[��ֹ&<�j�o\�wr���B�k�,�:�b���'l*��1k'u�l���}�7<������{���%v\cG�bRGDDS(Uq��O��wU1j<�Y�{�����;�Q١��nj������lE͹&<yQ�QM�hm����k�:�?�]��nS}e2[q��E�6�Ry��c*��uO���B��X��=�6(�i�صj��sq�������w�\��qn]���f߱����t�cp$%�T,'�^{��hS�3�ܶ��vL3Y�����
g�B\�o��A�(j/}���8���#�pp�:d%'���7�wg?þ���{�*|��%""�hS�C��sal\<2�W  ���a}��v&�h�e��B��������~O!�Ǡe������V�<�����6>5;7x�$Ц(�ͭ�<r
��Q���+��y���[|�lj��pp�:���ܺ���.���oL����in窘�b���~}&�^1�x�mQ*�:�:��	�����	{���O^D͹&����7�:߇5��h|e��gϯzܯs���4 "� ��b�͏<�W����q�����ohԌ���qv��C��6%���KG�Qc�������K7������йjl�7j���Ϙ�ڊ-3>'��1B��yc}P:W��]���;~U�6/��)�a$l�1�����E�L*���+�� �۸�����"d�:��zq�I����J��0��Q���z��;��>�l������ߙ�L��G��;�T�o\�״�}��e*�l-��R�+~vv=�{� t��4�mד��n��7�]��hvٚ@.��Q���{}�?�u�(��k��Jr�E��W����bo��Ϙ�׺T]|�$�������3WP}�J���f��ɉ��I]��N��E?֥U9%z��@������ZC�1�c���~��z�=��(�!�;��.���f%'bד�^����'8���?G���x�m�+�bp������o8��:�2;E�5�����=V��Y�z�\�۱�����:""�Iv�q���ҍ�K�B����Pvx׻�!?#�{��U�ńN0h�.�q�Wn�ij���E~'ukr3�������T��P�,����uX�F�,�����޴9��m�;vv�ϡ�o�}�f&kr3Q�s��ݞ�˺T���nKͯ�&wLf+�:�aMnfT�8��#""�d�'|z���N�� �7>x�_	�p�*l�i	����>�إ4+9ѯ�ukr3q���۸�6��?���z�x5Á>c��]Z�Ө�ݢd�����^�[;��Z�S���߇�(�[;q��E�X�����v�|�_�ŵuaH��F9�2�#""r���e>%.Bӏp���S~��g�õ���k/:���[ס�r�����1<����)����^qͤi{��8����f�9���Em[�y�~����_7=Lf+�j>�ؽ����)Z�)���8���[o�|��H�����c���ɋ�u��G�SA[�c2[E�н�p{	O����q:�&蛗/�����]+�pv��gn����I���ǣ�S�����y�K��S�6Q	Or$vLꈈ��i�3n<<Y{�`Ht��Še�GNy����f��e�C>_���?g ��������>�o�t�pt��k��E��!f�)����yڭ'&��c���V-�Zw��ޔ��q:��<���1�#""zhMn�O��bP���%�2���ِض�N^����VwMf+�s��yc=�7�c���'١�Se���uAٻ�S�x������K7<V�}�Z[V��������N�&�n��`&vLꈈ�Z����}�!���'>���)�P�ꍎ�!���r3`ד���k{���#ܺ.��� BE�}����D��)��L�;e-ݠeT�
��)� ����{��&�O^Ĺ[�x~�㨯��J&I#X��:""��|�8��<�����s&�}����{>�/��8���4j�=鲒��F}s+NL�����P�N��n��7��^!��p3#+9ѧ�)e�\غιf�����7�!q#�cRGDD��/�߻�#	�}�>�qJ���n�''>�������OIK�6¨<2�<�n�1x�as\�u�&�����Og����2��Rh�:����DDD�|�=���A�׋��n�&����Lh����۞�^���֮���7�M~F��]=Ϸvz=�-;y�J���Nt��mV}��-"��lŁ��.�/���XG�醍��Wx�xs�xޜO7�K��{��a���*�>6�:"""������rm��E���7����h����ـ*%�u��V��͹W���g����+Q8���uR�671��]���﯆.^�s7��V5皰E��b�*������ۢ�5�tS��H��4��S����8�p��/o�k
�6$$=�;N�$""��)Oӹ�g�N���ߓ�/��r���ـ�]J���{l).�u5�u����Vv6�c��+)�����K٠��/�}+��@V�܈M��)�e(�I1�I|����w���x�N�ӹ����M#�2}.�W>�}W���u�����"B{���je0�����J]�ߚ���sq��]���lG�{Q�&2$�;&uDDD>2Y"sO����~U0"uj�/�G�ur�ٻ������y�X����5�b�]�I��k=}�&o�0��[�9G'i�����:"""r�Te����Q��Gܧac�P6�&�/�y)����1�#"""')׶E�Ó��5�vEl��W׻��I�X{�I�EJ���N�׏"���:"""��s��\�ʛ���ͭX�s#�����BY�GAY�8p�":�ݛ��1��S%y�[����]��8��m4�v���7�T2)���qK"""�g���������� �"l��c�_��&7��/��0�{����u�ZG�д��}o�Y''�J~F��s�Ө�����-&3���<r
�+�q>&��uR���[�0Y��o���F�] �0�#""�o��z��Г��V����Zq��zr�߿_�s���������4j|�ڞ���_�z�����WQ��󾍫a2[�*a����N���66/_�|,н���F�씩7|i��Өq�'/8�4��������E	;N�$""�o�n"m��6>5�6�M�Qc������ƛ�F�^_��y�`&;yj��E����|�V9�vs н��F)v�.X�a��/۠T�-t떩Ϙ�]����B�ǟ��Lꈈ� �6���H�Ey(�ٹA��ʵ�(�db�2��ٟ���^T�<%��C�r+'�ي}�>q{,н�<M���ٻ���;��H���e!"8�Xp�d0�f�T�2"����=A�dfrj5�����`������cMrƐ��(g-r	V0Nl.��E�`ld���ڒ��R_��;�����[?���r�~��<�H����<�'Q�wK�_P!ъ6��  �"�bf�y�g������+�,��mј�#X+y������ӽ:`Ц��X�t��e,�^D���'��x��We4��Eya���F�;9c���P�/��h�� �+����;k�~�"��Ƶz���*��灻�g*<r��:?ҭ	��P�7��;^xY�O�;��������|v��dT��<sf<{�S,����7|�p�$;�����=�Ԗh��Ǵ��c������"v�:  �8�L3O5�)+�k��BvݺV�xP^F�v�yh������*~�a=s�����zC>�Gό*���3򔌑:i*ܼ��3�źw�ۧυ����|5��=q����w�=֕�ЁǶ�ÿo�-�Wh��"
v�:  ����}�����0Wm���Ѝ��<pg�ih�Z��f�7��ĝ_��o�ᕤ'f��3 X�蝹f+/#ݐѺ���z��>l����9k=Z�{ׅWO���
��.p"M}mF3���c�C�?��zC����p�`G� ���'��ւ���I^F�<�=��N��h��%���myံ��i�?[^8`�3�����Ϳ�k̺�x��4'�>�A�g�q�'"�jj��oה��4�y��9}oe͠ue+�Nen�<�(�����k�`G� `�h@�����*��{]o���L�ڞ0&�u:���sa�9=m�C�Dx{�F�9����!��}�v����F�֕��3�6�,�軤����/��3��̙��W<#b���ٜ�	=3�0N$fO5�kK�|��P �4m�����i�� /}垘*]:��ㅗc�s]�
Â]����Q.	�f����HK���~L���-}�7�nH���_?6�㼌th�mT6���j�H��_?�����;��>o\S�[W�b�F��=�ˣQk���hb��hԡ�C�`G� `��_?���n]kȺ�D��;j�+��x��ԉ�K��r0����6W��z^�륦k�<=�n��~����������״��A��������"��W��{oW�_�3���N��hǈ�3gf��ٵ�`��޸Vo?�+������S���#�{�o��b!�5Uj��%=���k���*������I��
��l۷o��X,�jPzz�HFFFA�������1����n 9�ׯGn�|T?`�}ӵ:;�S�a1xx�Z5��ӵO���P�ק�O�j�>'���}�����7]�W?�X�/��$JMY�~��;��f�꺽o��_��l���u�Z=��u��Ks�tq����>�=��>�{n�TinV��nS}M������ڕ�.-TEQ��33��ժ���#�~^�޻I����-U�s>�=C���r0��ݖ����{'㪜�=�ԵEya���F�/�^V��3�uin�vݺV�k��۔�f׈�#�קue+t뵫����ڻs���s׆�{��ׯ/���G�W[�����>���<U�j׭kuནQ��a��H��?��:���Gkt�z �L<��Q����c�o�lІ�Fx�+��<B���:0k�ቾKz�翉�o�?���~�E~k�Jb��tOD5N~��g�[�f��Q��Wն�Ks���e������z=��=�]�.������R}MUܣ�������k�J�|T:��U��ը�jK��Q�o�>�/,WF�~	 @8�=��}ݳ(�h��H�+�9�;�z��Ԟ�V�+[���_ZU�btRl�fk��̜j�oP#좩�:�ξ~տ�ꢙh�4Li��x����%�k��:�I
{~���|X��a�%�<�_�Չ�~}m���Hm��REa��>����5e%:��v�}ӵ1]����O��;�j2����nԺ���gS�Go\���ᾘ]g_����1�~����L��ghT�>���rm��ڶQEyq<�קW;>�ۧ{U��PuiaT���������z��.�^��FO�:uqHwT�Ϩ����麇����;��y�1W���?����~,��-U����Θ2��{'����bj�/˾}��V�T5 ;;�l~~~l�u�<��N�R� &�̽���*SS�JjY�x�+MM����bL�,9#.����[I������g�rS�{�9�	�j��%m�6���;�~���Ж�r�++�-�W���y���:���^C�_EQ�*
��N�]ZS8�SQ��'�U}M՜"1�t����̙��-U�:��v�e�����W���[,��0B�<B�x��a;Z�=��_?jHI��l�Z�}_�'�}�b	,�M�g�ߊV��SϿ~,��Έ>z��o��C|$����3>v�'T���'�YXغ�Z��dF(
��x�xlFp�պ���|?�B)  \Ů��z��]��>������h��I�t�C�����z����W�-���
sD��(O��G��{�^:ܡ��ް�N��V��{o���^~�d�]8��> S�e�1��oI��� A��a�c����k�D�%�u�����1��U����J�7_רS�S
������v��ۧ�E=ʹ�0�J���1������^��{5��,d׭kC���	}󧇴��
U�{ȩg~�֢�����+[��L�N�]ҁ��3F�������P�%�P\�#�tך?�������望�R�����ŢQϤʬ�����������d��D�����=8��!��]�᪢0O��)?ӡue%q�6�f���L��<pgB�v:������#ij{�[V�PEa��T�6$��R�>V�uh'�.i�C��X����5}���=���?���z��	�0�/$��;!��`���4����nB��Z���2?}l�IW_��5.�<�H�J�sT�]���옟c�Xd�X�i��б��9���co{2�軤��^5<�m�*��pF�����vEy�(��at"%3�IS�58�rv�x�u"u*��f/��H����v�?��g��7�r��ict��H֬r���d�Ŀ����gҫ4�'�j�ߍ����?�G��0��A��x=��H�O�����jo|(�s;�]T]�+j}�A�U�QS�5���
2jo|HY�k~E]����}���˞�#) �,�H�W�#�u~�1�R%Q�.�^��v��FB���W�����bڠ|1y���)A��SL��(O��{�*
��o��>�k�����:�w)l��p�G5��U�r�������{����g���{���W,�=c���@@���# O�P��b�U@u��'�-�: 0������oPS�fu����S=3^o����,�W�Oތ9Ѕ��9tV�.�QFf��)�)�[|ۦՋI0�xl�)<���pGB�q�ݓ:��o�>2r;�X=���{Be���[j���Pn�Z��¼�7�Gb�^���7���?c�����ڦIϰ���~`O�UzF�����R�q���X���5�c��O���O�z�Ԝ��7�q��?���"�=[�O;�W���u�����KW���-�/<��EO�-ȵ�,�@�EJȲ3B �Hǹ�*���f~��Ӱ�35J�s���7�����k�[7��z��O���h�!m�Xm��3%I%�*��9tV}���▘��L\Y�d:�wI[^80���b��ׯݯ���}��}4{m�b�!���t�����Ӫ��im�*׉�KZW�bN@���\{tL�n]Z���]j�y����e�k�w�~߫�փ���K��&<����I��ǆ���#�4��{2d:����g���뫵c}�Z�ר�'o��~��j�'�%C ���,����j������%5�>���b�6�u `2-G;UW�F;�W�y�65��MՖ���~��F����yNN���^5�xኛ�;ߩ�K��h�u�<ˬ���w�Q���3��YО׏�dDg��Ѯ�U_S�=ܹ�G�9%5o_�������ۣ=ܩ�����-e+B����:�}�o����GN�jW��9Ӳ��{�Zo�
�W����5��jxxX��.�ᰫxE���	oC0�u���h�%�[7�q�F5l���x�`�t�����n'�k9 ������l��F_x�EO�mͳ[�,ғF�S"��)�\æ�?���͡���fW|�Z]�=���ߑ=-]EJw��n��bY>�)����ۧ{��;ݨ�����K��gm�����s�}G�����j=b������E0:���A�^~�d���=��yL��~x�ywG���،-&��	�{n�F\�P��ٕ�?|����Ј�3c����B�XW�B������p�{|�����*=q% �t�#������d�    IDATu�Z=���q{��/��F����v�QU>���!g�k>?ӡ�wԆ��{��A�=����O]��������Lӛ�Vk�Ƶ:r�wƿ/����S�?]o���3U�����\Ymv�9/�\��UPP���jY,���,;�W��zMh}�l͇ޟ�~�?�Pæ��3[��T�Ԛ����>�:��.�)c�V_|j�)5�|co�U��w�&��	�<jz�jy�>�>����o����%��b���Z��z䛼�1���̑�jU 0w���D�%��{U�n]�g�ݔ���>:������,#.���~L�wLMI��Ji�s�'��[�jM��W��Kou��;qy�tO��G�{B�5��XÕ����w�N��N�vb������{u�T��U�umQ��T�Y����_dL/��j�F\�}t&��	�軤k��gs�jm��SI�s���ܢue+f��RU�-/P���Ϩ$���\�ۯ�wԆ�o����ޫV+?ӡ]���V� �1����{�O�5��j{�Ka�W޲z�v��S-�`�
K箅��[������wy�Z���Ӧ���z���{~�8I�����ڱ�zN�kj;��G��23���w��uz�᫟��~�5�[{��~k{��.��� ��h=~*���k`DMmG�ކ��J]�N�I��^�vISB�=�_O����7̎��=���;�[�s�v�?���t���=�_{^?��~��?~C����]Љ�Kz����tʗ��`��/�����go71=��>o�u|��V�	��k�TQ�7��#��ծ0[\l�Z�-aF�wm\��53�`�e���0O�gmi����ue+tǬ���j]ي9[`��^�k>�aij�qKUy(�Mn�鰇�|^v������E8�7�5���]�=�Iψ�3.j�K�50r�"&�~"Ia��I
��;�ھ�B��������}��k������� ��*��UwcE����	M��e������}���'C0�m��ӄN�
�GZ�T���k�+o�|�e��#w��)Q/�Ow���=�I���1m����m�茜�ۇ��u8�����>����u|�J��3��{/���+����<a��=�Ԉ;�}f�]��.�uI���z��M�}��՞׏���j����[uy삡�-�t� ӡ��]�Ѱˣ����V�B`����eFH#�G2]���>�ᗿ!�{0� L��������Tæ�P��. ��Z��e~}�{R�%��ͻ&imX��>}nj-�+o���JwTMM�="���Q�軤{/��ӽ�v4.Z�~���#�u��aG�"�tO�����a�%�u�IZ��T������-/���u�	��[%L}���g��qy�ďߘq<�����;Bk�z�FC�ئ�������{d��C#d�}����ȭ��}8r�W�=���33�����I�軤�_?�-U塯���P��S��r�x�==��7B#fӧ�N�{�k�v�릿�g~�������N=�ũ_���/���J��^�k1���U$�?���)+w��3c�w*��ڎ��z��nP��݆O�����y�.Co��~�5�/�k�B �PS�fՖ������t��M5j�����%�~�?��m��Hekn��s�9��V��V�#[nט|^��F�~���p%�}��� ו���Iq��3�O��m�EX*�jN�]҉�K3ʾ�*�_���<:����S��{�vzi[�i�{�\hs�`_x���:τ=���^U��8�����K�;TQ�7�ks�+o��׏�9^��U�+[!I3B���9>��h��������R�=�{n��\)|�'�.����{|�s��~�O����zo�{ZJ�N��is���3���SZUPF����;��L���݄}���B�4��)���O��f셧Z�a��^S�����:B �L�7�]#�@��YW�&T9,�i9Z]�Qc�^��=!ɮ@�+�-���IҤU�u�O�ե�C������42�*#.Oد���wΝ����FL�;>�ߍh�'��.��ْ����K��>�Ν�@��(�`�q��ר��t��\Fp�ѷ���z�ڱ�Z�[7�ն�<���@��ŧ�O�m�X�����5u `"�������4�o�w=B2X,6��W���MZ��Z�y9r��]y�*i�my  fc��U~�t�����+��5֫��Sr|����l�E���;��`�Y	�׆G��x�Oޜ*f���@@?OŴ��F_x�%��)�: 0����?�@��Ȝ�d���Q��g�TKs�++�L9y�dO�Qzf�` H���1]g�ٵb�M��s]�kt�3y'���M\��i�[Ԗ����9�k�[7���!U�ݣ.�a�'��ymyiT�	�o��}�D{�/�$�nm��F6[pyp��|�E�b��]�:#�$t/�ͦ�K��
 �Q^����^���Y�Z]�^�44����S�P_��}v��gj}�����WN_'���������F��9uk�f�Z�-i~kTSu ��4��w���C�G�bY4��e�Q8s���>Y'G��d���2r�W^�_���r����'$���� �����ʟ��V����r��S�K���l�Z��R��oC��?Sæ�9A���)�~�ID�.gk��k����y�uF$���/6���>Ց��G�)�B� 蛿����v  ���Pqh��O�d���ҭ�Ϻ�d�ov�+���ۡ��٣���W��Ψ�y-��Nijf��A��'P���J���e���N�   ��o�98��')i�Y����T�a�@@B  @d�wnU�j9ک��|Ֆ�������8w1��A��P�  ,k�?yS��^h�W�7�*�P��Ў�Ւ����k��Eiܻ��_F;zH�  �Gp�dI���"�R� �l�:  "P����?}]���uu}���T燞o�nij�)x?D�����H]æ����Xܲ�Muf���uQ���f  ��L_s5}J��a�G]#j�߬���<�n �A�  ��~�g��f�~�G���
���T7�T�O��q�F�%*�Q�d�X�=$� p�奪-/���~Iu�kTY�0�`�z KK�*),���t�4  �*��r��O���Eu�����R5l�YpS\�K��g|<}ۂ��fǹ�Qm���P����������!� �G��5顏�'s4�cW��snN K9ʊ�A�F=�*��:q��y$��%Ip=]p���������M5j޹M�z��vD�;��F�Z��RÏ~1�܆M5��;�]T��筴���y�R�^k9�*�_W�F��?8����FT����q�5l�	�D�<j~�9�g���HS!)�`��H�9�ػc쟟jMu[$��6D}M� 0��֤���B[s��W�y��*�,����Ue��(-;��X,Y,}�y4t�du��e���r;�WOU�tyB��Z?�DM��U����d:���}3�Nנ3���6��-/Uˣ��dD����T�,�t��~��n����v��ᦢ6n�0��'o2�`Q���E�����: �~߄��㲧�H
�/�2����5��f��$I�w�*v���T���h���Kp���G���G���Q������7�	{�VY����|��TS��<�,�W��m��^z��p;=��<jj;���ҩ X�F�;��� ��X,z����JϋOu���O�m�(����R  ���:����х�?�u��ώԨě�uA뇟�x-P")���v$t~pM^A�C��6J�褩i�;~�3u$Zjp��� ����BO�ӧ[����f�ێs��?M�l��ϓ�  &��%�xro��bm��RB �X{�C����io|hΈMp�g�f�M��n��?}=��*�M���;rUZ�N�׮Sz����a���N��|m��=�(S��S��s��pU�n�}��|o���.OJ�,�{��
gӿނ���h���a��8F ���b�]9�ػ#U�ϳ[�b��u ��Ֆ��Yw�~�G͇ޟ�*����\���q�b�HF�r
oP~�-�)�VNA���t��*\q��ӭ��i���,���٦����p#n�Ey��F����:%��g��CA�#�j���f�����*kKַ�&}���o��a����z���"Q��~���`�kܺaF�hj;Z�4�XGA�#4:��r��׬Յ�:{����UPT�tG��v�,KB��l�������
����N�,9��^K������_v/xn��{�0��o�Y[���:���p2������V|S?��E��'o��TO�����$��~s���TY����#	�XlZY^��kV)?7Sc����Z�η��(]�� ,N���٬�zroA�������v��=�i�A���	̷n���E5�QS�f5�ܦ�㧴c}uhzf���W�f��y갼^��m��iF�R��T�Y�[7�
�DZ�$x�|�۫�v5��>:7}�n��,�G �.����p��Ou$�9�ػ�귶��$F� `Q���-/U��H��ܤzz������v�,�����^�ˋ{�H���¯��n���lAܫ���t��Ia�x�����)������0�E��~k{���k4��O�-��Ƌ�6YfD��u �ht}��9�/���xhZ�BO�����{I	
rd�PY�M���I�:/$�ىڛ�T�UGނ{�Iх���B�nm0�|����)\x�Jiz���BdS�fISm&�0��o���=�b{�7���{�ܧ�6�٭�E	�P �\���5������a"�k��~�&''599)[Z����,�P�z�vh�3.Ir�����}Ѕ�?�;�pQ�T��7]��eO/RM�N�mܺA�;���Xmy�Zp�)��+f7jܺA-��q��r�30[p�{��`�kz�Ii $�Ţ���{���ܧ�6D�������ܧ�ט�����~�t���cM ,ӫ_�X_ڬy�=���@װ�&�~]������5u���rTV�gs��|�	Ym��y'd���3��j�Hz�����t�i=~J�WBَ���/�r�S�5�o}�k>�~�Ѻa�G�o�*�����3^�0F0c1���G�Pˣ���8_�;���q��� `f���zW�]�O���@@����uM?���Z,�JTg�h����}�: X��S�ZP-�ާ��aGꂁ@���9����u����b�)7�B����h��#��s�5��Ž���Q�h��CV�`J��z_]�N5l�	��u��Z+9��p�u���h���צ���8wQ�����nPæ�ｩ�Z?�$��1 `&��Xt�d�;�1��$}˳�۷��j�J������>���o�$�\�g:9�Ju3�����Z��z���4��}5���Rmyi�}��nPS�fu�����9��>���F�mGB#s�jԼs�T��W"j��}�Jݔ�ٌc���O٫bzO�M�����^������ׄ{0�z�d�������  �+���"�|���u���`�����T��Ֆ��=Zc�Xd�Z����U��5�/�I�E7�jK��M  `&�_�"���7����6ը�T�Z�����2�n�������oPæ�?u�i�N_��kg;?�urT�Mv�-����z���eM_)Gza�kpBҙ�� �rE��E�k`$�^���?W��ݡ���~v�װ�35%�J�pS7���/Å�?�  @��Kk�R�5u   �ǚ:    01B    ��    L�P    &f/))Y��������8��=K_q�D�   ,Q��   ���    ��u    `b�:    01B    ��    L�P    &f�t����1U���^��>UϏDFFFaFff��?�����⾧;@�N�7�M    ���/�גnJuC��>���������z�����O�    0\    &fOu ,]��"��ޛ�f   ,i�: 	㷧�U�2��   XҘ~	    &F�    #�   ����   ��T��@C�o3�*=_�P�j��G�   `g?PqW����Oߑt�a���    ��q�u}��[
�.���wT8h�h#�   @�4nݠ�m��n)� ���   @�d:����*��P���Q]�]���P    �wn��e��ڎDu�RtA�;
�    H����j?��5e�-�@T��;�H�S�9�Q_�H]��Ҿ��6    fm������d����:B]n���Wz/|��v    �lL��P���5����:9�Nus    \�V��U���7n�G�'���>5�E����f����T��^��qѰ��F������댮R   ����1�S+W(=}n����ٳ�
������46��ʕE�?�T�~��ϝ�P   `	����a��:k���w���+Q��ΟTaav�����$���    ,~������y���|��~6湉t�R    ���   �T?�E����0R    &�H   �%��%τwƱ4�_��i�}���<�3�kKK�s%B   �%⓮:qp�q�զ��I�	X�t}����<ע�Ң�<s�s�    H ��:I��}�8,�w2��1?�2��zn@}���O    �����#8�'����3#�>���:    01B    ��    L�P   `Q�_q}���4~�M#��b��P   `Q*Z���nKu3�o����wk"=+��	u    ����t�   �"�T���N"�   0���
t�   �I,�`gd��$�!w   �$*Z-�6�\:�����ut�   ���^T�k$�͈Y�ؐ&�u    �������+�͈K��H��ʨc�XS   ��B�����r/B   �Eo)� ���   ���]���P   `�Zʁ.(�`G�   �(��~��]P��({l �k	u    ���T7!��Ƈc��P    &�>u    L�s7��]��d��o�n�:O�׻|j���F�   `j��4�tj����ύ8�=:{�W���S���u    � �ΟVaQ����!��w���+1��R��?!�   X"���;/��?��?��f�
�    ���    ��u    `b��   �d�����8�f�+==mI>W"�   X">麠���Zm*+-������熞�л   @�Y�7XI���S��ay��K⹳1R   ��>>}>��|RO�x�l��   ��1R    a��7�aS�
2�Q뇟���H����0R    !�wnS�����sU���ƭԼs[�[��0R   �p�5l�Q��Sj��/B�ZP�j��vD�.ς��_q�r����ܔ�[m)\ӵ��   0\ݍ���?	vy�z�Ԍ�2T�Z]�ݖ�."~�M'o�[�Y1]O�   �4]�Ψ�_��.�@'�    ,rK5��$B    Xj�Ψ@'Q(   @U�i����;.I�w/X<e�h���T��;	ik��$B   �j�����"THe>�`Wr��K���m0,�I�:    	�q��5���h�V~�Gu_���G�   `���5�1��g?Pq���M���.y���[}�!��P
    SX
�.���p�א{1R    a
2j�T��?Q��H�X㶍��^�a�G-G;���n)����/�]Y';B   ���-/U��� ӡ�Ag(Ե>��j�KC��U�QSQ޼k�b�2"�1�   @B�<z�$����?�$5nݠ��R��T������W�q��mTA�c�=�r�������b�    n��jU�����|����su7VH�������P���4���z?Z�.���w�=6ӵ�:    �N�l9�:V��P]�u����))4�W��1��c�Ih��5>�u�:    Iz�zRܒ��B)    7|�-I�,�m*�c}��?�������nX��6W�f�?޸�u�<�w?�4�g,���F�   `��h\��jz�*�th��ju������.�<@s:�re����F����=۫@�؉��z�l�:    ��8wQ-G;հ�&4'MU�j޹Mu�kTY��+CL    IDAT��������u���
��e��Q��[~�_�Y}����	�   @B4��Mu�h��j�<j=~*T8%8B7�����3�^����;/��?��?��FI�s��    $L���n*>���G�P��S)h��B�K    	S��PS�f�U���Z��j޹-��#u    ���T-�ާ��|Is�T競�T;�Wk�~皺勑:    	Ѽs�*��`��ޜ�+����vD�5��f�3�]�pi|Ɵ��IC��+1R    �ר����EP�����5nݠ��5qmL�I���88��jSYi������zNB�   `Y���B�B�.,��&Z�V�����wqX^��#g�z�l��   H����50�3>>}>��|ROo\�Y,ϝ��:    ���`���ω$ b.B    ����X_}�s��P�26�:    ��8wQ��O�q�5n�0�y���O��U$e9cM   ��h�ɛ�,�WS�f5l�Qǹ��tJ�*��T[^���|u�����6����m�ڏ~%�ߗ�'�Ǒ�K�T�t���,Y���[g��P��   �IA�C��6j�-7�Y_�50��?Q��i��	{}���%�<�l���ޘ�'�E�P   �'82'M�H��-�`o���~	    I:�]���Dz�N�|��vF:�P    
2Qo&��q���0�Z�3*�I�:    	Pwc�Z�/�k~��?5��K%��$B   ��8wQ͇ޏ���	����bmZ��Z�r>J��R    ,Fl>    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01{� s����5=�RZz��2?�_#���T�   0�q�8�У���T7e^�/_V mT"�  `	b�%�666����T7#�˗/���?��    ��:bllL�������������@��   $��SZZZ��2::��&    	G�ò�ZT�e�l�,G�N��   +B���4�ʍ��YRR�����a�   bE�    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &fOu��
3��ސ���C���ci�����|�c��n  �]y��+�R݌��,�zzc�k��
=���X
c�����f  `W��T7!*�:,�>cC���   bŚ:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� �P�f�Ck��_Ia���/v?    V�:,�t}�q�%9��   ă�    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� ���Kg\~����v/    �:,�~}�g¸�\2�^   @�~	    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���S�  rm�Zlܗ{aN��߳#��   ��n�������F\~C��?i��%�n�=����\B   B�2qflB����o֐O��   @�XS    &F�    #�   ���    ��u    `bT��i�|>��n��~�l6eff�b���Y   @R�`J>�O���
�$��+�׫��\�   ��_�nw(��|>MLL��E   @j�`J~�?��   �RE��)�l���   K�����)�u�oZZ����S�"    5(�S�X,������D��%�   ���e�X�p8":�������۸�|θ{   q`�%    �#u0����R݌�ݮ���T7   H(B1>>����T7c�ϧ���T7   H�_"n�5�I���S�    a�C\&���-(UAIy��2��_�Y��n   ��:�er�u����W5��    	��K    01B    ��    L�5u �����A����n  �p\��&D�P ��seU��  ����K    01B    ��    L�P    &F�    #�   ���    ��u    `bl> �jJ��o�ָ�:����g:�t/p%¡? X~u R*7=M5��r��c��e�m)l�yџ  ,?L�    #�   ��1�@T�\�*�՘˘�YΡl��������\.��*��D���ONhrx@���2�{%B�k\�?9��˗��Ŏ4��o[���CǼ^�F�n����}�I�Kc�C�>�x��  ư���r��VZ�����+*��\Y�7�\s��ۍz<�(���u�~-��-��<E7����ؤ���T7e�  a)��:��~(�m����T>0���n���oVVV�$���L�C.�K����$��ŋq?o��d�gFF�._��,� ��lY����<���'�===��'�a��7���v�r�-��?�3�p�*//Waa�$͘&8��������&&&��ե���9sF��c
&�%�,������ٳg�D ��-�PW\\����<��?�?�KA�$##Cw�}�n��v�|��r8��H�|>���kddD:y�~�����O?���"�'  0��`�C�xV�������l|��SFA���Mx������!MK�XȪU����k�ƍ��Ϗ;x,dhhH###�����~�;���Gt]���	  �Pg����r��p�je���z�r�\���]�����٣_�V2��4��U�V�G��͛����@ ��VNq�\�������~��_GF�Db��G}T_��Sڟǎ����z� ��Y�.Uk���Ҕ��-#u���x4::�����s��r:�S%�P��&�dggk���)	s��\.}��gr:�:x�;����
"�'  H�e�R���D���JKKKe3�˥��A�^�z��������'�۽dB]��n�����׾�5egg'tZ`��N�z{{500����/X$�A$��|�ǔ��C ��-�!���C���EVV�#u&�~�����y�������D��$�.q" ���z��'��C�f��t4)�á�������v[(��SPP ����ߖj�4�����	  �[�i�P�x,�Pi ������|G��r�|>_[�ժ��Y,]{�*++����Þ�� B�  H�%�6u��ru����K�>������h�|������)�á�7�>�����"�'� �d�,#��E@�mۦ��~ZYYY�	 A999���T~~��y�egg�=���R��O���b~��'F�'  �:B��E@�|�ISoϑ���믿^iii	"��\;  ��	���������T61p���ʕ+<���������Ą�_.� 2���ҙ3g499�={�h||<�y�Vq�?��O  9B]�|>edd��΄&''5>>����ϛ�������7U��4��]�V��������$�.�Ad``@���w�=/� BN����VSSӼ��  H���b Q�$���g�UVVV[����*++Sqq�{�y�N�����9՟��'  ��X�2�� z��'URRb�"�*,,T^^�jjj�iӦy�+..�Ĩs�{џS�YXXhH ��� �q�}���n[������L��k׮y}a���5�\#)��	  f"�����Z?�pؽǖ�ͦ��2����'�H�3�[�Y�&��	  �"�����򗿬���T7%irrrTRR���r�[���{/�����LX ��u B6nܨ��k�O��k����Z��G,�Oc�  �G�K �Ͷ$�X,Kv'�e-##C;w���MuS��f����D^�W�a�=�Oc�  ̏]��b�hrrrɭ��Z��X,���,��V�|>ߒ�����jݺu���HuSR���D������ׯ���G۟  `~��
Kr��|��n�+==]�E�@@~�?�-C��v��o߾,G����K###ڴi��=��Oc�  ,��0�����˗5>>.��#��*�����5�\�[n�e��"��n�q�q݇��bT ���>�/�$��jbq����+�����)������<]w�u*--��>����  ,�P��
r��r�\��wX\���USS�$�
�"??_N�S_��c����)��  W�O�H
��/�˥��IF����UWWS�押�<�|>�_�>���ϙ��O  pu�:$���._����ȝw޹��~Mg�ٔ���իW+;;;���ϙ��O  pu�:$] ��c:fj��v]{��Y����v��nݺ���?�������X��	  "CiB�������f3������:+oKQk"������J���Ѳ��u��]��Q_G�k ���R�gI;�ͦ�˃�nF�


�f͚e�A�|rrr$I7�pCT�џ��ڟ   2�:��R	vf�j�*
z�#--M���Q]C�/��  �aA�ǣ@ @�$#����p(///�k����ҟ   2�:,���<�iq�+--M>�/�>�?�K ��갨�\.��K"*5�/==]n�;�u`���b�O  ��aQ	r��
)�����jrrRn�{��&''�!   )E�â������NA   ,Z��~�=`�w���Y��X��
��b��D��P�EirrRiii���LuS   ����7�����w���?��X��m$�ٚF��,v%j��P*vQG�W�΋�焯jܽ�(�!,��=lv��E�[���L���oþp�C�2��]j_%G�nD'e,%��&��-r�^P3�(��ΐ�~���4���cZ���{� l&r���Ƃ�~�踽�b�
���Cz��I�;�Y�2�eɿza,\�/�ŗ� �@ۙq� �~��;&udZ�t��:"�K�����n�0��,�?�����x��/����u2��u�_���Ů����,��?h{��X��v���Q-�`�K2�Z:��j����Қ��Y}��E���Ç��Ԅ۷o��1���ʙ�z������.ڛ�����8��gB�Nf�g_�_�y�,c:-Jn�:�ű���Q_�	Hh�� S�d25q���ں�k��L�ϬVVV��imll�b��4G���ʙ�zu�DU�?w�/!��2z �^'s{��S�1�����WǦ�����PZ��Z$v\~I��N����Oj"i6B*�*yo'糰r�^��_�k�o����Bu���y�4I��dV���+3������X��EI�:6�rn�m�İ t��<L�X<G*���e�Ւ�d����d2Y��8�;+w>�ٕ����P��ש��@"��<�H��WǦ���Z �U�s�#e2�ZY�Y���8��鬭e�A��Ζ�8���ʝO""�j� ySǢՎ�r~,$�}<���2�,��èK�D�h�Is���U�۷��~I��|���$""�&YƵ��c!��/�%���x�A����_��IH���U������|����<�̧����=""��TF�:��cqY�|�<�wT�GI?��կx`�L&���|��Ge=�����|�t>��v� pr�β��Q�e�̈e���/�˩�1�#jp������e�iii	{��){�W<�|�t>����A���c�,��~I5A�$��P�VWW1==�g�y�t���.�H������/�z<�s�T4�fao���œ눛��<=��ن�_���{��|�'��}������� G��� 89��cO�  x.mm`:}ng\���h���'�կ{���:^ṕ�7�r��u���W�cj�����ف��_B|-�_\�������9������?r���7��Kptv�s�-�#s[����q�?�v�^Ͽ��焫�K�Z��M&n�<u�#��R��ւ$��K�/-J�=�8Z�c��QM��V��������6|uiccKKK���X]]-�y8�YXYY���|E�Y�o��#��@;:;��4k%�{�����\���y\җ��w����7�:}����������7��<�^��$wv��:  <{��mq\�]����9z��7կ��=�n�w���I�u�f�/>���|/����aDc	�[���-�,N�xsW��v�d���x����W����z�����\���Ww�#��� w�͒?�*�ukFF���K�:6�~�b��s���j�,�쀩�{��arr�����/���}��������|fi5��8:;��߮��;ث~R�5����]�(����w5�I�_K!89O�S�R�G���l�;��0p�&����V) `j~!{��G��;؋xr���G�_wtv�7�Z���:�[��(�����$��������]=��ȅ�#��QJy��d���ϏB[ө�x_[MZKQ��֊,c��w��D�I!�N�ʕ+��d2<x� ���wiT��jm��ZΧ�n�Fpr���7@T��k)����-����!����a���M���ݥ���~���A|-��{GIDɼr+j����|�X��7���U�>'³w�u�f[Y]{Ky�+�'gv\�,-ͭL�F��[+�(��l�JM4�� ࣏>���߰��!�"���I���裏��{�5l���|U�����^�g� �ހۛmE���g�l��M�/l�u;{05��pdnK��݅����b::;�Pc�9y����jUMY������E�Z����lC��mDc���BJ}�k]iε��M[5���TSA�:��������7�7�,��`qq�dR�$d}}?��Op��Q�g��_@pr���C!O�n��$ `oi*�9ów�*���)7��X��.�#sp;{v�KUh�f~����S���yy��L� ��f)	X�����u�N��o���5��K�b����Nv��A���BU��_����������uki5m�嗒(�E��u��3�������D"����w��d2��S5��9�����D���|j;�;��4!pr ��H�^%1+�r�U��H���7���F)��I�J���CM�����Dpr�`���F)J�{����եQi#���MG89�Vn�#sN��7<��q
een2�u[��۟K����L��N<u��%��zݴ]c����ӨKت-�N�ҥKX\\l�����
���055���/Χ�{颱��u��=�})���%�?+�U��(��q{�S/��ei��d�ꏲG�X�����rM�1�����-I���N醩�2��Z*۔�ن�<?�Gm���K������J[.�<�xr]�v�sn.��V�s�����J}�Gc	��b�[k�V�tR"Qݥ\�J�.���X,����A,3z8������O?��������|�'p�fիc��&8:;ؐ��'gԆ��	僃��������V�$N�����Z
���E��q�G�mk;O�S*j�+׷��
�:���E��|�':}b[�47�*�� ����RI+t]9˗�zݴ�:�	�R�0�p8���Y�����O>1z8��x<�믿��9j
�'Q��_��M�N�@���-gw���|M15��=�+����=Ww���J+��BG�7ԏ�t������a�Ȍ|���N����Y����t)	���+{v�G�($=}�]�J}����.1����䌚�z����n[Z��^�6�ba��AJ�2�#�mdY�ݻw��3�`qqKKKFIs.�}}}�Z��/̝�D"Q��jΧs�؞(�P���\  BIDAT�)���\z+[�x�Y�#_82���;7;��t�������#�N
5J�M�	��	��4��f*JI�vJL�%������<�_��]R�YS:izLh:�����;>�����^���|C�p9��1�끫7�<����׭�R���.��:u��!��j�j�8�r� @Ū6�H��X[[C[[[��666 I��կ���s����E��{wnWl�o����G^��ֆ��&���u��9���Kx����o�vyy�}�[XO����p>����
�����+�������������/!�+��b�`o���+�!Kd�[��|�'���qQm�����Q���P��w��_��V���,����hH���hii�7��M������0zH{�'��/����ʾ�\���ػw/�S'�f[v�[K���t�;jz����� "�mб��g��X�� �U��>��/�����X���Ckk+�}�Y�ٳ���T�'����Eww7~�ӟ��+�q>kH|-���f4��c������Sy%"jD�\z"�#o�`��L�	�9ܻw���>[�&3% �������B��7��>rP�6:5��{#b��߷��;RǢF���̸W J>��I���j��ޝ�����~�ݻ�������n��	s�\�����'�|�4	Ƚ{����Y�����i��ԛ��R��WΦS����g�N����v|���|�'tI���ID�a���JkP���q� ��rʤ�L�V*u+++��ں����yҠ������hjj������֭[�����\���nA�$�A���E,þ}�jv>�|���z��&�`Z����o����y�Spr��j�o �'������59H������}�`��{N�@��'{.���\zK�$ˈ�Dd.����[�n��T� &udb{��a�Z__������o���|��)��v��N����x���ҎVVV�L&100��,Q4�@<���g��r�O�WTEs;{�9�=�|�\1�ȱl��Ko!��B��	�G����F\�]�N�;Ҽپ}�Ͻ��V|��1�ȜD���s���cSՌ���G F�}<�:2-A I��àH��h4�'�|_��W��_��Tg���v�����~�3�/�$	w���|�(p��p���D4�P�y�7����BprF��g��?r��.�Ԁ��5t���ߏ����lI�k1&�� tX3b��n\�W#f˹q�(��J��I���je��ܽ{�(��v�Ν;����L&������׿�u|����/~a�X���ԇ����%s�{����;�״>>����%�k���*$v-��]VI���R���Licc��q7J�LX__/z]:���b�Ҩ�I�ڵ��bdd�H���UMF����tbqq����*��,���	�P6��;d\�����X����<G#��ڒ$���_K!�,��B��ē�L,��4�$v�s�^��b�;;�%1XiB0�#E���D#Hg2�WCWWW��'�����'�O>�sss�{��f1r555�駟�7��M<��Sx�����Q�8kkk��Tr>wo7�[ng����-�=}N ����b��U�D3t�6|��>�ݯ��H#������`/<}�-�5���ݲ�3x긚P&n����|ϥׁ�F�$"��Y%1�v����~XVW����7�����.�:2Q��5��$�i�^]�������������a�Z��"�U��455��p����~�iX,ܸq�n��h����q�=t�f�Z�900���fD"ܽ{�n�s��Gf�g�K�#��������	'g*��4D�S*e�/4ѽy��|C����9�Mb�Rj7N��1 ���.���b�<�݈�DT�C���3=A�W�|mgƽ� ���FC �F��2:t�m�Z�=�=A�N�M��/�� �J�����u��˶�6����������9Ċ������!<xP�f4� �w~�w��҂��%ܽ{���H&�XZZ����n��n��'�@WWzzz��ގ��ܾ}��_^^�.�����c_)x�Q���c��/����l���`�����a��=p���l%+pr���o��{�Ww���SO�f��ܫ&�J��WA�:<u��v�A�>'��?�������VFDD��2�ɐ���v���6:��k�xA�i��)X�#S1CB��<�;�{�H$tODdY����YEtuu���v� ��������b�ǿ������}�>��3]ǘ/�L"��m��!]$���OeNͧ�b���>|�>��ABWL��M�:GgGv��?e_�w��f�nU2{K��6�5�#sۖ*�A��Dc��؛mjsV	��A� �+~,��xM�� E%���D���nA@ �:.&ud
� `mm��a4����o�z26����ê!������qUc���C,..b5��M@�������AI���:�sS��Y	-����=�F82�m��lC���o���t@�b�v���Ec	u�`82��tD�`˾�z`D���jY�F>�c���<"2� �9A�s�q�77��*��dRG�cBg�ŧ~�O����֍5H��t&S�18���G��e?���~��}�6���#����@ =��.y���S��Ep>���n�[�89 [U�7���_�xo]n<GgGիb�+�|�yO߲����D��0����߈ʕ��e����VM�}?
��C"z$&ud�zI�������o=��-xʰ���_��aߖ�#��8���(V�W��많j�4��M�g!�X�����;5���bGg���������*B�x7��^Q�2K��7���@��k�臈�:2� �$���ՊL&����F����ެ��T1ng�#�Ԋc�A�z%t���-q�J��\U;���Tٿ�r�!��7�`oiR�\��S�LIGgG�^�Qg[*��Wy5�Y�L��,R��.�߉�1�.������S7�ă�3�7���s"x�8��?�M�n���FШ����\U;�����lSv刊\�X�n>����;ػm)s4�@pr�n^�"x�8<}N�g�����I���z�5��]��=��9�f���}�M������D��_|C���;7��*����	�8z�hL�j!�S4�LB��� D�c��fXͩڮ�&�LWw/Z�h��TZ���*�ĵ�x�����9���8�Z�J�����s�7< �� ³w����X��Q�2�ZO�#�\�~8Q଼hgG]$;��~�G�!�C`�Ɩ9v;{����K�#�gD!Z'�~��TϷ��"�{�������c6϶T��*�� x���:}���۾noi��ϩ���~���^�瑲�AY�`o�m���^1���`u�
�YH���F�n4�|O���A&n �S[�+7��Ύ���t(u4��c���j����_�6E��O�3{�����MGt��f\#*WFV���;eI�N�.��3�*,��=z�>�#�S:�j�;؋���}�u�x89�k�LIr<��R���7���^�c�ów�9�mń�ϩv�՛+?�����f&u�+�ł�����;GD�|�}��m#%		��<|C�e߈���[Yf���;���@��M�JN��Q�j�j��r�\,v���I�J�� �U�Bϭ����X�X�����v�Ճc��s14�.OL�4��� L�y\�������͹��_���S�!�֢���oX��k&L�Hs��$1�#"]){E
-G�7G�~#�v���P<�bdoڪ�߬q�H��L�]�]��>�z�S�u;���P�Z]Wx��w�S��$W��٥�:�+�/�SϑT~F(U�����ȏ�z�5�{ng|C���sh:���F��	&��z�;ث~ �,�MG�+66_�s3&uT1Q��(�2��4R�����r�����rtv pr����_���zc���ܛ&=؛m�A��.u9dprF�O����/�8�ju��FLGgǮޣ�R%�_���q�i����4�k)�.OTe�Bٓ:}b����t����^/��_|��
��]{�������h,ϥ��9�.�ԓ�G!��=puw��ݕ=Sts�|��[��}�m]�`�*�q^}�r[�֫F�A�$X,�AH��l�,�2$IB&���$.�� �J�����u�t��(b�?�����vS������>�]N�s`w)��6L��7�\�u���O�7<�h,���}⮴�w9 �7)1:�"prX���	RDc	]MSI빂��܎�
e?[�+�
=�*U�|��l��Ko�����<}N�g����U�yV�{T:�V��7w�`�_�QX�����2��٣V���H;��|�o�Om+Y���tz.��pd�����g;�uv�]��v�d+�U����N�����}Z��3"&��B3��ԃҡV�_֣��N�7��5?�^{��6ڛmp�oG���sh:�=Ba��g5��V&��z� �1�#"������P��ܮs�P�JwKe����U��[pr��5=.Wi6�׍��g/�S ��<e���/�Sa�� �����+��_���wt�˸�B^[:?�eRGDD5���;�޶?G��f���;؛Mb7�f�S����B|-���͓{�m�YO��3�:(���Q�J(dj~�>'��ܤ3�Q�I�R��=���O��~v�2n�Q:��/�����.O�庺T2�|$=T��?r��~� �h,��郒�j�`�[��N�S���g�s�<0Z��s�'�y��LUc���i�9�������Ҕݧ��Z��p�e�Z�k�܄`RGDD5J�\�$����W����-V��(�l7��	\�	���j�,����ϩ�M�!�@v��w�WӤ.K��YT^_4�@0�:���P?��՘�u�����S[�+���
θ�k��F�O� &uDDT������r�Զc�����vـ����-M[lG�%��^B]���+���[�##�#s������Mh�D24��x#bc�9�z��89�P?B��޻�˸�h�����J$�~Y�x���r|C�r@�w���c��!ttv`�� |��[����&s���e�o�_������j�é��TZ�m3"f���T��z\>���P�V���.O�t�q��J� &u�bRW�����(	�rV�B阨Wg7�X�l� ���%L�����|C��l��=�[��4�<@3P�*���qT�2n�)��L�t5??Q����F �22����+�eYF[[���ˤ��teo�e�gy]7j��r��;��٦&����S�SL�`����^�r��ۆ^�3.��j\-=*������?62<U��?��Ƥ���H�0.��z�J�&� �$""""�0�ƛq�lv���~IT3d�daRT���([\� ; �-�3h�DDDD��R:�I���2�ɐ���pq,^�Ұ�l�㎽�Gd� ��DDDD��R:�I�)�2�eɿza,\�cSǢ)   �vf�+��������L�LE�,��/�0���-_bt<�n�0��s�QG����O�����G_ȸ�˸��5J��3��w\����������x��AU�~�k_S�<�9u5��s�V�&���2��ɛ|ul��'*`��q�1( z<?Շ}ˋp����� �2���D�c���#�U������f��f�1��A�t�,�����u�$��x��饌�ƅ���*�r~,�rn�m��0;""""s�4����j���Ts+���ș4�)$�[�_�� d��XJBW��&���M1�#"""2-:�I��$�3���CF����2�H[$���|�WǦ���Z �U��DDDD��V	� Iݣ��E�~{�Y9?j?{�"���nH��t:���	��={�0.�2n����q�;��L�J�ؑ��2��\)-�ۭ���0�QdY�Ç)$�Ɋ�KE8�2�G���q��Fi�yf����5�:����O?�4�{��w[!^����R�k� .���3�>Al�8��A��bEKKKE�H�_�V�uW�D�q��Fi�yf����%=: `[F"�2~��85z�Ƃ2�0zT�_����ʸ�˸Տk�F�gƭ︕�+���B���c�4z T;��E��/P�e\ƭ��N�h�̸��\z&t@/�$2+H��7n/]��(�H"�ЮY,V,..buuuW�>���(�2.���m[��3��w�R��LꈪOF��!�J�:6�~�b�S���)���n?����q�v5�<3n}�ݭj$t �_U�,��G<��M"""�ZW��`RGTu�(��C>S&�DDDD5��	��������H3�N� &uDU��6_Ǔ�C"""�ZcDB0�#"""""҄	�����Z�p=�|�$����IQcRGTef��	����DDDD�;Lꈪ̔	� ��C """��X� Q�1Y�rn�%H�0zT[�v;���vumkk+�2.�(�Qm�����:�*��}g�=+��BF� ���5zT[Z[[q�ر��J����ʸ�˸�5J��3��w\3��K"���)������ڊ��8��V�'��˸�[y\�4�<3n}�5+&uD|�6:�0zmgƽ���v��_��r�2.�2n�q��h�̸��̸��� 6�L���u��vA�ŧ�!Bſ@6�@v��2.���(�6ό[�qk�:"��3ro]�U��JG�!�"�V+b��2.��X\�4�<3n}ǭL�$B��w'_��f�}g�=0Z͘T�dY�Ç�q�����q�;n-��:"	@�5#1:n�V̖s�.b�Z񈈈�H_L�&�k���j$v-��]VIs�%Q�`RGdJb�rnܥW�}g�=L興���`� jE��q��U��A�M�,��/�P������ͦ(�CG�����7��O����v�e\�58�Qm�����8?jH~Ťn���Q5�2�eɿz~,\���
���C�����
0*�c�K"<g�x����k2��r!\��汶�q�^��#���Q�cRGdb�����uX�c���k��0)*	��^'�� ��p� ٠Q�1�#�������G�f��DDDD��/w�ҽMDDDDDT�d׌�ͤ���i��@DDDDD&$`ʨ�L�J C="""""2��(��ͤ�˙LPF��������C�q-��+u5��X\��ݡ�DDDDDT�2��72>{啡��ũl�x"""""jd2pq�����1�RW����f�""""��&���L��sq,���ֶ��������Y��=��/+�v��|� ������d��$��αfR���q{���L�������|
 ,A
��=�|�����I
    IEND�B`�PK
     o_�[$7h�!  �!  /   images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     o_�[���� � /   images/bf314729-9196-4b76-b154-4ab11fec66f9.png�PNG

   IHDR  x  �   y1�   	pHYs  �  ��+  ��IDATx���eGu ZU'��b��je@�D�1D���/}�`��؆��������4k�`���<x��a#�ƈX$�H���J�R��n:��f�
�{n|�V����sn�:��کv�r�l�l�<#a��o�l�<Ca��o�l�<Ca�	�;���Gn���O�͛7S�~���n�l~�����q̛�oN����
���:N����Nv�&Yg6��c���LDyF��B����-��,��	���'ֻ��	�Yg�U��x�W\���j���x��8��r�u:1��23���@w���	a#�8&[�l#KKK�Z��:���G�6m!�g����!�J]_dׯ����ݞ�����s�ya��Hw��e�1'�9֞{�u� ��ЗUL�Q�e#���kc���#P�5!�
�C6 N%!��/볨�I@����lD���ӄa��9,c.i��$5'�^���$�	��@u;F�� �/�?-����$F��p}w�'��Z�0��+_��C�^w���>�!� k&����s���o����G�Ւ��r�7Ά�nK�dzOB�c��O��O*B�N}J	u=B!��$�"µT.�k&��꽡@�T1?����q	�HBe��|��aD*��V�+Yf �1�}��|G��2��k���c�摓�'Fί!8�w�8X��0�q^#���~czGd�`]�ۯ��g`c�!Eob�sO�����w���|���������m?����͉������ٛ��ٽ�R��Q_��=�N��A�q��v�8�$I�}�*���8Ү�	���b�A�3D��p.��n�ڊjc܉H�S��i�S���H�+R�'�x���(�x�����g��t�t���OY��0��#�-�Pw?���<������sg��O
����]})ۯ	�y��­��ĉ��'Q���۷|}�����^��w]}�Ս�6o��UW�j�ā�WJ��pl�ȋN�<yF����:��u|P���S�v�H�Z��ȰH��~|K�W�'��wK�Qc�RI�����Q�J���ݖ����XK�����kӤ���7i�8����ܰ�ޞ:s!k��jޱ�-���f��W�s\�رcgA����n��?��O|�S���-oy˒��Wcxh<}ӛ�4}߽?���wC�.l4S��+L?��"qG�&n=,���<�y�ylx����~��LK�\�ez/� O���o �#x-�����I��P@DQ��GѺ���@�?���=^�)�=���s 8�����~���>���Xm�c�~�J�<���W���;�\ j��9L2�O�����ˍ��I�Ϥ�?�9���}j�4���c�`ĝ��Se�]>???}������W_��E���m����ɟ��^�W���e�aʭVG�q��igx&�ɇ���ۀ�A���=�!���,��ʾ�_T�U�H�߀��@���X���o?cii�;��MG��]Y�q�8�:��^�`���p�5��p��:�X��t/����Z��+�zի>�'�-$����[��}�{_y���@mس��`�� w�9�n]�V��ҵ�a�d0�aD��dn�R�mC����~JC~��U�d���9v�T*��8��j���}��}���I�:��ԩS/��l�Pm@���t�u�l�D>[p�_�S} ʍ	����O_F_��y$�t�
�ϒT��_��=�9jS�P��7��~�l�}o[���Pj����2C�K��3��w���'W��܏x2	��LJ^���K2b+�*���T7�<��a�.X�hOYh��摸�A@ڭn-��=�����k�B�֨������ �Ǐ;�������m��j��� �7��@�B��	%���{�#���[��@M��]�F>�|ҝ��A�)�ɸ�<ۯU��n=��*3-�I�J�J5H���������v���D�i��H�eЅWjn����"��߀Shn���GQ�,����|�y��dR��~iyy�¥�ŝ�f�у]���S�+6X�Z�۔� �p�k��"乿����!O�G��*l���	W`7
�_�TR�p2(�n�R
��o�@�y�t���f)��iX��g�y�B�3_�T.�ڂ�}lc�i#i~z�)�0e+�\�3-lw�FU�Ht؅0����+'*����1Ǵ/=.�$PvIm�v�tzB�8��r�reb��G�v���f�l$�����WAYW{�=�ҼOXO�4�3 ^�2Ix:��z�e0��OY$�R�HF�X0� ��Ab	m��|>6���Vw�SFg.]�#<��x������P�<�s�ݱ���j.��l��QB/4��d�V��@�Խ��5 F5����h�[.���V{>�]0n�*���@���_fi䠍�y�^#�:!~Nz��� x_��/|�K�|xT�������tr��A!l#�N5l�%ж�333�wG�Ѹ���@��g'��퀺���~��������k_�y衇�5�\#���w)�:uJ�3����`���u�MX�r�>��2S���Y.��'�!Dq�G�F�A=R�uf�'��C"��-���&�p��D A���J��r��І��>�a�*����J.�2n_�Z��jQ�Ў�D��ԣ�*���#��_�
�eh|hc�]�!v�
�Rf��:����"�}X�=J#��oG����'�:�Ƅ��l��{i����=IP�|�O���X?�Y%\�����C��L��S��%�Y�M�J%*���tNK��N���a�,�p�0v�\�%.Bq���N��i]���!:�j��ҙ���b=�t��~���&Z�<���7�(	ı+�>��*��L��Sg�{[��6R2�V����#qO߅��:��b��1#Tt�$���,�jI�A��a(^ 4�J6/�z|(��"�yF�vx��>��Mp?V����[��������>�<�����p"�4������W^y�я}�c(~�,�(������[���گu�F�^�ϧu��I������b.�b��K����&{{-��o�O_X\#mY��0�+'̳e���~���5�����{�m��s_�73�^^*�� �Q��bá ���$4�H+���
���`1�Y�mp/�|��͛7_�җ��� �����	�=	�D��6`6`0�1�ךg=�7�����
���{�?��G=��V��6��[���8��ۅW���-{���7r)i(�隡]�j�� kKʂ���'y����_�ћo��N�Om<�_�s��痖��}�� �}�^ܦ+��+++��V|�R��b�|z���=��|t��E�'˃��7֏iX�#R���}�<�����vY֗|9��+:1-{�2������b�4[=���>(O�s-��`yX����Ԧ�o�i���x�㦷��_���XƤ�������lP�Є��Ф���J��	LM>m�{4=��?k�'�e�4���ەϗo��vr�j�o����L�k��������jE�~���Q��������� �|+��3�.?��[�}�=�ɮ������8�Z1[j-��б����^�������?`���>����?�������;y>4v3t�l�u�M�@G*(�S�Mޘ�+�\�FS4�x�\��m���h�Q�p-�c;�m��ڕ�	�קж��L�Z�3B5���yU��z�j"ԃxӆZ��9�f�wv�KB]^͂.�s4GA���1�3<����JA�4'<P��
���������h���P�p S�?�nA7v���(a�*����ȩ��L:~����x �ܽZe���$pH�R�L=֋��:���u����r2ܪz�ɧҍ0]��~���J�4�r����S�{�~Of�i<~+ R��Aa|�o���zcyT���9"�j���a�M�O�cH(㸐L߳lli��>�O�n�h��18����wC|����J���,��-[ڢ�i��|�6Q�R87����jj�b�4�7$�L�C|��h�7Cp�N\��Ӧ��o��9i��sU��ǧ-���`���1��:�xC;)�{H��8p�q��_Rvs �(������_t�9G>��O6�ſ���8�����c7���}���m��؏�ZRe��tCZ����C	�9�������ceH8U�s��چ�^�W|�W~�W���B���L���������]PvmI�����@�	vg�M�u���CI:꣺"ͪ=>'�7�v�\�	��H�qr"Ӑ��j=#̫80|0$��â�S��D���(��-ևx2��;��P<�nl~,ȧ���4����f��b�J�:2
�׭rK��MI6�fqq,? ���,T�8(�t6��.��E��-N�������R��"`�'M7�EuS�oU��l�>�^T��~#%�!�1���ƬDb���si��Z��c�'�߹��}�I��<���s�w�9�� �W��m�{;�E��<���s�l�T8ı��y���U�~p��D'	L�"�|����m��5��}[�K����,:q�ʵp��-��˴��`�֏�1i��v�)M�p�����|�]?��7��6BN�T��O��c���C�=���@u)����5��>{B�#��"���yf�þ��l�A�9����K��ɾ}�J�^{��`��Pw�;. P�a�D�C�q@�q��m��Һcҭ�XS�u��wQC��=���ȼ�`��fS)��ϋu��l���U�ly���u�yO%�Jby8Q��C?������@��q��
���q�����f�*+�<�a5�Xk���s�f�[�w`���͝�f���9v���Q`��֍!?�A�Z�q�VP�20P���sA�m��w�܅ʁ.> B���~�]F�������6�g$%�[��Vb����E�:���/��%(�W���{É'�o`{a�� ����#1?�l�� �=��ը�45��������'q�Xaj��B��x,R�Wq�Y1?Z���xz������
KP�x�8���d�������u���<~�}f��+�y���nc� X���d���ݵ�s: �NˤV�>$�vN��h8�H�@����l�>SYYY�ܯ����]3ܟ��L��;��_����mG�_5!`좋.9��x�_Zo�?.�=	�U������}�c�9r�� ߳�Ν����݀؀x:�6�) �/K���T��\��Y9�y��m�Š%n�ߞ%�C����瞑�{(��5+2������4r��/��{n��������Б�mOMU�qT�'��2�px��6����!�^�;Y/�Z��Ux�����o���\s���%H<|g�#K'7�؅�Q��$�����w�uɦ7��3J�ҋA��Z��������؀؀�X��5���R��~� ��{/x��-��?z���8�l�Тǩ�?�
v_�w��$���/�����|�|�#�n��ƽ����9�Y>�ώ���L��!�������s����o�#ʇ>���[n�s������N�y�ZCJ��0�����l�J+�v�z`߾}������M�r������tW!�h���L�_�k��sY^XX�B0�z:��,o~�=���f?�(�׺���q�hF�oݺ����Z���+�_��_o�۳��+�â�ݘu���a�p��OE��&����ŧ�*,�:��sܜ���1���j�Қy�w�	{r�^4�l�f�J�h�jM�^��R�i����I]�
�����ٵOąո>]�х0uzkƈ��{i4ȞA�o�)�#^��&���+'~����<���ؐ�|��a��p1q�7v���u=��<��7�W�$�����㹔m>���&떾듣�h�	;��c�+��
,\(�!H�^E%�ٴ>��MA���̟��z��8Չڳ�eq�A%q���`�I�@&�?�VW<�J�����4I�!�p�Kp� wq�U��e����b��.��D,Bsm�{
�#l���zW����υ
(�`���c�g����ףO�������]�,q��&w���g��q���wא����{IL(��	��Ku~5�+Q�4q��cY�1t��}w#��ru^�o��L�/u��X����z�z6��NĄ䉎T�"7I�HQi;�3�y�E��d $%P:K^��C�x|�qWܡ���e��#�g>�H��i)]�+��᩠�1Ȯ������d�.����n�| ��#$f�.Dw��U]��ꯓ́��h(�_��&����(m�G����jE��
�g��$	i$v�%wi}Za�#=�sJ����$J'��%b.D:�+�Kѝ�� ���}��S��ab�P�a=&.�7�R��	�Iߚ��cJe,��2��S*�<}ǟ�O+��K<��8�c;(ɢ�=-q���]�C%�;*l��*��l�' )�aI���G�l;"����^髂��hr�����i���A{�����h^:�Y��`�h���T��"6i8cV�C�
�MAJ회]�>��	i}qc��H�
/�9t{�.�8�r�]�Vj3N���t��~�.|fO]B� rP�ԦX4"ZA�ɺvї����qfq��w&�+P(���t082�x/LL��mW�=�wϞ=z�0C��j4��Cs�<�V�VoB�]xy���J;X�s�O8�>I�t�rd����u�aÐ>�j;[�5_�cN�K�yb����홑�����vE�C�]H�]�O����]mnqrIx��ƙ�헱y��k2	ᮐ����R*�ۡt½�O��U�qٻ*�ql��C^�֓Us�|U��m��J��'<F�앴��)��ca�oj�[t�$LK&�g�O,H҇!����S��&�>c,O�e.-����%�U��ԏ� ���I�=c�>��c��5ƺ���&�(0�ɯ�ی�֋j���gԫ1ь5�FxI��Ә«D.v��"��u{�d�^Yo�N��ʢ���x�F,��a�l� rU�a�J�ѐ�y��L��<��O歂��� �/ޚ�����5���a	����@��%�H�}�Z��ޓ{�"�<��ܭ�P�'?F��Bb�J5%�������tz�h���J��?ƘS���v��z��X4�i�H��d�*�2U�H�5'�&���S��恧��0h0��&$5�g��PxǕ^��'l�rq7�5��R�jAv�	�2��Oj���ϭ�D�r9�V�E�-q�r�,N@]�u�|�]�L-Q0z�q������6-�u�L�v�g�ړ2,��+�#w$]ow�`kV�יY4q����
��Z��D���M�~�߅8�����S]���t�s[�B�����x�룿(:�'D:�G�����F��!�Oq��~f*&��p��0\�扖��yn���ES�=`�`��cw�-Y��b�Ԥ�(d�	M J���ۘS�N��j���5�D3e���p�#gRH�l���Z!r�G7����_�z������R�*�)R���]�a���C.=_�U(fF���C0HE�g�u��Jh`�Gҵ����U�T3��v�q˳�Ί�Z��f=���r�s:�=�Z�^,L���+�+�W9E��rp������L� *���M:x����)������@�Q0:��(9NY��B�X�9?m�n8t�D8�$""��^m��8��1�D�3�3�0}M�B��Ƃk<��� �;f��u9�Sh�Z��B����)�.�f�Z�Ŀ5�u�7��8�u{�J� ��몀ǁ�v��{�'��%<��m�M''lw�F�f�x�D1����L�6	ꇁc���l]�:1Tu�A�G9�(S&�RG�IMG��AH�����(ЀT���՚�r��-��a�f$7��O��w�k�:j�P����E�%i.�&�-��|��w�D!��53Z��u����xH2RD�qC�C�\��D�:⑼�L벹�+�����L4^yZ��Ig��R�[�#X}�9�� �'�$��i�a+�LRuUM�mc�I��\���x�u�Vyا��CY�-T�my��\X�z����3J�]�F�$k .��4�%!j���~�)G�r�R5v�9�6E����s+1?s!�;����0����5k5D�	������&��+�g�p��.�95R�1��,��dz����{�V���mI��?�!�3G��|���M:0��9u<�IN�ܘ����i�z MhLJ9�� �%^Đ�!����vN�s�F�{�(I(8��cH���Pq�{U?�����x��- g��"��~�`q�ұ����ڵx�೼`��ˇy����8j!/R+�]�qȌ�&H��+%�'�����v��"V�#�k�|Z���X�KJn,� NĴ� �SO�K�WԝI�W�uL�_x��#�J%����7���*݅z$sus$����zLy
��<hZ�t �\N�ڜ�8t@��+��ҵ������>j��vsg�}�҅C��,����%	�����Li�=X��X5F`#&��ߴ����샒�-�I0��b�eY��8�j���o(B?�WW�7e1�ށ�����߃��r�*��kx�!��\����NS��f�k��\8�,�Y��=��"� y�G�4TR} d�=m){w����u��e�Q��^�.v���C� 
�7���b$��[+��:�D��t
�^�]��L)p��	�����X���c*b#�h�p�=���2�Z���^��������+ ��u�X�:c��a"������GI����1���R���H��e���f�����0R�g����w�"����'���IR�Z���w�q�s�Lﾩ4��`��1g�.�~�X�w#�fK�
�����h�M1�T� ~ُ��n5N^��.�G^+b1��C�ne�q=����ឲR,EG9�������Ȋ�Ĥ㵁���%VH��;M�/#��pZ���J%I�4f���;E�8�r]���c`|l�HDB��L'�W[��<,�s�o������z((W���b@L] �����7�� �&�2���ν�R�z�M���o��_n7OtX�M3?p��2�5���#��J�:�ë�.���v�;e����ca#jn�ߠ��	��Ͷ.�#�0��-�<%��g�?�#�0�h� �P^]��1u��,�'x��,A�x�%�8M�B��
_��1r��O�ѱ�+�-�������sI{�c���k��Ȃ(P|����3���FP���׿�����׼�E�[����de�4�����#��>x��o?7G�������։�W&퓻�*��5�"�c�3�Qլ:dy{ɻ}w���;+�vy�O��)������,Q���HD�6�`�`�$�T�S҆/ޡ�}���e��HhGA��s��t9j�	(��%�͕� �J��^��&� ��,�0��WE�B㣶c1�X�~7Q���{`� Nǁ��Y�ntdYT�=ɖ�u����?�/� jB��.��y�_U�P��k�F�hXjc^#�^qcS���B�1���[���-{��g�/~�O��;��3��=�v�W<�����D�^y���t�4 v�;@0�Y�V��4|^![7�!PSO�%̉A �јL�yV�� ܲ�,��uK��� 
g�$�1鴥L�Āք�B�D.�!h���lJ@Xe>H� ��V��b�T;��#���,�� ��d�yr��,޼��~d�S�V�:'����%	�~ϗ�D�� �#Sg]��m�]v���������Ǧ.���;��7AB+���"����V@	�ȃ� :�8 -�S2`x
/��:ٚC���E{��hN�o��(Q�s�g�T��'���j�č�� Ϡ~�L)+���Z:a���He-�%@^��w�����e5��+A{����T W���	צВ�4B^;��������_MO�����߉��$Ѳ�I*�j;��,Uc�D��s�Ww������gw�G[�����Sr0+?�e�JL��$l�B�O݀$Ǚ�pA3��	%XB�9�I��A�� %<��6۲R-I��4���}�r�s���w,=|�}'��;I��9Bv@�i��ق�D���Ͻ����ߜ3[tO�z�.�t��縄{%ޚ�h�d$���$ B1(�0������D�Y�YF�	���@���{_-��3�n	1+$�.��)8�#5U	c�T�is�eǔ���A����������GO�s����M.�'�+�1��G�8����Q�kf$21������b��`$�cN�nY�Oz�v�t�9�|t��Ϻ{z��Wәs~�TX~I��hP&��H�PaU��Ip���D�m��:L�%��bӳt�촞iw����e�l�Z��^��DJۥ��h��{�b�\�z�Y���+�+��G�S��(����v�1��9Mg�ޯm�z��ӳ�s;/~G���y�:��I��!`�S��&ԔM{]5�����A����ΈH�e�Q� 4[2ci�����t�d��8��7˘]�d�C���H�{�~��V�qIL���������Ն+�~����!�����ک�F��ش��on�������m=�e���oqj[��q+S�|�wѠ�$�p�Z�mˑ)�E�!^%�(��א����>���+w��%�T>$�����e��Jӫ�D/���*�}�xU�U��\鬐Ʈ;�J���!�t��ڔ�M{O���w����N���<���[y���2
K$OH��+����~p���?����=S�_�	ۿ;�r�Boeٍ�Ir�WA�I@Ĉ��h��	�	�JA���q'��!�]_ܱv��V�O���rO]���d��Q��J�_��bY�+���,�����IR��K�J�O���l��g�y�<ԉ�B��;,�k 2��.�s�χf�	�>���|�h�8��b{�_>���IR7��fw|��+^���������xꥋa�{f�&P� �^_J�E�H_V��[����KV��&r�U~�q��޷?����ؿL�6�c%������^�~���G�en���+��-���|p�J�{lv���o;���s��"�w/�ٖ�!Lf�Lb���:p[�z~h��mYvS&�b1ץ~iž���J�p&�|�s%C\�S_��
�11�͘t�3���o'3'��M�t�'��S�����-����[o⹒զ+Mo����/��󊤼�y���ǖ]r���*�	(h��@Z�=Qb��BO*�	%�p�w�+�Pc��q�GR���V���
W��X���6�{Ƞm�����XY�a�5c�Z�M$x�<G�fs�kϙ�t���(�?���y�w���#�l�;g�ʑ���H筩r��_�Tq�7�����g�Hi�MJ�o4T.����s�Q~U���@�^�*�9�C��@7�� Ф��E���+PSL����W����\D1�o�)Mt��4h9:f|���|�-o�>kv���)��M�=�����]�.-^��|���(X�)�bg��ɺ�h(� �+��lv	�
E���3v�:�˿����>}�Im۳N�"�[)��0j2� ����J��d��� ̱��}�O��<_ز��$���T�� ����jy�����7�3�|�/���o|����Ti-m��~]��3u�{���tf�T�מߡ��P���ȱ�$�<�\-,)?iV�i ��*|3a=x�yN),��e�/7��qh6� \*-JSU��l�H��Zy��~ij�/����~�����+՛Qk9��������j큟���?<ј��Vw�M�۞��2%�Lj��KH����V��D���Є�M,��@��5��"�;�þ��_��sM@���Uw+��g�y�	�吔� �W�l����?�y�s���黿���<��,H���Z�~M��_�u�ܻk���U˯��삸��D�X̉�0�H�+��q��7}A�J��I]��Hv�߀-�^-���ȕ�����ک�a*��[��V"i-��,
%���o� ����>������;�w���݇�.�,�ܤ�$��5;���49�Ǚ�n�w�;�@�?�����(J��(!�}&&����Nח+��T�J��S=k%���`�D	md���告!�H�����9�0��{^\v
DƸ���g���O��}��R� ��,�ĸX*Uݠvƥ�?�r��[�*w��DY�df���GB�r���'�թ���yg�Uv:�Q_u.��c���Jt&v�'�-�u1Ƭ����jZ��*�#���/�H|.�$p�7��&���I�dC!�HAb�d��2	��D�2Ss��6��e�|����E����b}n8;��@'���ڎ5���V�
�K�S љ�2wV�>j��gڣeR�g�/���k���S3�I�W�5L{�g�<�}c"�X1��멓���49|j�2̾��������wK���w�&�R1b�%��+�V�#+3�W�Qq9�<宀>�x$�uʵ�̄�iH�ٲ�
�gD��_���KrX(�Ahc!K��8����Z�"CD���;�t�;kM�\��n�]�ԩ�س��Je	��%jɹ)�Q�H��M4j�KA[-Bns,S�DG���	ʓ�Mw�8�?��;�8u���+)�I��eo�f�x&hT�0;xB�7�옉�&��(#�2Q�n�UwР]\���q�3�)C��Mj�*Ni
��4�j�Y4͸
�DᑚmQ�$9�t�nx���ĝ�2��΀�I0��U`p�ԯ��(hu��s`\Qv[����	�u����h�v�C;�X�$�+/?���؝�1�սJ�ՆO��Q��Rf�"�[�6;�q�����A�M?� u$��cھ+i&e���t:1�3�Ru�M�_��3�?߶���F��׬F�uD9O\ѡ�ྋ������8~r&�m#��x5})�a��!l���tH�z���A��A���E�M4M��=��q��p{�ظՎ�w��qw�9l�y�q�)��uaJU�b����5�����'�[xz%����5z��j��K�Y�e��v�.ou��t9~��I`	.�삇��EP3�l�$��� Q���l��o^P�b'��)� 
�a���ӡ�B�F��K2��U.�@�B��T�)��3_yt�`�3t��>�'���F6�p�,���v�̠r�W���3�+�������[��N�*�`T��]W�+�b��fԛ]��%i��0��x�M��N�x���z=-*O
���Am������2�B�	3Lq����N���{�O,*�m�iV���%Ɔ���P�w]s�ZDd�vѮ�Z�LjEI�Y�Xy�WmwW���6�k/]|&��#Ǆ�@�e;R�k�AruM~e�HɈe�]pl�@�JAP����?��&44�1���������S�y��*����Y �݃IE
��s(Q���D��U���B�Xt���&�@4(Z[��9M�=�@g��Q_��A�#����7���ȾB����>��=g���s�RB������˞ ��B���5������r���7h�Y�[m��u�u���_���F�Q��I/qV�%R�n�*�K:g�$����[���iI�_��b�a�p$@%�'"L�]����5��4;�N���#O(��S�'���:�]�-W+&Z���U\�O��F���ߧ�w��0�v��T��{�j�+h���m��ʲ5��g-�M���AWB�](�*���EɽǦᚅY��f������8�����k%,(n��3�;8U
99M`O�[�#��ٺ��;7��dqz��4fJJ��3NY���֫�E��8R����j--���̞7��L�H.��Q��i׳��+8�u�?q�&*��K��ȹ���''���&����!�9�@���6��H�=w/9��;�	��8j�����)L�p�*�G.�)O���oG���%𲀿ޯ�1�Q�˯r!�<iG����,��.����Ui�l��	���͸��q�I�;c{�0)�E�A����HqQ�f���6����҈Dly�>���m�&��8���)k�ɦ�]���;ϲ�$jm��"��0в]���&%뚼B�s����0��ì~䜁|���������?K�F@H�"ؤ��F��ļPEbV�x�$��Ψ�������z��$Q6s��_F놮���8e�)���T�90%U�C��ri7j	L�ͼ�
��Z�%ƃ��P����<a�֖�U��Z���e�W�*�u���ZѽI���YJs\B���v՞�5�~3�l�EPD�Z�]�	x��]sB�"_,wr#�r�D}0�d�'z�z�X�%�aJ��'"er��`{o��Цh�&EL� >�����`iZ�Dנ�S�"��u���t���nO���o:�dI���.����.W���D�RMz�3oB�^5٤��H4j!˼g�i�+�^B����#�@t�Q�?��!��~yq5lX;�eՄT��úe��/�C�3��;ه�6��/�:�*�@ #���Z�I=�8�	cє��\b��p�����!���$�
k�,~>-�+����ha�ELM)[.]����V=��������;�'ݻs�b��D\&ڛ�C�=���[A��~Z[��^X���P�DM1ѝ�ϫ�7i(�2S^'�6h�w�C�S�T<��|���S�!>�H�A�Z.�%xQX�x��1�(X\nʤҴޮ3奀��5(�}���"F@��oB2��K��
M����.M%u��w������" 	�(&3���M�2�GW������ے�a
����^�cSƾa���e�j&Tlb��|qP{�����͆ �ِڭ�n�kv��<����7"%_#!q:��6AU%�������e����*�sj�!�=���p�Z�ZYrh��̊��# !��h�Ĉ�Do#K\,����]����BQr���
�MS�HT^���'�����qx.wF����x��M�����jw��u4�ZNl�7~�c�
98/����Ñ�5*u�Y3�n&�&�6��v�{:/~�V������"�-�eQs� �4��D3�t��2��l`�D�qr�:hW�@5#��]/e���sD����*�Ձ��L�5W̹ H�q,c(�jC��R�M��"�M�Gŕ�����g��5�͸m�A��]����JL��]����;ٻH����4�ki�O�6���f�t���*,31�dH�q3�/l������z�D�Ԗ3at�b�N<�њ�Txf��a{��z�HW�	�^�V@�Ç�T%���NH�J��$���<�\ו3[2Ĺt��)l@p6]�&��%�� ��c�A6���E-��M@o��46x��MN/�M����w�]�nC�����W'ϐ�Ҋ��t�_t�#m)��.m�E�RU�WmH�X��D@2���9�Mx"�m%�F;�NFcA�����܇�Y3�"�ы�nB��8�`���
C-u��z��o=�@X'%J�YEeO�Km`
f��4�.;�T�h�Aٶ磍j4|>~r���:Ep�o6@�v��>|+��LT%�&Ƹ7'сzr$	��^U�em҄���mRoSL���A�NQw0�!��&4��8a(^����0MFj��#
 o�H�%�?XP�$ی�-���0V��c=GrY��Za��]��r����e �ӕ�$i5�I���L�ߖ��mCXU��]|������K��:��[�[O	��C��	9�§ϔ��s���G�i��-����	�+F
d�$@��[R�R(n�F����i�al��n�U0��<4a��'g��_Y�P���u��*�"u��$(� =�ݛ�)��$)�����q��F��@�@\EU
�ч	�:	I�OPʳgJ����kW�9ax���<E�\�
��D�m��~�*�K��yΜ���~��z�p)�u��S�~����s�40ӆvӹ�0!u��YRR�4sd��(	I�A����G�P��&+��oÄ��w)��;f�h,J/�h��������9��d��hB*�"�7sb��|���N�P*%�����6�a���'zq8IE��y����O�ax=\��]W?�a`��l�'R�Q_Y*w5u]/6X�����4"�2F��I��jG<����1LB/�{��=���A��k�v� ����}��R6��>t��X&1�an��n�[��VA�I@r���C՚&��ӎ�m��&h�S~��K��)ǰ�N�-�k�8&�c�m���5ȴ��؏�0�XF8��RiE��yn �(�7�9���)k�)nY��T�AS"��\M�a>�!W�)��J�".�y��5�W�k1�0�멎�E=Q� �MO�0�)N�ٸ�m��{ͧ��6�I4�h�k��N����
W9�/��l(��s�W�w	�#�1p��Iɦ=g���?ڎ��Ch�h���%c��#��j���]N� �?��8�H�F��_9�\\�$�jQI,�m9��6�2I�iw���":2Sʂy�;��n'!�+H��Q�	��%}?~�����5��Q�``�"�������=�\��������N�A< T���!���%�?8���z�߇����4��Z�N�3q��6u���D�@�,e.yЇ=g�N���J�:�	�����/~��!�;ʙUR<�	T/��K��nh������hK���j,""H�.n�RY���R�9Œ��t�6}Wyݻ)k��3-�/���s���m�1�-��*���$=��zt��5�l4�ä��h�Q�
N��O�c��@ �����͵SOs�w�q�Lv��J��F��_'��T'SYgI>��x�%�*�al��zntꕒ�H>>�vap�]0�!��c��<�W����uDx���Wc��K�mE�0�^�\hx��C���#��"��N� ��j�S�����G���c+�+!���g�]�PHļS�y����C���-Y�}��z4p:�ڎ�%TϞr��,4[���:���&?{����X�B�T#(<0f��y����ط�P�bѨ5�׽�]��ۿ���J��V5*�	���e��Augx��F�� *e4q�?��葄/��27���ҩ�e�\(KD$�r�:�7�nD�S+�+���s�Z����d`�8f֝�X� �k���JS�h�|��S�!p:	���,�U�t���J�x(��w�r�M����k���k��οwۆ�?�Ձ7�F�d]i��DO���wm-@�z��ס#1���g�D�HZ��8X�;4X�7�p�.�p�輠OF+��I�����ϖ?�ƷV�
đ��������b�$ ߅��H��Kj��>��/
FL0IR����|�y�h�0�p���r��2��8i�~��n�zeRY�Ҷ3g��|��޾ݓ���2�媫����3H��d�i���7r'�����<>/��[�+�;hD�?s%&4��Й�� ��0$3��)�	{�z����s	�K.H�s�P�`ؕ^���Ýen�m�.��
�,nvҺ�0�H�lvF���7��d��H�/�����眳e�UoD����oX�`<���T�����_n/�F)^"c��K�ERs@�(�N^n��O��jA�h��`YVS6x@�wj�A�a������J׹g�71|O�xw��꛾��[����׻?���XwE��"
g<�-��(��^�>�gO)kg���v�w} 5��m��-�Rq��\ߔ��2�}��4$D���(E˫
6�8�MR�ɂZM��us)��ֺ,�&���ib�)�F�@\0/� �i����?j���>���'����JRsv,v���:�0D!�����j O蕉��&��$1xu�C�kq���#d�a�Ϝ\�Q��s�a���a�Q�a�B���J�>ϴ��;�l�O�_X9����k�]�{��6��8�O5Nl�yѩ
'��%oe�]�w�%��߽����#=�X���;I�&	�(3m �DԢ"��(��M�&�<���\�C��MR	|��|��m �&ʙ!�O�Q�Q8�y�vB�4�ʤz&͑|��%�+���1b}�H�Z�ݠJ�߀��{eI�z��a�x������f���;/Mn��;����g*����&9U&�Z�4���[ë�G?���ny�'�x�s���sf]�s�sH�0`�s�d��u(B�e2Gxi�r{R��ʥ��?�=��L�>�A�8X2���LP�%O����J�쉔��x4ญ����������*�{�!z�B^uU��_�=�s�����g�f����j �t$2��=���؇l�����%&D�( 2s:��·{'\�z1�}F����2+Nl�W\y��2fqO�ݛ+z��
��G[K���cf�w�3��]�R���Ss�0�D+$�z �9J��w��Z��W�L�k�b�~����|�l��4	h��2��U�}��v}�����v�s�x�O~"�]9�5C d�z�pT�_6��WgSkq,�aȂ��M�-ip��l�^�oey�?m=��{.��ȷ��N<z|o�D/c���Re��|��J��-_9����z���&^z)9�G74�g���,��ߡ�?KR�v����ȣC�������X\8��sR*9d�2M�V"��������M\M1E�{'�	=�J��'����:)�cJ�K�����t��ʁ�a܉O}����_h�{�t��[�\⺵=A�u/��X��x�^y,����G����+w �<N�=����yy�m�-mn���mA���c%�Ijm��w�v`j�M�A{�w{��kx��\OpAy�Wm��Qx�5P��!V��FHg�!&�8�!x+�ܟn��Gν���旿\Qp��������mz�u��w`�ܠ
��[N0���k<!7�96o"`�UP���
:��
����Efќ�Uښ'\MF��*�d	��QR6Ś�6e�S�����s��d��\��ǏEg~o���AևP�p�qQ�^�̅!%�V�za�l�"=w��.R�K��p!�*�(���2�%�vx-��L�P4�y��c��<�8o�MD�]�g���9r�5�w���%���;��b��+��<��zT�ɡ��������Kw�k�����@��|�q�2�g�.]��!��� ���@�+�-j�+L�f'&�!���8���$	���I̓ �K�{��i+z��v�`f����.0�q]��P��Ven�v_�7��7���E��_BX�u'd[�J���FTg{KS�o��-���_����P����.�?~c���ωN�%z�POy2�W������N�<.�p�r'�xbm�t&'��v?�j/Q�Wk��o�"�4��<?	�z�wrf����}���|��n�;����׿���o�e�/}���詟PA���hNM�˄4����N(�Dz/�b�)�`Ɖ������1��PO�L�tE.\0�C�R�P0�M���M'���K}���&ʍ8�V�T���ݹ/aџ����O�U��5���M_P-��U�ow�;K�E��:�Cd)��I�m|P��]��Q��1��fƑ�ʹ"�s� ���x���t{R��Y���)7��Ӈۿ_�г�,=�/U_�����P�[^��T�oxfA�gS��-���#_x��}o8�Ⱦ�����t:�e�LK����+� �	1�;κۚ�����R��(n��cc��y�= U��Ro~��J�m?R�,�\VͳH���jS��[�b�R�����JRYh���$
*d�֟
i5�-��E$�oy��c�]/�7�E��:�P=���H���N1�n��P���m��M�����aܬL5 �;�6S��*z$��^��Q�����⩲�h�	w'�h����L�`�cG��_p�x�C���ۯv��_������L�=���U�W�0775�z�6�`dDK��>��$�:�Ϳ�����|��b)�} ���i6-u�Ym��~��P���{�#�^�I�L�
D|�uo�:��o���\z-Ϳ�����Wݟ���ջ��N$(Jeh�k6���\���ތ��L�Q^4��R)�X"ҭ?G�q���w��Ҿ�AI�Bﺴ�il�:N�>�)̽i�0{��b�;���g�9߹҉�)KaⱲ["A��L,�;�Nq��R�U�7m}~�>��9��NBW���t]�JcV�1!��Iz}m�$�b�4�C�/xPEq�;�&0����+?����a��"Ѱ+W?�,XZmf��c��3 _�{���m�"@��/�ЩZ]mCCH�����8���C������Am?���D!u��q�S��2 8t�0=o�~�p�z\��G�<��|_pr�۳[����<�Y!�)q�4_����_�3��}b���zP��e.L�fg�������{�k��P�|r�nǚ|E:=d�����&n�I_����q�I��6��	�G�c}.�b� ��O�k��_�EVbԸ|���Qfb��m�b,<�T���5�i���_���W�+Y���!�0Pd��(���oM�1��<�O�����z�'Zt�!0�yK���n��21�EFAO��
�e�	X���U��K/ѻ]�ZVm�ur`ia�ys�V,睗��[����!���h�[�_'���1u�3� ��FB��\f딶�܃��t�a�E����2H��a{E1�`��Ct
��o��T�E���$�qHb�\����U����0�6̷2�Sa����?/��RG�(��၀����7�2�^��6L�v�8�Vw�����^�I�D��P��U�WCa`8�:[O���&���G�b�҈��[�y\~��-��cK�]�i"�y������������bM��r=����]dD{�z��4�m�0o�և�#����k[��P��}�y�u��0��Q��m�fX�5 <.N�o���/I�y�h�}�C��m�bϡ�K�+�6u 5P*d2lj�m��kĈk�+�F�`X\��c�0�#m�}��Z���:�UҶ�T��'v<�n0�,U�����Y� -�!i�b��5Rg^�p�f����KN�4Q�wl�=���C蓼B����������p2�;j��s.y�:���l4
���a���V2c�݋��"��?�y}d.�6��fDv����B��@�f�Jd�ف�������J@��@�m��%�Cׯ���{��l.�q0U�e���E!S���#g�0����Y68%s�LM4}^��Nq��5B��i�5s2��]�T��3�Q������(w���ge�go�^�-�(�֢���y�Cﺃ��?ւ��'*o
O�({]3�3뻰��1l?����cܱl�k��*r�A�O�G˴ E0e/�Zn6IEz,(W^�X�Jb���E�;-H~�Vj���N`�6�F3!xbz��B��bhA��v�W�M�\�g�Cq��Z�"�I�-�R�E���܄��f�� a�0&5 N	H?�OU�)�8C�� �j�ѸAΪ;�����o�R�
�ڀڣ�Nd�q��ԑ��4�q���0Ȓg�_�Y��$s̥(;���F!d�R*ƢQޅ��}ya�.��$��i`���^7�|rb%!�JM�㋋mR��i�R��Z) �VB��Ou@��ΗX%��/�(�(A��9��b<�
�>s���q�T02o���j���rYn��.��8GD:	�PF�R�܌��WM��j�9�ǜĴ��H��� |y!I���S��狭�TED/�;�
�~�Ԧ��h��o߉c�������1����\Q	�����N��.��o�C��u�OH�t��\�.�c���n��-���0��9�����z����M�������or%�Gy����5���FN-I�ǙRh��%�����4t�me,Z�-�OZS^�Ȫ�: U�r���~0��k�_�ae./B��P�å dB�Է�X���[JE��ō�42�Ȝ^dO
b2c�*�k"�f�6�����ʛ�"'�@�=��2>��	���L������I�Z��)�)�N�������#�C4��x��-0(Ւ�֩6���/��{�����[s�b*�$"�ѩ��kNn�c_!U��h��2�b� ���Z�\��V��a�ee��hW13��h�x[�p��Z��m?Z�{:�͜���*�w�HP4�p�p���t�6�qՍ�A6x#�	�6�փ�ض�D&I�t��3�k7��'�����t$d� 񍳹@�"�eJ�Ҥ�xν�>����/�o����w1������ӳ���s�>v����	�_�<w�ѣ8(����8���K�1����:X�r+���T�%�K*�����H�➓ǷCQ2p�+�3Z�M�ŉl�Ԙ(���c%[y�\<u��(Ԇ(�k�ȩh�r�	K�%:��,�#��U9CM֖;��q5_��0b���"�uQ��=�!�P�X:�Lת�[-�0����ͥ
Y�m2Ub�Ƥq s���;{!T�m��}�/*�rȷ� �*�4�������{������]W��ɒ��aҞ�Eh��d?^c��m��2+�懬�w��<Z�*�J\��Ԇ Bmb�v�VA�p]y��ؾe���]F��,���t�ԛ}pE��H@�x\@8l��c�e���:�������9o�+!���3Cb�EPF��3c��oYP�p	½3w�� �d�5+�zf��W�p��
�H���-[.��_�P^�����O6��ݴc۫�+��d�e�SFXr�A-�J�z{�Յ0N��@�#'�+Q��;(%e�	<���jǉ]c�Im�6�@���&�D�ˉ��E3*$K��~Z_˲L>�K��u[i�V�P��c`���!�a쩣��ǆ�_ڞjq��-���^(��"�tPӻA�y�!7^�����<��I�~�ę1�_9�4�>B�q�ML���0[�bT�%�1�vH��o|Q�W�TH� C��4E�
^8�\���~�V�rY�'�e�j}�l�ԧ-iF�vvE_����K�L���K�;m�z.�1�w"ٹY6���o�Ԧ����r曷$/Xh���+e2�,`�m�LiLD�B����V��E�	rXv�w�N)�kc)�����uDB�"��g4���6o��Ȼ�����3~��~����Pڎ:�\j�Ci�շ�ඟ^v��|p�k~�������WBI�1|��ۇf�i����и�8���0�"�a�_�F'tH�	:ԟ�巩��^�w��1�A��b�TI�hB�Z1YVc���+�TIG�O�	O���(͍SK�G�m��e�_��,F���B�X�2�/�SrA5����5Pͧ=	������f�>?y�ܾԊ�������|e�b���Z�2=����y�!����K�mN^��u�+�'d�
�� l)��Qg�ݟ@��@�X�e����l��\A��QA�@u�j<k�V�_���P�x������ց����;w�Oݕ<J���&g>xh�F���eR��x��&�D�[�j��K��p�^�l뎭;���2��4U�V[�*��ҝIMN�[w�FZ29��y��7}�(�������3�l�(/���61и�͕�������>���C��fY/c�8��x�{�ے�LpG�����|9gB�I&�L����-`���)�U�]ZK���ի�H۵��ҶL�B-���%P"ʠ�/!�Lrz/3��7�ӝ�ѱwD���s��/�ʎ���{��ĉ��������}�����7��/l˘h^��u�����ط���<k;����XB��']�LT�1�M#y�J^I
��ɱH6�`��:ϓڶ�����f̖l"�df�o��'�Fg&d�1�(��N�`\RӌB_�FIH�v��Y���a���&�5�8�ƱS�O��F�Er������?���}��H��_���p�K	W��g>���JjΧJ��|�yf;��n簪뱒4��z��VWfy
s%5�XxX�[�p���-�G�P�BCM��LV#��P(�# TF�$���ev����_��z"��2�������?�S���ޭ�.��ou_>(��\~�n�IE�rE�04),=%����x`����|�(�$bE�\t�9��N���J��0�ų�J#�i�I���\;CxU����U/��調>8}0��_[����a�<�v�57�����p��������%q!�ٚg�M��,8h��+.)��.�\1?�U�T[���ھ����vd�)������k�|h$��!�l�<z��`b*�ORG�[_��Z�Rj�;��l�=�a�h�	t���ڐ+<����m22�����	9�F#qh3z�g�_9�	����.��j�����>gPB��b��=N��)9o�;wX����,+u��62�FC��@68?��8Ip�|��`Lo������D�6�7��J���4����u?��� ���c�#��SR��^ȣ��~��T��n^��<�s�M/*P��"�C���dx��9�s�\A���ݶ@�f��"��j�1���@�G����d��K��}�]uÓdQ����hT�;���C�c�,�݅�U�l�eW���K�'�aw�u�C��y�w�����w=�^�k��:�������T�+"��A�;�MF�!	ڃ*��./�z+�0CH����8��r�^�Z�	�_���G�X ���yFzז�R3`��X�6�\I�d����>��VB���3g�P�i'+~+��Q���q�F��9]8^��õF,� ��	��N��s�y�ÿ����_|Uv��?o�R�׿v���>2�1�(�����nos�0~-�Bi'Z���I��.���	�d���v7D?���I�)�A���xo�}�|���z~	�>��8L^��'F��"{�0�ڭk�_�£�q��n���>y�5��K���ko]�&og�ڧ��9����T�6x�|2�^n��I�g�@�j�1���y������q _����G�u%ϟ~ts3�[[t�`5��=`�k�M/|�_����9:s�g��<�)��k��w5����80�&0��+Ӭ�h�mK�Η���e>hSDD�Nʽ�� ��^Vb�)�zRԮ�^�U@m�"x.7�Z�)ʐ� $I���Y�h��,��uB�Q.1~�âqnr��NV���	)����c�8�Nz���V��f����|�����M��ϸ����XI�tYd�B��a���o����}\@)�����қh7�!�J�fY��R;�n���[��m�i;^Sϡ~�(➫	zdO�%ڌ� {�
[1Y�v@%'�$WZ;��d���v原v�O�����{+��wM����B��b�ߖ{�c����,`+Y^����K�|?<q�ƛ����N<n<��'�3wߓ�Od���%�� /��Ccs���ѯ���e�$|��ݘ ��� x,�j�R���dBO�e�Ib�:�G�}3��������yN���=o��u�G��g��⭓B����d&��z꭯��'�������G:-�@��cP�~>�Pz���a�SH�2��i�\�ޚe)I��lL_�2�(�#U������tu^�:UtU�e�*��ѹ�9��3�$�yK�N�3fb�-c���V豢-���E���RqS��g�14Bs�$���@��ΰP��Mh`I�����q��odQ�k���W�M���)d��=�N<QcY��@c���3Ғ�zE��X(�g�n��v�g�-H����԰��P�Z�}%3�U�-� ������s��W?^�k�/�W^8R]��W������х�:6>O\��/c�mKQ3L3^D��D�>7�,-��w~�q4�ی$�Ԡ���IRQv��}$�%�8�
η.�YQ�k(�\]:�:8�L�ɕ�ncG�a��Kk�e�%Ļ�,��Qn2�v�q�;)�����!���*�����쉟��{��+�O��U����ăcB�\��;sm<�*� K�&��l@G0"q"�JVJ�m��L���M�J�W`�V��[D�	v{���m@�"T3`�F���Û��Z��������g��R1�o~�L�=��M�C5���d^��e���N?�{^I��W����}s���,ϟ�1 ����YI ���8�h�eLq���iƒ-F�O��L�X���(���Y���
gS�/�,��e��7V��$�i"d�`l��;@6�Xo�Ul�	bU�9NV�%VĬ�{1x�QV��S+Ɋ�|��#s#�ˍ���Q��#�3��f�m�A����,	Y��<�zУ�=;�m�M^+Q �L-:�>6�v0[�݆,��͈\���zڭ�>��!}�/�����?6�7����\_Y%�;vl�����a�b�wWzV��*�F9���k�������;���;[m˪xD��Z��Vo����j4*F/<����Z�V<)_��p����\<��&��E|�B�[�
�+%_�Fb�"��j�?�9��'O��O�U�����x~��х5�Q���5aa����a����V\Z"-pq���rm��r�JO@2�!��� �E��+?~�y߼���p���+^��O|���/���3ꩾ>]�����I�����7���[���;s���a��3�wQ�K�3�+e~אR���r�����0�
����Z�"��Em�	�0�3�f�5�<�����t�ҍ�'7wV���0I8�%�$���X��{Z�d�X�<�2;-�$�G�!6n�R�B�yR#��u�Mb���L�TMx�ז�#R��UV�"Di��O�V]�Ƶq�����{��ܯ��[�����;ȿ��y�Z�j�����#׮��>���=S6Q����;4����r�<)�2��:�C�`xz�~���~���0�q]�A��i��KDk�1E���{��k��B1yFׄSD���$Is�}{�Rnԡ�������"j��1��.���#'��ӯ����<z�����Z 8B��KxY3ɤ�G�.�(���I1Fg�)W��&�N(	8���n����s/�Z�)��H/�#?�щw�+�m�a�SQ�����㫫�/��<g�67��;!z�ސ����ȑQ�_�����6�<K/{es�[�1_�����K�1���D�>D�_tk�Q2��q�h���4TZN���Ji�h���}b���"��~=`�a�0O��J�[�r���%H�ED.j�YI��l�d��������e�iɒ�lc�UV���X�89��D=�gl0�([3�)�����C_I=�>��~����������w�����?��?��*�M2��FBNe�[���7־|�Bh-D�WY���B��ڡN�������^򙲜����l�䢎u>0L����o#C�}^��l=V{2����Z�Όj>��J�� a���Ba�3�e���{�WPI��Qo�{��nRd���C�,�nu�+��,��l�+>�W2�&4�R-��Qp�=6�L���z��Ʈ&"ZRz�V������=�?��?��~c��W^�xv�c,=�C�rG�����>��D���N�Ů=�����y���ߘ�����}����ܓ�?�m�5�)-=� �W>�F�`�Tf�R���/ٗq!�n�L��0h�	=F�pf� �Bz�����伱�E�Օ�=*^���.�崾���d�4&?�4���v�W��s'����fB�,u���h�)<>Q�ax�7f0IET0Π�px×"+�r�On�gx�f�w�����Ge���@�
x�½�����0P���r>3��
�d�z+��3�?�����YїW�wY�Cḑ2��V6u zy(LtB��D�j�:�%��!z����ƌ�}�<��e�v��sB�l)EjPfm?�d\�����mtWB_�s��cNm\/��e����{5�d��%s�Ī�kw��E&�a֊Vx��{�m����������v��V!e�Pd#��-Cؒ��l���x�<�:v4G�)I��p���wj��#;|�h'緩�1:Gv�
6���]�ª獈xʈ�X�o��$[�#7G9�}f���軁��Sc��snV\mSt��MƶS}�U�RB��w�*�1��f��E�I��t��C�<$~��\�5�vT�=Y��I;7�T��)]�D=/J���v����mn���?�������[�����O��+�֡��Oot���2Lr� \9P��
��TtI¤ŵ��2��s	� ���e�}(Ip�*Rz/���
(>ʚ[��Ԧ�{�a���իh�9s��1l ����Ŵ�tN��	q��;�W�Aq4�K0�S!+�@��k�Z%��Q����F�e���B+^LΟ���MF$M�+!��D×���Ҝb��^�2|��P�P��ՍG���m�}������~�P��U7���[ۭ�`Z�C����?V�w!WK���9b���:GV^����	�'�}���a�A?�Y+ha��n�|9�������J�J,a���-s�ˉ@_\���B��Aq142��.%@���Q����ki}�;��fZ�f�'��Lv}����';�mm�(�K���Kn(�_e�^~3���P.�hZ�R����$]"�k�0�8U�B+WO�a�(�[�lW�|x�����zR��w����������>�w��l㍻yz{��/(��}�Qo��B��܄WR˪rC�c)��5w�}�ʺǵ�MiR��-:+�s����D�e�zxSy�s�f75�n��=J���'�߆��4�Ad�w�(,���#�5#�0���aU�v�/�x�o�)�/�B6�<g�:���Y,��m>����4?{�Q���e�oJ�#��n�\_��2h����~i���.~�g_�y��� <kt�\������#����� KH�M�Z�8S�v�3��cA�pC���^q��c��M<��~u�P��to7������J5V�JK�".W4\����I��XP��~����6��Ƅ�c��˒y�����<g0�����&:i���2�>�i��zQ��3�gp��E^�u��(�0�C6�d
�|Ҙ���&����N�g�[hz���4�د�2�q�5��K]����3��Ŀ��#�E�/>t��}�߿����A|�ןP��ڛ��ܡ�[�O��,�7څvҸgyAҵ�6��2�4�}���g�Cra�_��:A�	~n%���=��$QZ^�o��c����Tᷬ��F�F)�_�*&6t��Bf蟆2Т�@<�S��C���j�s�\	�ZA� W��d�7���Mu߫�xN� �zē���;s�j&�w�٬�v��xK(�(?��6�7�0�0�g�����j��o��zx����<9�o��*���/T�Jv���D}6��ۇVQr��x��{o���cp����I�D �ߢ�+@�-���\E�1րZt��R�g!����$��N�K�MQ�ezN�4��0�D��1Ӕ����Or?���X����<Y��&��+M|�v��u3��d���vn���c%R-3
e0�c��S��F-C&)*�x�Z�=D{�(�Ɵaܦ[���Z�6��y9%�:%�u�z��vURm�<f���0�bhwW�,W�{��c�k̴���P����7����%��	�x�ԷE��Ⱦ�-!�`]�<?b0L�p#W�<Eh7|�zu��(㸀�0�rA���)�[�_m���*�+��-�����b`6v9��PYY0_��2�u�J3~@���@��~L��mQD|5q��4"_c��#u^��!O�E>S�3$TGcm�j.g)����P�4�G�|7
�������3�BJ_���2���av�R�>/�EyW��X�<;�5�g5�8��=w{u���;����z�����r�N��d�0 o�������^����ޖ?���]�Zߙ���ƾ)%��]	#�zMG�YՄU� ~H]Sɚ�H^'�m�����Ub}��_����u��8*E�0�pQ����:��+�NV����axv�\U);��Kwya�������!�����',��N��~���~�<��A_���َ�ׂ��d��%�/����&����'���/O�����8�Ш@s�i|�vh�)�&LĀؤ���pU�e�c�_��qθN3av�dÌ��惖>Q)G�,%�:!��8�
�b����F��;>���^�ҏ�{�_�e�x��|şV#�n#�$ s�h�������F�T��O�k;��3�����ŝn�zʋ%����?�/�'&@M���((N�y�ꥃm�D
E��x�c�@,#<�`�qޗ��B�He¹�U�}5�A�z/OvU��]E�=����j�]�Y�^&˶�kG�\n������G�r�y�� >��'��#��gpC���Z�F�S�,&}�oNC;$�CI6���^�H}��wE)<�O<1��b���
+����ϸ�{7�zW_�uW�ſ��wo�%,˴CA��Ċ!T���"�Cd��Zg-�����f���/�����A�������J��BM�R�����e\(�7+�MM��6�4�����c<	���\��� :���[`#�l�9�-��&��6��q��	�B�`�-~σ6�i@��*I�ɋ}�=uY=� E[,�;��/\,$�:]C"��T�c��sZQ~q�����N��9c��}��k�_���톆���)��L��^β2Rtg�R���54<�����4z�V�=��J#DZD�[�������6���SA'�1�VTǻ�p���n\%e�� ��ڔ�I��Ӿ��H��É�-��Z& ��1��{>(�F���6�\�7	�:���n�2�cY���#G6��Y��Û�WnyƱ���l6x�[�w�_ȣ_���u^q��BI~���S����E��O��3�Y�6O=L��/3�19��b����_�ۜS�}���/�lj�����M�ɯ���x��_���$91�Y��9-��0�~�(M�yek�2��e/�C�-�|��Ȼ�>��}���{vΞ�R+d�Od0��.�#��vE���q�Y���&Ȯ�ju�h4��a�TX"����V�0��" ����Lv��̓Ɠ��m���/ ��Z$�����3U�t�،,����w�аMbv��Nٺ_3DxItqT����JE	~<P����W�HD!v�<��#F;&�-]��ݘ]p�˳��cu��u��?��g�è�eR��)(�������[[!84�����~��XF����B8�&1fJ��"��S1e6#l˚�7ױ�i0��N=r��n�E���m����[O�c�\�>��$	�3�M�KL�SJ��Ar�3C����O����8}ko���[���[p]�@���d� +r�e3	w�O?�����Jt�B����,qɕ��r��c�}L�h���ą��R��s�;�K�{�?Ԓ�V��2�I�b���]_TvxR�8����F,��љ'�i�)��V��V�(d��v����!\�Fdjo�	*аxr�����W&~�f�{�s��r���h�x����#�ϊ�Sn���F�V��$�L��;e&ˤ���te%y�u�ԻF����/���O�q5?:��L����C�8v��j*,?������ �<![�uR���,uWh�m�(�c�r�^�>�	�_8%c<��j�wV}_Q���k�� ��·�}���O��Nݧ�j!��C
�g"��?�+�6�~ݑ��߃U%.����N��?���3/�+�#�����b�P��yR�����D�P������v�W�Q����๲�����n�K7����od���u�˕G�ky���r�Չ�y�����k/E�_�7md2Y�pE3�@i^b��L��|��1_�Ӹz��3��V���'{{�׿���#��?��tR��ro��j�aqB���g"�L��8[e քE|"B	ʠ�)��k��~���]���}�k�AH�X�j#�y�B�W�i���l��Q��HZ�]�����'��m��}JJWR|v�\�։�D���6�l�tᠽ��k(��@&��/tM�:D�(���������~�o$��BC��U�@[�T�/a�t�N��sm�m_1	T���/����/�H�8)���]tn�_�_�߱��{bEY(��I�Y�XΔĢtOF��"�$IA!,>h���#��/"Ų�Q2�H$a�eKm]�;v綱l������ny:`4ѐ`�0R$qՕ"�9W�j�Rs�/7��3�*��PJ�u{��a�҃���v��	�?����<?�w���zw����Y6� ��V�K�O�u&�������7�ޖJ���a�a[ p��.�vֈ�����Y�0��[��)3,)5I�d.\���̩�aԠľ�,9������j��O~�������(�1��ܨ���bE�[@uU�A6m��̂ ��c�.2`�rp?ֹ����g��_��v�����d9��+j�%i��V��+��hq���������Sm��n����������%�hZ�1�2���}X��X�R�A���y��x�=֐ix�Kؒl�3R���>l*����%/J�~-Y2@���-L�!�����ؿ9�2/Ӑ��$!���E6xI�S������ְ��H��UF����\t�Hig
�q�/L�F��@�����R����#JZ�E)![��Ha�}H�b�X|��"�Sr�����8Ψ핊�l��!�����Ń�{/���q{�!5L���c&1S��Үj�0�eL;���DL�q��b�i/9�g�H���vv�TI1Y�{y����`�|����4̋��FK�ȶ���a��q>B2R��7��
C���<A;<�ɵ9�O���݅� [�s�$��m�ř@`|����zS_#r���'ıd��'h�i+�w�,J��JX�
1�1�]�X�;0����PL���{�����N?�ߙ%��� -���1I�&��&/;������M�`��f7��L��#�/������7[]Z�$U�=��R�\��aV��E�,0�YHK�mҢ%�Jj',q� N�˩R12SC��e_�[n�b�+yB�]�>� ��L������5L�����PQ26�C8���am*���B�Q$�g�����;W�Y��Ӹ��a�3M���$P/��!�z)t,@b^@�ow��;�E������(O���'�ʥz����ơR,)�B�W�B�����:���I`4Z/������w*o���d�!lRDc�P#�Ԝ�+!������"E�|C�\�h]Q�\���/���h`B'� �cq�p�l�A�]_�UfL1�S�#u�K4+	U�I�Xo��ū�hV ����
�z�+/�����+��u9�C�g���Yjhdt ���I�5��5'���$��4̋J�g�!v5�������Do�:��V��X�d{1���Ei
5�J5���U�ʱ~������UK��M��o��x�������T�VJ�j�Ah��'{8��ϖ@�q�p>��(�QAXRUg7;�1���e��#_��d���^Mǵ�j���\�� �D[a�e�0R �院���T�ƊF�LWRB������"
�����eh�y��IBA�_���8P�6�i���F
��+�����i[-�ߐg�3�X�3=�"H�ҜG�0�v��K�ϮE~=qrd��Z\9�鉔)�K�	%��:�0��ªl�&L^�4��^�
x���q
�|D��s���S���lr��6N)�S�2,ЇZ"2>t���T�
�u(u	q*12�uM
S�(`�3�QѤ��h|~K��r�N��c�Nj߈:y�E&Я��V_Dh��|�;3�P�R�M��B��J ^*�Rz��Z�P�^�Ydf���	�N�f�3Vm��>��Z	a�ț�6/	�5�	s[f�`u�G� �
��)衵��H�=5�\1Ք�[��2C"Kjs[��h�t��%�`��<�9N}����0�X�y�3�Y�WW���2.%C�J����W��0�м*|]T5c^A�{�G۷�L�{!�h�[9
	R�����あ� ��Jb ����J�Ou�����j����~n�ݧ9	5<���+�c_[u|^��^�m&���l��އ�b:�ς%�IY:;޺��M��ڠ�Ț�T3l�`���`�1����>�0����'|�g��ewr�t.sҿ�8�jnj�e���Ď�D�����1�TIL!��W�Ʈ=�E	o(s�|��L�AN��0R��@�t��ʐ�#f=��%�6�������7��g���j��qBK�^�0I�ݦ�d(��W��*0��F#*+�	���E� ]�ڂE�4DJM�Hq�Ki
�}$���~�'����Rb�~
�,^$gZ�A�Jy".|2�p�y�oa��b�2
�v.� 0�q8�eSc��bb<]�N���<�������%E���X_1 9��E�ľɆ�K#t�#h��D�Y�_�f<�w��(a��X��ω��a**1&+�ʩV�D�n��Bi�X6�h���"<xp�Xn�'���c��Jn��>�ig�R���>��2��Ŧ���׫ƈ������ᗦ��%�e�g�?��R=���G�D4\���3x((� �©�Mm�A\;>��4�ތG�l�Xy�Nu��B���IGJr�[��$�u�Yy�M�ߦ��4�#���"�  �ԯ����t>C��g@N=�&���1��Sq,�f�Kh+�嘑j�~���d��څm$��]Y��7�ZI��sq����m�B�.B��I�RҹzZz���ӆ3�d�� s�ŉhA��i��$4�7R����+��̠MA�"<��	c��4zE�]J}	�3��*���f��>��g��7@֦Bm�t��C!#��s>b��D,�����3	��π����a�Tw�Y\vO�CO��K�Ͳ"���\��7���$��sMX�'37mb��x�l�G౤ͨ��x�5�ˋ�K��ϗs@b8H�J�e�����5NN��KD��0Ŧ@g�G𬒾�jN��&W�J�}D�XcU�����l��+b7���t����M�F3�أ��
N#S�19�	:�z�$O��b�#��U��r8�	�Gs��Z�/�2���I6�a=H��ҳl�~��M�s������L'�&���$�l8��G��nD�#:R49�v%���UA6#Q̩Ĥ%q*h:��[X�w��\�8��1���ZC���l�|n"�������{�:���3Z���#�4 �Eh��Q+����)�������qN���m;��|��p���$�j��/��a����_~�V"�x�-�F�IY��EmF.��%�qqɾ*\��<]���	��Q���P��Q}2I�ڒ���H4ѕ4��y��qIX���Ǭ&�x7��%�ym�1�0�R��'��75|��l1DcU[�o�]�;�ka�cZ������+s����./�UN4�r�=¤�,"�������/�%�	��gr|�ѳ1]�U��#�:C�;oy:��'��c@]�@uo� ��+��h�Ԕ<�J����(��`�V9'�T#��4��Eq�0>o���~�ƫ�l=�f�C:��L�����Z��И��� �Ӓ@�C�+4�/��+}�!�0)�0�3M��+��u57�C�Z�L�ː/�����ڲ ��<|"� 2��
2�k��x��R&�E&x;���Q�
2�'��D'E�=c}�f�k^\L8)�6�`���>��6����ڸ��=����}Q�h�;�d"w�H��u7�M�B���,���J�ऍ�F��:���:4�00�Xf#ࡺ#�!\��]��|�ʳF�)5��� w�]>�i��L�D�?m��(@�[����pU&�	�k6�U�v;�+����厡t.(�#L���o�����@'�J��w�ҚB/�[-)�N���9c�7�O�}��<��)1��:B��P�=LtB(22�ؽ�(1c�z%-#����in?���T-�zJ�'�-����$��=���A��|%I�Ѫ,|�8)��i��z���|yY~R.���hؒ�@i���WVtU�y�Y�b�IO��� �R�u�<ڡ�Ԅ�hFEeE����RJ�&{F�ci�D8pR�b�3�p����26�[�w��Zt�x�g:8GM�\I����8�7�qnYq@�0F�ӅX��|�%��H�qm+��-l�MNaZ�0R1[{z�s�m�\0>��Ǚ�H���t67`��,���
�kL��1U�3+A�����K���>�_�>�*��8�f���,���Y�5���uk�
ǤqmNt%y@J5�-;A��e+���c�i���l�7l�6gz=퀗4���Di��\rćt�Œ{ᐳHp�R�aD�zg�ݢHnl,��9����'�o�)�매`#�Q��(����V�F��u=��|Ţh��\4I$�����ě�D��	���K05���bz�t� �܊PP���
�|M,�g�z�Ձ=����h��|Q_3�t���0m�uI���Faj�b���>�2S��((ԧIK'I��:��I��"J񴨈��8F�sM\���#MG���jIzzU��;��[����ߝ���$���H��������υ���� Za0�	�L�����fa:��Q,1P�� R�4����Pn�Ff�5��ڻ7V��nM�h�ZS"���fv�"4��98����Z)6U�Ə�X����d��i^�-�~13��H�w߼� �(b��+�Rc
�(j��e�ʜ)��4� �aN�i�&�(B��`[�)+/t�_i*��0Q4������'�H&+��AP6��>�\G��!�L��B�`I>T��~؁���8Q�cGG��!�%r$�86���Y��O�H�8���H2�hJ8�Cfr���8l�9��-0D���Jh���t$�t��rm-Y��c/Վ^����eE*�5�2�J��DѠ-���tJ�4Б�:�ˌa�s��xv_-:E�G��v<����3����"i"c�E?h
��J�0�g1y
����� ̸�̾I�9��-#�Z9�(��D�Xw���,�
���=]dc�s�(��\��Z&?c�R���T�7�[�H����d�"Е�}տ<U�8�$�ig�M�E�9	!����U��l�13�IB[�N0[�`���z���\V���i��Yr�θ&({��#U���O^*���ZIV�B��;�?0q�a�b�i�VhĻ���bRK�aufb�#���gEE}r�ʈ�?�Ť)���ߥ��M���%����]���ir��>2��W(B��@�d�
�R�F��̻��*������d���"<!�b�]����r���	�S��͂Cv4�Gf�&7S��N+�����Fj@y� -��(.X$��o�v�Rj�`�~�)k��Z��H-��Bf�:����~�ii��˪B	Sk_1�6!�aRK�6it���I�p~����8Lo�?��q�D.�j�^��3�6�T�MG�"�Zb3�$X�4S"���W�����&~���o$)M�R���湙G�<�M%'&�h��8;^�O�@��z)M��k�j��Z*�+��er�3�J�({�4j�5��.y��$C�b�$0����3Nk,5�s���%�D�C%nX ZQ�&����h���ԲU��1C"&��ĝEH�6�'��)-�;U��$5��o4h���<��c����KC� ����@5���E|����hjp˴�+ӏz{%j�X3�eD#)�Y�(39l��%)�,����0�W�d$�h��G�T�RV�I� �\�>���~�me.t~'�`M��1o�8�������Z��ra0�e�^�f^'��Nf*�9�\���i�M,n�h���j���x7�~R� )y�����n���}�����љ�~+�=šB�)�+A'��= V�l��H�5Q��kn�!8Z�?�:qu�����pǿ�u��n��w��'G���f�V[I���K��[BҁH�V~�
��eM�<��s��z{۽��`�x���\13�:�j�TR��vЄ3�uH�d������D�*����G6~l9|��?c�ޢ`T���&�[P�ײ@p:��}^(M���Χï�G�w�:T= �i�Z��,˄�ٞ,v��`]�?R��'��@�M�C6���UX+��i����>�@w�]��;>6oc�V��Hu�ݴ����fK�4E�Ŕ\Yd����BN*����iZ��%+� P��J���2� <�%v�B�g���W��m�\fsU\&�Z�dI���2�s|�jc�Y�}lM$�d���n����&%߶�v�1?�15��4kN�%��/�yXE�q�KH
�Ǡ���*�M��7�w�����W�z$�}�W�G��rs$n(�I��ң2reR
2����d.�$T�cF���+9I��`���y�(C$QZ��3I��U�ms5�[�U��~��*�d�4KߙA���h��ǡW�=U]���Wl���7>����������Y�*�1�n&��Ao��n�|���2��&Lh��3��t�GF�$����h\�sBK�����m���40���36j�)��Wi�01n�{�~���K�Ef�Es�ڹ����sO��{�$�^*,;�Ak`2����׿�=p&�p��Ɂ���Q��H�#h03�)4��1��������m�2�d�Sm��X��2Vk�w�:��!b2��&��> 3�pR�!��G�q��}N �D\�.��ì�W�Yr�l��}��?���[��o��}}\�:p��{E-�}��PU;{�sL|_������Y+��c)�rsVn�v�Rȿ�_�c��v���W)ܹ��0�U_F&���7ݖ��_@�].�h��,��$J�i,O��ޥ�[v��V�����|㹇ZW����v��o�ݥ�ҞǸ&�`S���j'��S�!�N�ը�цjl���
�	�3S~�3"���ƶ,%��R�����qa W����Nd����LOv���I98��k-�,����KO�=(�?���>w<;��+}�qB1a`��l�h=Y^-z�m4�xO������~�:�g)镊����Xhۮ��MV#���V����)j�5f�8��w0ω�Ra=��X8� 7V����Y>6N8���)4�b�߼w?�y(���D��?��مG������o�}���p�k��'���"�z���H;����W�,����RPZ�ԻRQY秒�'m�8�C���a*JH�Vm��9N��q���Gz?mA?���o:��j��'���/�s��ڱi������3��s[�߹F�� @�?, �������?y*L�f5�/;���!�h�j�����A�Z�(��Rj��&B�&��2O��Ϗ�GJ�@z�8��5�̊�<j��|n�3�;QD�6`Њ�<:~�?1H�m$�z�����#����E��|��H�S�I�hp�s���{�9��׽:�t�H��=�M���zY��uG���+Q0g9+�'�I�+XA�v�O��hmF��p�0��N�ct4Nt%��ncH�	��G�%���[����c��RK�J?���~�Q���X����-Th�(֯�%M���[��`<�i�B�}�T�O��
.G��'��|�wGO�8͆��g��+�d��)?����q5Z-/��p��c�(z�k����߆W��w%��׭�u�dA�dd�T���+�� N�G��KD4�PQF2��{>�X�h��ƴ��!�H߅�=�[x3�o�1�X�
C0t"�2J�~�#!�q&^�^���M�{��h#=�lQ�	x�^uc,F�����'vv���ҙ������'��ǊB��0�^9tI`(D���s�ݿ���}�g�����t�e�]U� 
Ct`
"���1#��>\30�a0%g!�ep/E�0c:�QUL�mnсrV�w�h�#�y�z6�(�]�P�Ʒ�Z���Ef��m'�Լ%<��}�㽕X&/M��w�D�64����FF�P���������kQ!ߟ���V~N���y�&���>�W���B�~���I�&.��(�0jh��ě���ua�63�����;��L�0K׻�8+�{K���k�B�f � �6�"S%�9O�I^fg,ѮH�ic#�&A`3r�8�){�������DbKɜ_��?�W}8n_�h8�m���XM�!���@FJ=PD�+V���)��6D�qő�=;������y��ӮZ�R������G���U��D���$������7|�;B1�P)��)ZkyBl��c�}�s�d �~���z�1c�Eb����Q+j�త�m(���޷���>2H_%���������o�=y��Y��б�RT�ܴf�Q4�}�E�'ٛ�G�שּ䓝#7��Z��A�8n�q?@[_ZJ��$�>ce�F��y�x�Q�)ib��ƭ��m�@�(1x��cF��Z����j�c�s�xի�A���\Q�D��Hq���oP�Rz,�O��(r1D_�����!E�X̺b�(�q�a1侢��z���}x�<�T�S>qYP�j:mm���w�����.>Td��yS8����Ǐ�-�r��.*
�b^��}������a𨈯���������<�-����Y2��'�KGfb� �'���Lpf��,�<�~%��d>m�������QQ )V�җfᔆ����ir�HH��$��h�51ݪ>
���i�������l��c���{�K��}���p�:�Ja(�7E�N����[���]�m���|}'b�Ǳ���ë�O�y�j��{�Nu^.s�`@K��������)��:lW�9��2����y���}D��܏3�Q)�����7�oԙMH�D^"��h���l�����=v������3���a)u%cjT'q�w�T�D�� %���$�_�/�0I�m�rƱ��W��.�~��'�u����CGo�D�m~!_{���`�x��ȋXK��>Pn���Q�%�yi$�^�Ʈ��0��@`�uV�B��B����ȏd�T�=��%�2���V0(����(��I?~���W�e��M*S�
Y(G^�(_�K���B��꾁L<h�s��z�k�.���E�Z�_�p�1��/���HI2�,�\�ج,�v��H{��p�Ƞ����'��z�yj^�����6w�z���K�����&�w|�?��f���@k�Ag�\�1�z0���<	G��@Q����a"�P�cy� �9!˔R�J̊%����gOFà~����y�+�j�B��\i+�W&:�p���W���s�4.|%����!^��U�%0^<E�ò���y����=Vc��=�<�|����
?�>Js�����K흋��/�^�]:�����I�`�,��{	Z�1��n��+��n����x5�����/2�uM{u���8K�|�6�[�"B��R���"� JVЫ�.&��\�[�Q��H�I3�ԑ���eY�Eu*2�(�J��-����}�T���D&=,��y��,��uN`�>	^��O������O�}��/By���n���Gʽ��Rwk�X��{��<�{,-��]ȳ;����b���������E<V|8�"'���C�ҁ�vJm�+��7�����7�3Y،m�0��3�����̽X`�Q���H����3����C�\9b�^��y	�7����o�Retc&��X� �{b�v����(����S�!���^���F�("�W7�NV�hm�4�B�;�������z�����m�8�trWQ�b��}�hJ&���x�_�H�4����^�u��D��. ՗�8v0�8=�^U9��ى_{�!�}-�>U8�c�r��-�/���Q@9�� 6�*k����t��D��MJ��JQ;�4�Ң�F�(󼴗\��N�z��?;�}�;�_�q/��n3?wco��@�JthrY��ʱ�)/�`��g̢��������8�_�y>���s�ʜ*5Ճ�T�=��}X�ւ�$�T�kBE�<��LNdV���2cy�p:�==��y�h��`����~�]6Ufh�������n�������[���VF�}����tم��`�k��;�i�7- w��6���+�7=hl���lb����.1���Y�lk� �{�mVP>�&�]�����!UBPʎ����������zK�ߺC�-Q�J�R87��X�֔���3^y� �o������(��_���mA;(h����`�H'��i����<���ѫo��-��<j��hEȍ���w�X&��:�<u��n�a���(���E���W�d�T[�@T:�Rt���@�W�@�q,l���|�8,і�����9��U�:��`	K��4�ޥ#�l�|��M���2��*m�$�j�(����cD���4�!��HG�H��U�����yIV�CU�z�@��V{�'�`�z*W��JѢ)HI0�`�Υv()��Pk\�˼8&Ӵ�f���!P�o�Y�l�ɶ�ܴ�l^x��J���ØF���GU?��Ҕ�&�-�2���Y�JE�j<ǦÂyV���6�6��A��?� *�M��PE�y�S�y���,?e�"�R(�'���D��(�wisP�/�ӽ#�s�ţ�͇à5 /�x�@yQ4@���3�1�*2�j\wVo {�w�Չk�l[���z��=��d~ӏQ:�[coT��nF%yy�WC�r����
k�VYSk �":�p�Xo��[[o/{�OWwkIw�����u?,�d* ܖ�A�~���;Q����`��G��^������&���-7%��4-ߜWX�3S��
{�%>���J'�8���-�B}Y���,3Z�6��:�r����w)N�悲��?���4��X�'���w��L�����¶��
�)C��JN|�N:���g� ������� 䩳�kSui�6�:��`q#_�!.��K��j҃g0���(a�����06��^��@�]*���)����	h���Lg�L�+��D��H`r����9�:w�����JDa�b;h�K�����i��P��؛�Ft�0K�\[���[�����
k���ͨ���q`�1g��E�GJ�����a��ķ��to��}=��`YV�g�C�_W�ϺʨT�<���?i��ڕn�r	�c�K����N��f�<p��H��ʔ�):Nݔ�a�~_H�ɧQ���o��b�f���/L;jo����/�9��[��i���}Ne'�,g�":H�����K#����V���f��D,�GԷ�$��h��M�&LCS�xu-SG|2��6+9al�{f�ފ�9x)K5���"B�,S/����[�R�|{��<V�G3�9w*aM	 N��)��{:�<��1�����aV�f������s�q����3���>i���|�qd�w��;��&�(�d�c����j�<��<y�,�����x��d������%q����!��m8L>��Kե�f�F_�FA�F�ub�u� fP�u*�USwg��^ҝvr X�}�s��c�69蚳��IO��ײM.��=l�N��������52�[_�e
��ϥ?l��c��h's/ ���2[�3-9Uw/���
Xz��g3Y��̻�4c''w,�~V�����0YO�M��
����mm�;�9֖�ac�y|���<��4 \��M7ŋ��F��Rz˲6��m��9��66ȓ�}B���gY�YH�%4H�2/�9T���u<�t"��k�}]�R?��Jp��f"kU�����Xb�_m�,\-��o5ͤs���5�`N�̊��3���{9��DMqíYN�sb�{��}?����*���܊������q�Č<㍡�P��b<��֢N2`OO�")����&�am��z̛��1Lѿ�zn�q�~O�[{�e�_��v9�1xc����������L�	9����P)g�C���|x��ә��ls�xrN���6��q�Qi�i����b�4�=�*�m�eS��)a�3w���q�ݺ�W��Ye{��ֻ&m���7qJ6)¸̖5���b`
�Lo��f�On��d��?�w��[G�l@3��ڔ��.�Fhb\�q�Gr� 9�����B�92�}���ݺڃ�Ʉ��s��n�UBɘ�˘*�l��.��LsCL�s���	��f ����i"Hk��aE�����훹��=���@��c�F��d	����g��� E!9��A�PN=�>���>���͙]v�-\T�@f.ĬL�ː����?J�d}�]�SX6�{[C�]�u�[Ƨ�h�����	s�J��dT���3�k�i&�F����n
�_m3�]�uܶ!��U?\Z�w̼��M���e�h_�%��x��A���c��j��:�b�s���B���g�K�^)`��~���29� '�0kQX�g�a'����Fw��	�5�S����ܵ�'U�L(�	7�����Ў�y��>��ae�1S�/X���>:Y��H��UM���M/�Y؝�֑�pڱ��0v��i+�?��O>C��i�>������󘒉}�5ea�ɞ��t]Fg#�J�/Ox��6Sq&pC[V�8(�u�����
T�4�
"���D�1� ID܉è��!a|9:��������X���,<`�+L�#���)�q۽m�x��?��B�'�TҠm�H����(-��;��d��Z�Pω��1ͳĜ�������ikU����q|�w��~a@�����x��J5f�$�Lo">����F�s�$�G�Bp`Ť�i>ۯ:���sw�e�*c�2�4�Z��2�����������h����l\W2~��0��Ǽ��B&�V������yI�$Uĝ|lx�5PB�⼆�81�Gg:�4v�Z3�.DG۳��"V\B_b)9s>~��D��ҽ���j@,l&�醰g��#tw��x��E
���\(Ϧԕ�pѢfU #S�g&Nk��_֖:�U���sTV�*T�d�d�Y�3���L(r��%��-d03��^OL(ʎ��*��Øμ؏�s�2}ȉ�c�ho��p��E�L�>�Zx��̾������)��$�4�X�9�,���88��S�,���ye��e�M�lm�!��>��*�v�"����B	[�O$�t}E(Q����-���H^NPZ�"~Js �4���HMV��:p�`��4[a�wy\�F�����Ԙ�Uejl��.�S��B��E����T[B�c� �#���,��6g���?~v��"��8����M���O��6FIU��M�h�UzNk @�ybB˞���'N���bc�l��_GP�A�?��ج�67�D����h	��p�+�1�i:��N=�����1_�c�!"O�F�8o��H��%x`O)��b����aY��]�C����.AOSS�R�h)�&���� TH�#�x.����<�JkA�N`S�-V�l0�B	�b�ҤyZj)Pjd�a�����
ep��/n�(�$�@Nx^j�n	�� Q��C�(|��O�\��1m���P��+���1���;j>zk��,��b��Q�/�,/�,����1Fcek	W�ٖ�=�Iw����2�?����
G]1~Ң
W\q߂)�ǭM���� ���۱+�3�d��L���;o��T�E�|���iG����z�CC[��/�X(�L�K�$�y�]5h%(M��d��ۺ�:I�7��8`�p���y�����׶u}�	,+�BGT@�*�?�D���0�Z�q��q�2���^Z�FϷꊴ1x����2J�Re�����"�,��^��ϵ�Y�1n6.�i����lsg���"ȆC(Maqb�߿�V��t]V9J�X�|��y�nLJ���١6~I���&(��[]��t���bd�Cٰ�{3��e�w1_�۲�Z��*�;k!��pN���n��o���s�*a?������>�m����g���}�΃��'�F�_�n3ԉ's�r����h�J�/�_u��YV^�(���RUʚbE��u:���](�⊭M[�� ��
���*��*\	1�(T�B:�2͡���_�F�!^q���SO=�pt�R��<�!n�%>���T�1��"��̏�,=���#�(w�d<�V�����QC�`e唒�O�1�7��Y����1K��@!��5���x����m=nBZ�N�@J]`�߄���ZZ���T��|oڏ"S�LV��J��1߃V؂~ox��b�𨨕'=�E��<i�"�,���e�W�Pt��%��!�F``T&Wc:�:1�C�,�f������K�4�(SJL@0[��F�[AUV��7�`��[u߱#&	|�wQ�)���4VϏŹ��оw�~��2]Uh"{<��L'O�o���Ą�^܏�M�`P��L|��;j��խ=���A�olA�}i��d�s�Z�Ǣ!��D�k�,�!/$��վM|�/΍p��s��9�����Cėts#\�d�rM��a�/zG���?½��������ߜZ�����&��|�$�ʯ���"O��� ������H��U��7��U����n��װ�fK��E�g~F��m�҉�.�B�����0n?���+wvN���S���fOV���~�%ɽ�Ó����8z͇}����_�=���?�'�ꄢ�4F���q��~ꓟ����?��"���E�0��c�p��y~>H��!s��w��+�{��8q�D�9��o?������vv_��}]��z>��+ ��!�u�4p�~���H{��=+++��~4"�@a�5nD�W���`�Ub�1�(d�m�l���|�	��7��P+���*D����`u0�]�����b�w�}K�0���zk|Wxo�*E�����0��ѕ�?[m��ԉ��\�,�#=�C�P��3I�� t#;@@ǲ-�{R�c�5�X���QGG.��g�����`��]�K#�� �� Rc_yJM߶-$��F9��eG�Oۍ�^.a0��nEk2����
>tۋ~��u���k��|��ϝ�x�����W�����-VP���y\������������͏3ol�J�������Uh�a �[�]rqυ�y��41��"Ӫ	W��s�l$9���a~�KW�PP�SR ;��R�}��d��/%�
�ڛ���_����m���<�ेN�(˳!+=DՖޠ�,{v�"q��y���o���Xt}����_���w��������c��!�!�"�9�����=�ko�~F��>�LM8�(�ڎ�C�B��d�u���/|N;��q��֬��Q�в�hU���ě���� Ed����l��e���=�Y�~~o���gc�e��1Hd,� �@��ʺ�J7�ԧÎU5��U�{w��s�9��Q�kW����� �x����,�Z�_�4.�}lзp��d�J(�Hī�:��'��c��'|��z��{��:�?1#xN�#ޡ:��!��c�'���;/�k���_����oKO�	�[��fy&��]󾘰͸����6��� S�͎a۾��s�?���-��b��\�_{�]݃?x���kPX��W�cʴ0�ڲZ�"F����6�~�l|�ҙ�#������x��#�35NX�d�V�Y���9���o]��U������8�y���&I�P��--O~e�ߦ�3�@+�O\��.ē��g�?��_��os�o{0���tZ�w�D�M��\T`u��{%��?����dF�N�*�F�t�H?�T�$G�h�?��AA '����;���W��Y\u�K7��o,����\ui!�Z�<�!��_���e\�V(��6��ԁ��&�ʜc�0��tI4�T�}����Z+/Uh�)��e���ª���t�d����١�|FK�V�2
��h�f�:_��{O=���>���n��}�7���3~笋�+��CZ�&@�섳�ʩ6����7�һn���<��O��33g]�F�uV�]���a����SLC� ���V��+
�����F�\3�J�ហ�
�Th�����;������6IM�ZX��Mfr��~��+@k�8���⨍C<�E�;�������_����{$�(����d�WJ^��j��~�F��q�ߨ��λ��粏��<���~�k;)��xa��]��d���')>�{\�!=��-�8~`l1�@��:�0H}�%U�<���{M+��/�`�ஂHJ��9���%�g��� �J�h��n��K��,�]`��1@K���ΩV6���|	��
Zȸ�d���0�x��/��u�����>/�S�����(]��WdY�S���X5�����A���,�?�V��夕\�^�X�����4|Vw2��3.�Cx�y�xR��DZzZ�&K\�-F���k'���g��quƴ�t�@�<9�FW֤�ʋ��2�Y[���|�o����;o���c��f.l����t��v�U*{�M��43Y�j���Y�o۴M�t���~刨����۞���O��4�f��+����\������Lz�>U�f�ϡ�`�X�V�0��6[�Va<# S$�e�
 ��h�{�c7�o�i6��su��+[Y�u��q�}�����&����8[?{��#/���a�^+H�r���o�������_p����ڶ��w�'��B���:����y(�rx���
S&�m��W��U��L�Bm'�3�G�������,\ᅋ/|<��?ͅs�NY���}��g�D�c7��!��f�t�Y�ۯ�x:{ŉ�s��ޯ�.���4ء�o�X��H��
J<�U����(�O@J�����t��@���c�$� ݠ�,����W����_W�����)O�SM�_@�:B���t��za��B	㗺�ZxZ���@鍩�)V^Aj�{�\���T�Y��Cz_��x���9�뢏��Ȏ_�����|���ꨫ���鲻�bާ.[�n�u�S��(�<�}?���+e�zǔIX�h.7e���8�)77�o��6h�����J6��r;53��E���u�ל9�=�đ��'��|�_X����<��d��#��T�2f�3c����*f@�:鷍�A��4Ө����]|'��}�����׮Y>�!��P�`Rha�� ��-HjFER��k4��:��#��[��;��lHҭ�&BN�C� 1%#�9�9j�?k���M��^����;����A����������xy5[��f��B�]�g��ͤqί-��ss0��hba�P���`�lD)�(J��KB�ɱ����P���J��-��L49␲��U�7S2�F������}�/����Uo��S���.��;�J��6w�i�1;
����ַ_�"ܻL�.�鞿�k�|n�0RJ��E̖2��@2R7B�3�ը�����-xu!������v;�5�Ǖ�V>k�9&,K%�V3������^�u�{��p!�V�=�\<�����a�?t�����x�zf����J��ĸ��T���o�3���Πv���S��^F��\_'"�d�d��C� �7�B�%i$��J�TIu}�쌼��SiO�~�^�z�
��>�+�,X-!h�G�=_�խS�۱{׹���<��Ͽ��_����?���^�^����l��[�N�m!�<Z�B���#M�8�����y�bGS�G��zsy��zۛ�]���}E*��S��yw9��P�r�D5V�'�(�d^!��U[y��=1ߒ���ݲ��0w\R�kj����W��F��Ϳ�λ�ySq�wV��tz�&Gb⍬r��D������]{�7��.?���,Q�0��@�Q�!7L�N2c��t���Wkԭ|o�sp���":��$t��P�ޝQ�|J������_��g?��k_��-�ɃIo��][n�Z�V]��4�{nx�/}�GG�s2g���$|N���e�;���+�"'��#�2�A���� �a�c-_xEL7��s�vEE��G�J܎���`;��A@� F���Ăi�֜�Ftu�Ͽ��3�xֹ_{|���D��0-�4�3A�d\�Ŝ��9~���^���2��wi�P�S�S�N��k�a,-�8���ïsLҲ|����*��j_����*M������|��D��M
9�����G_�U�I������E����˯��+������ʉ����
��BA����clNSͧ3c�ǂ'��e����m�U!�Q���V���[.��_̘�\�d��f�1�eh�`��t�hb�-y:��	�~�t��e��q�ݓ�����[n[�&�`���V�����g"ߙ�~�y�{�m���Z#�BB�-P͝�	��Lkn��Ӌ
Ǜu�+2��KzJ�6)QZ�W���=w�zF����1�R��M?i�i��m"54!K6�R��!�������ۚi��N�ަn���i�@�:�7�֑o�zw���h�s/~���������T.�*�Rg�z((��Sy��(�^'mG�~\n����q����n<���C�ry�Y��ބ
YKw��s��5���}�^����H�hxF�2(�G��Ł��k��_��^��#�S��H���N�kS;�{���Y��l��-z|���X�'�"���=3.��>�oWj~FRV_х�%d��ҍ�p�U��V�&��󳽥�}�x��U��:�w�~��d�m*�#��YU'kc-��)��+�}��\2�ɥ��E��v�D!#8�D�� ���u�[X��k8O�<��׍~Ȭ@�P��-ˑ���o�1�����ۏ�*6�y�+ߪQE�,)���Kc��!�Fm� �t�a-6`4���ff'�$tM!()rr�#I��`b�@b�H�j�~iL4d�uV�}�o�ÊY��jq�"��|0�~	o#��4��Xr	��=���i�jDz5��C���$�j���|�a���m~]��M󌸾O��q�%i]JXp*
�~��<�iZ�l��$S2/6'�N�a_��v�ah�ܗP�G5��]R0���a���mKi''��i��?2>�Iб�N�z&SS3'^M���܀�����jW��t���lO��7��L�'?�GBj�F��A�w��	=�I�<���.��Ǥ�Bט'Ċ]:X��4 <r���4�2�r����ortpZA�J���Tp�u�\�@	�<ǚ�N��D������W�&I�V�Z�S�
7�U��DH���t������1N*���u:�LN�z���Ʉ
ŧ�*}Q�Qw�nL,�$ÁyG�����T����4
�x�J���J�5�77O�w�'�P�2�7{_xL,����ꌆ��=ɉ�ۓ-��v;�,����8[A��)d@C�WH�IW�	A��=x���<�Z[c��1�)j���	��hV�J���ɮ�A�.Es��¦�k�:���b3-��13�����$ٸ���!�H��P�l�>TK��{a�O��e_��C����}G�{� Q dNKQ&9���n�[�M�޸v�nֆLs���t:�sn�\�=�yGQ�I`���&�L�k�pfh��@�V��4��DZ^������c�6�,J��y1�&	�b�!����k�l��0P�hg�E���5���n�G�A�
�3���Н4�|��.L~Ɇ��m�*`�������D�=�:q�͗͵��������Ú�X�6G�<�s䴴Pϖ�Rjr���^�A};�����
c�R��!l�܈�h�|"���k��B����a����Ʈ�V��sl��0?]Ԓ(�d4WI2�%!�~նtjlG�_9Z�/<lK����=�l�IP�p������<υ���%������J��!JO�L�fI���'�I�ث]s��dAH�Ͷ0.{�Z�	y����JI���o�Z-qd\�1E�9/?��>�m��M\_ &��\К��:&#70V��5�_ɸY$<��d������Je���az�b��B���l��lqyC��d��)�i�\���� ���2�����sV��2ch���3fu�aB~�#�/�m��>��iW1Ts�u�Q( <��*jM!��0�Q�!�������=�z]��w�3��3s��g�F?�?Ǹkk�@/>Z"I �Zb�>���^Y�*ll�}.@+��J�b��A�BOp@�y��AE��̵�M��4��V�7�~������߇��ah��䝾zu�#���_�3���m�Vi><��x��-�I� ͙Yp�c�pSmѱ}b�$�-{���K"��[�܂�j�sˀ�&,2��V���4���WW�{1 ��ѐF;j"be
���[cE�(�� H(���\:t��]q!�L=��i^����қ�ah��i�q����6�F-�N��`궵�;��6J���0et�B��~ �w!�Us-|�3����)�^-YB�L����=NؖN`9����F -����o���6D�TO�,Z`�ۜ'6>��������0�^�	;];*�G+89�1Ӷ꿪�}�[�z���
�ķJ�L%Uo�w���V-q�D���辐nEe��@�@L2��f�������ELƇ|�T�A�`j�m������`��~���9��&�|Џ��7��Q0��Dk�>��]���V���$$�b6�W
��1EK��T��:v�����O��lc�3i"�8f�K�$+ӷz��ks�H2�u�M�`)���bږQ4b
F�j%���7:ST�k���E+,����d��Hjq=3�q����V~����l�:�����Mj-?o8��{�ͪ�KU�W���Qj�N��W|��BT����h˯<2fg�T`|4�s~&֖�����H�Mm���#��J�
�k�2�i�AX���7ob�n�y�?�e�⑩�I���q��*
����&x@�駰x�e�����Y"+�������4�4�0���5������@�����Ew땻Lڌ�ݓ�E�06�axцPO�W�*�	O��n6��2A9�K]�_�pm�#��JWu�;��J��}l*�|�mS�X&��͒��`� B��|)����
��T2Wʡ~ܚg�f���c�"�Ü��D��V|�Jgi�Q��ڪ1�<�J����
H���C����dP�gRI��� /���	Y�h�C�8��&ÔqYH6�?�`���X�U_? M�<���]�"5
��wUa��P�aO��i��v���JHy<���8��h�EK�,
��w�Q���Os~l�U#��D�
R'~�2O8J�;$�ljshU��h��
Ċx�r�ohp���U4Hip-�ӗ��Z��@C�����gZ�����N�a��J��li���T��ENR�3c$�Pߚ��� �ѭKIahWt���F���C�glv������	F6�n�gq�	wF����I"Q`�9�}B���Og��l"h&�(MS�3�����a��'�q.mT�G۸����I��%;��qM���XJ����F�^E�&ꃘJMX�D�X�i�-��G%~.㠙#�U�۞˼�lp�i�����T��c����%�T����E�٥�����6�8��1�L+�e� c�s:�GjQ�<��޽��!�o��*/�Mg��e.E��a.y�)�J�@c�ep�*,5E�\�R;�cscE@2,*�b���Z�.k!�1��I�y���ɸ��K�"-�{*0+�@��ZUq�{�_3��0� � e�B�<ɹ-�FL��Y��8���r�J�m!�+avB!~��vcU�}���D$0a�����B�v�06<��`���wu�oX 6�W�ީ���6%C�	0�Ih�0h�w4K0D֚��rT�%%BGV��L9S>A��L btG@���Ê���6v��,4�˩�/��/5���6u�n��)�߄�1����GL:LԐ�G�fT�/H�ޥ���Ô��-���[���>b&������|�J���x��!Z�I����X����I_���ce���7���I `��5H�m���ݜ����?4��|7��Ꮳv�����=;ȫe�'t��}ҁT'4#
�����L�͍����s\1��(�8�����B�ܞ�c�HdH�*�]��l�j>{��
��-��b������7Y�kb��v1�P��/G�L���� .o&L��[�fS�a���ΩCj&����)���� s��d*a����<t��8ƼR39iYP ����Qj��2#0��Ȥs8�Ml|%�pc����4�h�B߲�ׄ��JX�:-'&�o����(�CG�B��I�f:��<���`�~�|�Ͻ�%��ߐ�^WV����4Յ]��ʁt�r��s��2}�Ѯ����i�#H��2�\+X8��D�j	�:mӨZx.p�&T��3�u�gb>��31���J"�oC�	ͱZ)C����A %C(�z��c�W�����fj]�Sd�;�\�A&�9��_�oL6�`k撥�0��ch�k���jĵOb�_u�3�XD�&ըX�C�j8�6�!6G�Z��$8��pR31B�o���v���8�@w�s��Q�
wy��AB��d��\��&��u� Q����)9�ox��F]#�3�̪�������z݂4#ЏI[I��-����yFv� : 3;�B#|(��>�Q���6�&l "���O�`uwi�Y�1���?��mꍮZ��HХ��" u2��Z��b��yK(3���J[�2�ai�>yJZ~@�$1��"Rd�rB`*)�Z����qf4ea�&�8j���fgT�W�J_�x�dv��]�z��۸�|����IB<�Q�T��s�o��k��R(c5���;E��1VT,Y�ƙp�$���XA�`(�p��3���2!�  	d���2����8B�I����H�^'q��i���`;�<7{l߀!u������7ʂ�ƥ#|g�e \��Q5���^���	|�1�"V�MT���t���c�z)h�p�s�����@��,���~G}��HO$�$���#�p��_`[����s��2?T��:5H[��ט`%I�� �gLN���# !�P�IA��u_'���JM�љة�Yja4\ג<}?���C���!&�L]����`�Ì# Z�U�m,24Wj��b?�A�(�fFQU�kb%���iuap[0� d	b�w.@�B�UɅ��c\&���
������H͇�5���T	���Toֈ��X�a�J��$L8�o��X��3��tvρ�^���
~�3d�q�S�� ��,�!����i�B~�@�0�j���X!�7}��\֔$�=*!��#s/ _%㕺f�E�6S��ͅ�0Y+��#[���FQ�f���c��P���Bs��q�ǔ�2S�ņ���AL����� 4��ccp�Y1q�ҡ
���ȵ8%s�	@��k����"C���`�(��n$gL	}u�X�q�blŁ�N����>1���������f^!����,�8j-z�1NBHȗ4T+(��0^�T�M���Mz����M����Ġ~w�t�ij�E�ᐛ%z�I�V�j�]�z�K�7�u��z:�X]w�w� ,t�JG�5k9��Vƒ���"�z����?	� �Y�Np��qӶ��d�4���^H,H0�b��1f�LP=�����c��VP3�� �f
A��A�,�ryN����WY��ۙ��t}�&�R�Rg6��S�M�<� z�0|n���dZ�~�o���&4�D���n��6+]�J',$Z9��p����:>_M�y*��=2~��JWP���fJ�`� ��  ��χ�"4/DM2g���ve����L�
�i�^l)��{��������'��������~�/�4M��>R܁n�o�U�����t8�g�>��k ��G��B�m@E�4�ȕ1\H깅��<�
�E!F֓P$�ϡt�Ա�%I
O��L�W�k���ϥ�W�J*7[]�<�g�����RVv�,��Y��&�Ha�c�H���Şۥ��)�M;]��ę��b͗)-������ܳ�Ѥ9[���.
UCV�O�X��z�f�" Z#f�3Ӹ����<s���F��.r�ll��,�b�&7f[2t;�p =�'�*7Z%D_&F�b.���k3�*��V$tĚK��q�^������߽�jw�k߿�vV�{3A���yB2��j�F���FG0���6ա��:�4Zu(�Pyk�_�?���`.q�V��3��	�����|'���f�Gk���J];5&��<����J;�f�4�/WJ񻕎�<(Cf5aa����	�IN�*��6��vJa����b��Olxd(:�.�SS�b��eh#$AYYh�P��¤Ih;<5g�+���l!P�Z��Pf|�&{��V��S?�T��z��ц�P���f�(��}��ש��Miu(ؼ�͵�q>����{3;>P�LW�d���Q��ӌQ�?����p��	�F�M�ޛ�y�{��q���,�$^R��>T����Խ�������V4j�d1��d�+�ܽ�.ѽr�?�n�c��7LT����יw�ju�����7���!x=kNiū���WM����REҿ��<Yk�I������{��������_V��9I����W�>Q����:�KR3�N�9�*}P�WO��f�YA�_�)3Ӹ 6��2S�djB%�s���-��Z����K�.y���ɜ��*}���K������Ќ��__���Ӄڷx1��,��5�>�:*���C':d�l��z1�����C￉1�Ep��7M���'݊�rR+m��
�E���_���B]��}��"������m���0��^h�;I���lu���U�>B�.� �﹔n�Y*��d�&��p}��5[04n��f�
�Z��@��"?����@��D��,�R4�s2��Тᒬ�����O��[���ފ9�r�~F^�R3ξ��%�@��{�#σ���2�{�"�į�G�|��'�7_!����@	Y�fH��V���QW�K���O��LΗ� �L�z�ث�_�H�*bUӬ���2"66QF{�ebh�Gr%�"�h!�k�H�?���/;��{.'�o���Eu�Kp.+�\�F�+�����@!D�/��mN��MS@F��v*����(��Y�:����o�I�B虰�d?�����#奞�y���b.�R�
�q���歧�s��|.
f�����̈́(CDu�!����
�I}�s�I�L�82��d/}ޏ�����hn��4J6��LC��`��TҚ5�-��b3l��`�t��Ѭ�]W����Ģ�	��j�����5���W0mHX0��i�����/�9'����}����{����E���b0��_��>aC%d#ߛ(@*Y��̡87/\Ρ4��ީ�c+N�CW��h_�UQ)@��/�_���(j��+d�~���t�k��]����ܗ^Թ���jI%}u����u�?���{[Q��4��W��,��I���J�OO��:z/���jI����E�Z<�m
?�	�e�M�~�d�I&��ݘ	a�ޖ�\��}�i��n�/�y��?8뼝��y�t�}߱�N����|oMm�Gj�n+ �$�{dE���:ͬBf�bpL1"ܑ�oK�h��M�R�NdۓƦo�ym���|�����[M�wz&��_����Di8~r�ݒ��'��l�%B���p7� � �:3pf�3�v:+��\��z��˂�B�C�$Xou����i�RҪD䚪 Lo��gh�s�fS���8���8���Os��W��J��˧}�gg����o��O~����w�sh����~�o�������U���Ok͵淫nO���}�`��+x��B%�Aѐ�����~�M�VN�!|�i���m:��1�c U�w�ծp��Z+��}���;+t�+�{�酤;K�>��+w��^��Q_|�\��j/�A��˵(��?~�����c���Ƕ_y�#��WB���-/y�w;O=�� ��W��Q��D&������B�ш��vF�$���7�(�iyv��|���K�B�����`|��Fn��@bȠlz�2럿��sz��ֱ���;���]|7l���FQH�j �i�`6"$�!�m3O�όZWp>�~R�P5��
��6ZTҔ(���D� ��z�|��i�V�#s�^=)Z�d	�\p7���Xm� �?�
U9-�,������(q��\�/�y��o?�U��M�?�ڈ�ڍ�"������O~�����EN�d����?4ό��Z���U@*2%�g�^�(V>���_�����᥄��O��򭏾� �^�O���Z�Fth9��|O��<�̫�q9�Il�}"��:,u�6:o�N֑߰�L4t*���P����$���I���� (���c&"��S,e��%���;��U���:��t&�$?�S��[t��-?i�n���<���O|���z��=��_�ƭ�|-=z�������V$�B+
Ƹ�L��Sj�j"F�gş�>��8�2��s��8xV��3��jb�6�=�i�+
iЧkb~�EZj!�M�m�T�Ea��D�R#L
ᐆ�Pw����ߜOS������s���=��΋�4|�t��,�P/Z^k�䝌��J ����}�R��m�X��(&�dڼ1�UX�s��P��P?�{���Q��P�[E�H�����!�C�\&?�x�B�x!�0�TȸoCx/r�9�Ie�d�o��&�Q��m՝��"GX�-�Bj~נ�a���B�U�o�|�ż
�W�)'����) y�uˣ��N�@[�z&̔��`���HwLêN���6���6��/�P��A��?��s�{��4�_=�'������o�w'a�K�d�e&{���>�A��E4����Yշ1N��{6E)M��s�p���>�f.85zIJ�4�
0�+-�������N�yh�Ml�X���Z5Xc\�J�<�ګ'�]"z
�>������>ĕC��k\q��]R��5u��?����|���j����G������p���=E�3`/����9ҏs�Л�z���~Z�z�`���Xjl\HM��m�S��D3P��_�gE�H��Z�9�B]g�ƐQ(d��bn&�k.�}�?K���#��v{���¿4M���������Je6�&���dJ��ez8Ja��/m��tBű:����T�i�t�����u3.4�F}G��8O�6�u\/�x�V8Di�Xt�v�LF6�?Z���c��1�GF��#����yի��u��隇3L�»Ɏ�e��
�6��D����%s}��B-�!�
-�����>;��g^Y������z(J�s��Z�f�o�+����fz��{��?~F�'��#d�T�v�Vy�Ӎ"��!��C�)�V�k��i�:����Q�ܛW�B�Tf�x�~= ��6�G���u�m��V��>���N+z���V����oZ������Z*0�@I�:$�Y	|�B.�s���,'z�H;s6xA�15�l�Ш%��q>f�X�2�4�>�4����� ����"]�f�'Ev�;v���"�����Kɋ�ې$.;���D�t�)���$��H�˗�Lu�j�肛�l�%����Ӵ�Cϩ�#O�~gMW6�Yh�+�Ry�8r%�S�DE:�Ŝ�FÙ�$NX,C"�X��> ���3a�xx�\�'u��<�	V5�Y-�U�w�<�z���Ưo��op0�$��ݰҨ�U!^���f�J`2YFt�j|��	SB.��O1���ٯ>�" ���������8�'����;���"�ǒo��q����$v�:f�W#�N5�M�g��1��P�N�m�k\c� ԴN5t"���*\-��8�2	J-Њ�V{df�X=��z�Km����t��Ύ���v�i"%�|aǢ�z���u���3�f�39���mZ��: "a�ч�Vo�1K��Z�D�ȵY���v]����:�����5�$⥏\v鎯/.����vu��np�w�z�],�xV��/��Kj����2׀���u'
�I-��>�jǂP����r*<�ᥡ�Á�l@�d61Ia �n(\��$��<�qO�uu��Y �/G��a�,�9�L��fG��@Pr2�j���)�vx���L=[�|�;O2��
�J�lDj ����31N���_��V����Y�,&�~�(������O4:wmPs^vdI����\����V��Z�!�6*3��ve�ȯz��q�PohC�j♶ �"���o���	�o:�l�7�?t�.甉k܀Њ`NC�Ӗ�ݟ�&!o�#J)c�Ǐ�֡m�^�H��|��t9T���3e݌��h���gTf�3a�9�(��m'�TǞ���2n����A�T��T��Ȩ�@J����$py��t�+��v���e��[���9���o�;����{�D����Щ>�R�ʎ�A�<�\��+�jZ�(��6v;ZF4�(`�L��t��g6�R���Vk���u�2w�uB�z�j&�F1�[!q��)�2"(�� Q�.�ye�Q�����	(4�A�z��
}j���l�	���%r��������6J��W�M+Ջ���1�"�ݙV���v�(��-��� u^�dJ�	e��W�Wǅ�'��@��A�H�hWg2 �4ަlս� �;w��E�D$��	��ǂX�h�����{��'�m�<�^���X����Y�>	�#�I	z�f�bX[��}��/6�rw��m'\tH^p�cFb����7j���c�t
r&<�iL4��ǯHk��� ��s�{o�k�����Sͬ�'}�>R�^F�=��i�p}-{��hk��$�n��Bf�Q?�W�j�Gj�>�*�6̏B5g��l��IN�j����	�J��l��l���%,R���,w�BR)ڐ���#��6,�_^S
P�Q�SK`����n%�c�Y:��g�g����X���7x���W��<��B�܏�}?@�o~@
^bEVSu`D�٬Q�o�^"x\�8�;�!�4�=�����7�(��������S�uU��MJ-�k�4�V���`���d~{o�M��Jʭ��{��!˨Z{1�~O���Tll��E�d�AɅ�������R|NiQ.ouG,�I�q�
��[
�w"%��B�k}��y���6o������y�D{K��,�C����L ��3�@,��C�铤*��d�3c�?���ȳ���UuEبZY���S�wFT&��Z@��#�����lBYh�I���3��?��Żx��YviAZ?���s~���	R�ytqv�<N��S�$D�3
��L	}�a���4U�G�8���(므�q�CY]g����� �pu4Agr�dug���0*V���#3�ܚ��1W)�J)����:�Μ��[�
.\�&�Az?6���bV�\�@�H�w������Q������0ti�ed�6� �T�mʯ)�(��vb4��id͐�Bɬ@�q/o�t�/�O4�����Y/:��'EBf��Vr �
@�ѵ��C"Lp�tFB�-5��8L}���I5t2kzJR��8�t��B=��h�Ol�i��kܔ�R��_�'������U�l�h�r�y�GjR�-���-(2'�Nb�%��y��fF����o|cc[&~���.L��,(���3GxB�3�	=cB��3v-t�e����Řh`��BLv�I&�`6vc|��(<���e}07dJ�K�]���5&n|�^r������g�[���1�� "�z�����G�:�����}S�(d��@0;����-�­��4��3�Y.&'%�<E1�Ѹژ	A���e�4��uE���7܀q��9�}ֽ�<t�&�캵����pW2Vw�w��ݛd�E2u�U}{�J.�R!V�������R��u!JN����t��Qc��|膤���	�{���P}ҩ��p@�>n��}��Ō��|H��o���y�.ڗ:l�Q�Di6y���2;��7w�s͉��ޤ���s�#q���mn�H$Ḭ�����PpO��©�,���`	��1�N��:�v�m��N���Hف��@X�Kɩv���*�P���t8�������%d����Ŧ
�{;w����d<�%Ki�G!�/����ɻxmG����/���������J�P◂3���k�$�5�U%��.'Slk/���/\�W���V7�����<�/�yC&9��Q ���Ή(�S������@6���d�fxi�L��F(��c[���s/[��]#��?L~5��O��X-�d9��,�����\f�Ӕ�,9J�S]A#A`����1�ֲP2�������L�?��`u�Vz�DlV�f�{ �N5�^/'!��G(�2�P���q+�)i���%$.byų�vn��{����.�(坫�@s�A�%5pWrL��Q8������=�<~"�Y^o�\����m���e��_�)��%d�ڻ52ɪ�5_5-@?A���*m]�?��'�m_ՉNdΫQ���
j{ԕ܅$L"I�V3aX��&
CC�zF)��JI,�VjBpkf�A$6$��=W^$�h ��x^u��;��D���ܳ�����xd���@~����H�G�KV��z�5W����/D�%Z5=S�F]O�M�p9�*�	p�T�m4���BD��Č��M��p�$�)�5�9��[>�2�wB��4<���-�yYA`��������7t����<un�ǹL��V�&�!��Z�f'����{]��f~���}U=��K/�'�N����f�t:��P�����Ix	԰7�>B��������f�o��@���[Wy��%���i�)��ls��;�-����CZǿ�`3�VvT���)�Vs?�AT��?�;�Z�q���5I��D{�4;�w"�����R �J��b,��bd���v�)�U�*^�' �j(������+0]ܵ��6xt��7����M�AX�%E��rf�ه=�ƣ�㫯���;������^�\�y��]�)����U����m�zt�t���f������/_=�9��[�y�e��L�6'�x� ��F���Q��.W*��ˌc��0�����2%�Y����������V��҅�`X��ez�8�D���7�+D����s��������dn�����\��cu���4#��d�so�,]$ꨰ��߹㐼�c�[�F[���9���v�4�z���B�M��k�p���R��&����
��h�w�(�S��F ��ĸ�	�;j�d�Z�1�	^�v���0��6�ǯ:����py�����ճkA:����;	�W'dM	��^G�`O��3;lhq���U���%��= Ni(;Aj�ҍk^��;T`)�/�Ј��A�Ma����B���[��|�4yח��E�U���[!��m⁂E�B�
H���9��� �؁���hn���i����Baubl���&:s�\��O,���,t��!�eȪt�	��dVȖ��c�+�T��,�Z"#��  =����Sw=��hA�o��|@]G��������<՟9��ݝ��B��J�{
<���!:��1�儔�An�����I*������o!e�&�i���R:�J:�JKT|��^�gPq�1ԇ�6�+=`5�:�^�G�>v�����od���:W牼z�o�����!3$K���n>*������������Cl���c���x^@2��(@�$R�lø�������y�8ݐX7�!���QYMt��ax��O[�p�������qVLp���'@�߻�0��{W����zw84��c��֣Zmy���T�ZQ�=��EFt��3� ��iS!�����ʰ������ ����s�(�	���R�!;y���#�q��ߺY�:�|�S���L�uQ`���9�֊"!ଧt@��'U�@_��U�c>MwU'�8���M�JW��E��"Y�	q�8�񽦸M���5<���t&`�B��gғ�(��)�%���T��3"���r5jԮ��?���]�%�|۷JyD|$��X��R=�B��(��1]y���GU��#71DyQ��BMZ�s�wȓ�n˜MH��<(5�I���Bf��Ǫ�CN�Uն{�T_B<�-�wd�a��������Ǟ>��}��b7f?]�?t��w]���q'�i��w���������o�8ҽy�c���� �$6��ܐyI9��ce�����5��|��4]�z��6�QS���l���h�����!��=�w_��߽�O:WJ��fJ���a��q�Xr|~8̂'h˻��7�p˭7}����j����r_*N��¦K���TxީDߟ�&)[����rZ��m�C+�RLX�U6��|�Jjꀑ��je�2]s����6�Dh�Տ��ƭ��G�ѳ/  ��IDAT�����_'�ґ��I�^�_�3_���� kH(��B(����)'��:>㎏�\�-8m�g��7�J����B���2�T�%���6�U��Ǳ�%��*Fs����13$dz������_Pi�F2��H�1Էe&�>�j����~�����+�;�p�w��z��M����G�o8t�y!��qI���_P�(�m�,c�Ũ~���	c�aL�I��/����N�)�O��P=	�t������甋<���u[A>u��a��]����)ġ���<6ǂ�/��������k���]��8�&��O����ǹ��c7J���&���l)���M���S�T��&����������5f�~`�a��h܃�b8���
ɛ�7eA�f���{����W����4t#��)�|*��nz~�1����ܭ�Ó�?���^��{�<y����<O�f��t}��B�)�P�U�}���&Z=�ٟ�x�M��h��`��r[XF�8��ʀ&m���aU�Nx�@ �t�Ɯ�Ƚ�P|�M����w�������ns�7<��~�9�;ܥe!k���=��T!�<�E�Ay��υ�pz9w��Wc�Z�٪o+�#�ncw��'+�v����S��J,M�Ft!�T�
�>�$�<&h����:�O;+d&���'��\H���_z�r����W�{կ��]�O�������
R���|�\.٠iX��m�������P�
4Ӽ�l"? i���4��fP�Ǔc���}L4!6�1���\�w`/F#�d.݋��_�s�~��Ot���B�����$V1�p�G�8
b��<�v݉�=
��봳�p��_-�Wí�Lu0��r�NvH����M�Si�A�B��ss	����4`m�&dr�t���0�}we���L��&sf|��y��Z~�,4w�hG�y��>������>禛��_�����Gn	�Y*�(� I/�lt�&���g����<��)O(%�t�E��@���	�8H�NV��,�`��A���P l�!D�PG̲⎦�?�+��q��(�=k��x&/��n�s�ݦ��ۑ��|I���C#�^ϡ򈽆Z���y_m��Sue'c�)y�R�ϑ�p���(��ӫ�>�w��KaȪ��[�hj\/D�L^VK��c�azR��v��
�8('5���Ai/��!�a�P@[�	\��l�]
�L`��B�'�N�'-��Eu�po��'����y�c0Z׸�=�ݸE �Mh>`�����fD��{�u�$q�(R�a���v6d(mL6r��S���$���oP_�\�ᕣ��u˫>�ܽ<w�鑧;���ˢ�G�uRS�S�JY`�����K�����sjbu���'S�V�|/�9����6U)�^}���	�VG��@��P�P���i�� �K!t�R]���38ĦqA�#W]f�'�6M@^�� ��e�X'"�̋��+,��s����m;������Ï�����"%�B�E���\s+�]���Nd�(8v����d}&邧n["x���[_(=��[�]�m��&:�:Y�6�ᎉN&(Ԅ�2d��=�`& �/?={OO�JHG����s0D@��d:Q��1G-�뇬�=�fy���#���T8��*�)V�/��5�6���c����GY[���������9��BZ���8+�J�JՕ�`���3��̈́��TI���GV�i����Z����uM{N��zi�Ē��P����v�Mjr-CJ�iE�L��8%�zD�4!�R+�������SE�ŸUH�g A��ܛ�X'��+��"x��3jHմ�l��fW
���/�$�b;#���dY��h3<���uu=�k�s�Vr�߬-�D�S����}��ɾ�T�胕�2�Uɑ�.<3L#\m㾃��h���8����pS�6�U`����}�$�Ŷ�/�I� ,"(K�b�X��ޒ��5���O�>�g�]���w��>����,.������v=�t��6a��1Nx=ht�>�J�t���T\Q�Z'�H���$�_���Zv��mu�a^ИBB�I���j��b���N6�자K1tM@�%X�^�����'=`�N����)�����㵫$��5�26�,��~��G����9��,���4�~�q�jh3	�d���a����"��~-�tW�{�y� �e�Ҋ\�p]��}?X%��\���I�h�-nF�'�����<K�9��U� �'#ciX�LX����Y������V�Ў�^p!�����4 �3�9��4P�j`�1��2 ��3Ƌ��j� �~8�K$-R���K]�_�/���P�4�|*�X��r<,n\}��T��4�LuW�SQۦ��Kyh%*��+�P��jT�����T�_���9a�w 6=���P8��\����8�#���tD�E&����x	����VÌ�[�I�ff�ȕ%m*�)!�4�ZM`��I�TO��9�#�I~A�@6�_��?�z���+~p���L'։j�<�\'�ߖS����i�O�7u����Ju��r��["x=^���n�C�C�&|\ �bf�������W7bC�f���Y���'���ߔ��.��f^$�Ә>xࠫ�'�P��-y��;�<����ʉC'>��:\n�_��	Yy�����6�ḥ�՞}�J<<�Ǫ��{.4j��3�ԑ[�z0˸F����:�N�4ۘE�N/x^ �^���f�D��D@�*���p�`�Rv�C#���zWm?�
Q��3��Ot��B��(ՌZptR�^���x2�@x�M22�ϔ�L��?��wI���h��@6V�vi!jGMD�9B��'=���P=�s}��rLxN\o�>d=}*Џ��/_����B�֫��Sq�Ug�#�}�Qz,nιю��)�� ��}uÖ5N�O�e�]�*mk�aMF��L4 ���*u>�����W���4'�u�eB�����q��'��}��z�����N��\�����Ş�D'�mf�;�&+��L�`lrM-g�?e�&���	q�m�n���PYr+ �,m�6C�uptYB&��Rq����A�8�pg�o�s	N�$s}���RD���8�G�+�>�"-h�E���޿P��>,r��N��+ȯ�:�E���zow��9�z2#��T���A3���0��=�yYO�L�: Owf��X�
��&��b��fC�˅��X�W "�JlGj�Pi�T}R;�%����!��k5�z�`j���זZP+��B�w���I������B��i3�3M��vR���(�R����|���}���81�}\/�mZ&��F,U��6k]�`hs�� 	� �9�"?�����i�>Ÿ{�[H��vȒ��0��� �2'�F�h4�u����کT����I��B�SR�Lj�5JMcV��PRE��5���6x���)@b-ai̍Зp�e�6��5I��\�|Y�O��P�n=&��J��4#��j��m������"�����?W�fmu��|&�1r���M|��7�-i��"����┉:f�h�[�5{8��5l@���^���ɳd�9�k���� 0�x�2uA�%�W2@mG�̓���&HP˻+ݕϨ�}��N�9{/lwɕ��D���U�ʂ6)��(gw����i��L�h�t�
�;�����I�6.��ցd.���k~��X$[�)�bd��$sL�P<�3*S�}��B�z?K��#�?�x�c�����C&�3Ё�soՒ,#s3>I�9�E��TG����(�Hf�h�봂W��H՘�p��A�"I<�e�T���0�����JI��Jbg�=�X{7 ���"y8I������ ڽ�Ɉ��9a&o�1Tu6��*Ѷ�r�m��~���_u=�n��W�Џ��c�񀸫Z�F�p����Mp=�hnfh����o���@���v��M�L�ӨZ�n>�}QPO*<.����P�F�f�$˫j��N�F�U�j�G���]�v6$���_���<�ƻ-l��γ�^�w&W�9�����:,u��!
iȄ&v�t��u]v�%�l�#���Pu�"Mlr�~�I���*��ɺႇ�'�N����#����1�QjZ\�H�Th1- �$��D����5J�)T��8��N5!;�u<w� �� ���s�$�lC�F,�(���|eד^�ARپ�|4�Ԅ�9f�Y�HH�c�����Q�Q���S�@?N]F9c:�R�AVᆐ68F(�S9� ��߷k���_������8����{{Y�z��o���s�4���1��ǵV�'�j����0�H������&'K�E�m
AS5�Qסl��w�d�L��a�󌐇�@oh+��b�����?�o��k���z�]s�w:��ӭƜӆ�3������
!�������yŵ;�a���k��{r&�&P{�!u�FJs&�HV}A`�=ߧ���`�tO/�x!ƒ�W����P�\��;���+�/.:K��$�d~0��M��T.�����$;v��J{;���`��^��Y���@q _zN�_9z���^�Q��|������O��muVc���Vg7Y����并D�2�F��y� �1�� �#`�:L/�N��@]<�ِzo����Ҭ`�fL����"��NR�c�j��T��Jj�����ШP@��j���ay�Y��D�1�$50 �Y��ns��qB~�^���S�9TN2��o]�G�]�DS��v�Z�E����ѡm�Λ�5��d���e�89[�k^ߨ�/<H�Q2	��lĲh.:�պ��>p�%Ͽ���,䍙�q�ɕE�8)�,�9:���-S�+�{�5�~s�v�t�}��?}#�K>+6It���y�R@J��h~>ɩ�9t�)C���)L�-)}��ݦ�^��[�������\2����=�g��Ƴ_�_��5��ƫX��%3
�ք��X|׼����ϛAS�/^�څE"�Zc1�a�>��}���Š	�k�"�=�Z��)���ScL�pU��N+H�H	����5��w�3���m�����b�N��9;h���"��};�أ�7�p��_��ݽ��_���
�[?�>����	���&�KwJy�Bh�|���!���?�B0�gS!J�m�zS� ��������:-�T08�8'k鈕��J&u��6L]��8��H����2K��4��Z�I�r��*%�[��5�K�Wr�� +9D���R���Opf��Q���K��e�f.+��M]�%ӕ5����>#��q,��#FfH��֡����8�.>�Dq�:�s��?W:r��G5���ـ�ΐ�c,9~��ݱc�9O��j���Ͳ~����{��Y��)U��%�:����|��<uy�N�^��V#P�T�3_��4�RZ5ь6k
���D��
��}�ٹ�&Bc(GS��>
����{Ld�_�/�ta��/~���7��{?#���C�h�Do=�KwĲ���CG(�J��b����+v��J������r�����Mݛ Y�\eb���m������w�[��F�@B�4�d������Ǝ��q��1�!��N��c���`���ǈU ,�AH$��Ւz_����z���e��yo�[��{�Wu7J��[�y��<y�� **	5��B��~�;^�=7���^�J�4��@�V����F��Gd��4f#�M�]�o�����d��\��/�/mR���e��g�Tv�x�{c_�'�h�S�w�����]��/�3��_v���Ǜ�wn�9X`���7q������=)^k<�����Z��d�
�b�Z���p��U��ZLՠC4���wݜSp3NV9�?ĄAdWn��C��h���*���	�2����C"`ϟ��e���4Jn����>��R �9��`)�YE̹:�1�2x_O(��� ���L.p�|Y8d�%y�=Dww�c,�M��l(-��[�3�@�ҕ���%n|�w�����'�������7G}!��'��J�o|��x����O<̶�Z��f볟������;of���B[�8�ߠ��Z�JR��i��٫@[0�K�^?a�iaIƝSV���Y�V	�`��L�����
��HH�Ɓ&c�p"���7�]������W� Li	V�V���K��Ψz�����G>b����^�;�ޗ?���t䛧ev�Ѳ��r$*���~���N������C{~��go��ŷ�&�%��y�N̼[c�uc��ͅ8B�$P��tEq�VH�A�����<c� Cއ��E��I�9�tշx�?�gك���/��>��'>�Ϟ��wΟ3vb����u�}�n����`�������Ŀ}���7 *G�rS��.���ئ8����z����@z��#�����}6��>��
4���3@�7��Ʋ�40)xl㚯�LÇA*��<���]��ra24���H��4!��Tqr�6���
�T���?D�-���l����L����گ�W��mMd���L�1�	y��;�i�o��h��ϛ:IQA���5�+s�c���h]$x�a��:sM_M�PI��� 
˽�7��;�x���p��,JW&z��.{�'?�>3:ͮ������h����F����l�=��S�o�>�9�S,閆:j��. ���M�Sm+��a�C^ߏ,�����������������4N8�8��A�������K����K��5Ta`�@� �$Su,kh����j�e;&��S�_�N�?v�)ֹi�o��3����O�g>�_��=���N��N��������'����/bp�e�~�<��.���>;|�3��N���d�L��!�Xa�8��g���	�f�m��E,�#��"7���H,W%�7�Ш��R�Rfy�l�έ&c95�e�c�3ށ���;X��w�11�D�j������>�E�oa3?�c������~�7���w�ܛ����#��^���(�4Y��ڎ�<%V0z}�,f�.W��
a��<��(��2�󤵹��*:��X��,X�I�:��оÜ�M2LsCj�I���{����[ ��l'diE��R�On�ک�`i��;�+~	�s�$���#�jB�n�U%�Y���yo��{ȳ�ɻ;g�qմ"�m3ݸ�}��(���Q�'�I�ſ��b;ϳ]�y���C^2Ӌ���[��/=���ҿX��kwG�k
�n�&J0m�;'�}A��;^Kk�ͨ��;8d�Z� �o��ﱷ����_��V\�̭��8���$� �@���-4W����9+es��4N�.�j�B�^�rg�7�����0���f�_}�{�^����E���1��+�C�_����L�{��^�i�͵��*N}�߭�0�栍�v��ճ�ϼ�f^W{O��H&��*���^ͥ��f�>c�Z�,r���\SJ�qV~���ۯ|�����r���������X�=2ݩ=�+�&牒qYL{����D�>=��a-�Y�)s��{T�q��9���-k2���b�BB�,nK��;�0ud���O
�Y-TS�'Jo�T�^�Yg�?6/;Էv�J�ؼ��0�À%��|���[���4N��ļRv�p��}��vXs!zX���+��}����ȟ	%x��FiTΟAз`ʒ��i�ڢ,_���M�����\W��Ԯ�SV�����sy�~��0�L[�7J�r��pۈ�$�`P�bK,x�%}��k)Dm���6`��]�%`�,$�@!7�@|��(ʩ>�z�?z�`h/l#0?v��g�U�����ʰ|��n������������,[+�e��"I��{م/?{�[�2��bwTV�ȍ���]�c�G��>�8� p�e�gƲ���"��$�k�'�Șr�_d�Wc�}�v����ǟ�Ɲ瞗�=��r<bk����FK�z�dGZ%f���&�N�U���٥93TL~����-aZ)��s��n9��$�53�$���Y��A��b�����a�������3��1P/�B)-&UL��D�;�ƙ��#�8�����9���-~�Q�"�EQIHbg��Zr�GƜ�V�[��C]Lú� �e�To�cܝu�bH{��J��,o��o���k^{_X5ܷ��Ե��3��k�~�Ϧ����~JTh�Ts�獗lg� 	^/����ݕ�� )��9�c�+ZZ�T���z��Ck=����b/�ѕ�����Zˊ|���l��{&�ٸ��J��㞠d2��v���1�.��d
���\F�a���Rn��=�s��@�=����K�7��$pA�0[�yf�秺`2�Y��lg���@�'U�@�}��E��jʎ1���A>��,�ɐm��c���ʭ
�n���:ҷ;��������C`^�!��8�8�4m\Tc�h�,U3��%��}^��QGی�����R����mݳQ�����8��L�Lt �Z1/��8x��}V�.��0V�1{���l�Ճ"t|	��U��	ZN9�#�!5FK�}���� ��\L��+Mc^�^���t�ya�3ߘ�G9�N,C|�{>�w�{B���S�!�4$�`��i�.�0#�=�Tci��Р��>��o��h���d��ss_�j����!�Nc�^�Ǆ*��^Ɇ|<x��h8%:-Z�Hz��$`��c�'��F+�:��������%�7z�-p�Zb8�K����
E��\jN���$w��b��L[qQ�5��ي"MQ4K��oc��W�Ǐ�	���j�˸T��K��;���e�~kK,�����U����5:R1�#vhq���v�� �h� ���h���%�"���'U#���_�Ą^���!�T�c�}M}�ha�Hrd��ᙻ7mPV��1��Y<x��Q �U]B�pHȚ��������o2� � j��*�&����e��. )`�Sm\���fX��qbڗ�!
`1��6�rJ��=�7Ti��<G?�Z �V��(�?f��qq�r(Ю��!�����ފ:�Ee9 fUVƃz�+�=���3�~��@�Ԕ����u��e��e��ᬱ�Ji�%+�+HP���%��I�Ӹmt����`��aB�gޡ��_$�����9��a<K�(����Gh�?xA�E�<�ن���>h^��AH'��p�|@zm$��e{�����=��-F���J���q��ߴ�d\��3Z�n��>
`�b����%��>X94M,q!(�>��8m�����7����ZV�䗵HBMֲ�۠�s�U�\<�0O)&���b�9�u���1w_h����ǧ����>�� � �O��${�"r�u^p����Ֆ�O��4�������������DLh��&�d~�b�m���Uc���B�f���7�2�$�£aĬ}E`�tJE!�P� ����!]*��G<T�x��9[WVW�sN���+�C��ٴ,��
�Jׯ ��l�Q�μ�˿:�;{�g��@�h�vwoB���w�x���F��@�o[�kK���営eL�G�x���#����"t8L?j(�����twy
��J�eY����X�h��7�(;�	����+qwo�M��~Q��eߞ|+�Y�!}s���Aa��4i�,[�* k��4��*�9n�4�-���<�IӁ ?(�B;��(�$Ovz��ؙ*��t����<g� �3Zw \�EF4��
dR�~�mG�f�43t�320��2ђ�s�=l�v����y��A�9@�R�KƛN�Y��z�?C:�.��r��߻��JQ���?a�{�&�ڒLV+7��>�:l��	q��Dx�5�D��G'�������nO�[�1ų��A#�{~߽3)TQ�����v�����{z�2�~:T�v������1�����h�K:�h@�g��ut(�k�0*�/8{X�#x�[�+P;uߘ�E��q��U��݅�#dzB�A�]��L��	�-��!�\�59r�@�+�1�7�3}8����rMXt6��.����[�0� J�Ql�3

v當��,�<�(����(�V�/ۅ��Yd�|�e�LYкd}p��F@F�D셵XBTI����KM%vl���hD�MJ�:x#<��d��ڥ�	^x����ĭo#MʥQU�P̀%���i�q~Xk�1��T�׈J ��/���9�� .c��$�����%S��)�U���Z}�.kh���{�!����~���>�c?z�vbq�l����Re؀��z=�gV�Q�1��=����p6���-��,c��&ƚ����QMP��G!�=�-�m���3�A�'H**@F�#M���!��j��ss�EԌ�4��dΤZ�]{-�5NSH~h��1pz5S�� i�x�;|�����;��� 	>J�d\��� �Bo��א�j�]��X�s�*)2zJ����p�>��c�,���%Y��]���!�u�ȌǛ ������t�T�HQQ٘�pp;���j�I�r���:��X'<1�5�2�򸛱hyC�i�8�W��]����Џh<��"�tς�
��Z����<lY����3׶�2�M&f�zZT�I��8�Z��JqD��n��]������o�Z�Ә6�	��?k��Vi���<ϸ�f�*9I��Eˁ��4�c�Q)'�d�$&0�)�T�+�$�bf�hs�z��1w���9�S�$�0A�����v�k���)�����l�{vD�dل�t�ˁ�4�p��o��ν�3�eE��x��pr�a/ͻ��<���&$�t
�܂͎g�!zW��S���M�C�w0� �{Hp��~�#�c�H�G��ڇju���mA:�X��.rex\��8�ň�:@�D�;�r�-.6/2������xKg�BjBƪ2�������>�*~i?�?�Xs&F{��n���;�E���J�zE\���؂��U�����=�R�y���wqh�Sx���	�X�s��K�%6a��p��PO�������CE�L�i�K��0V>	��1S�f~��Z�h�s5i~�o��,�L��F��Q������?�����K���hN�d2'�F��L�W�Z4t�9Dp�RU4���b�!���Ȑ�i\z��g��C��o��,�N����X��5��2����T� ����9�S�ὄ�v�hh'ád�AĚ��e(����	F�,k$,���
AO�Aܼ("���҆��8V?/#Qk�̍�,���z�$_5��Xw�R���W�U��N�o�e�}��N�ޜ��`Sv�.�;o���_� P��:��(ݳ��5bS~wW��@"����K���W���Ԉٻ�/�m��%)�T�k�uq&��y�ţIL���k]�a�S(�[&�����G�����ϟC�k%��$�\s����6xD�3�f�<,I�'5�E~��y9��q�a��LX��Yӥ�@x��7�UC��d`��C��@ډ
����d�)�G�wlf�֣	Z#��/p�Nz�3M�T��@ͣ��xB����Q�� �6��K�c�,}�
�l��_�<�Wz��ޕmE��{�f�x:��=�>�0I�rd������lf�!s�F���8��7ƒx��,��=�1�i] �R�!�Mҍ�i�W�U{�Ca��3 W�|	�y��V�0�>ksp�C?�<	lo��L�����e <��b՘�u�.��1EQ����5�WV����4�/!_o3��ƃ�-z6��R<V|��!��(�c��-|�t���\^�0��+�`��ey�b�U��lk�/}Ù��D�#�,��:�^�{��c�Bc5�:�>����{:L=���^`�:�!�2w����1Zn�!��~�R��8m)\pw����BWh��ɪ�ReY���W*���鈑��P�&/�C�j.�a��0�n/D�<��s
��9�	��Ef�U޽��j<�#]��ɺ�~�|�L�Y��?��k\�i)��a�����ҳ���C̠��D3�ǈD)	j�O�F�s���z	K�G����o�W�]n�!��c�����UZ���O�6v-j�*�
��dGa��!�K,��K�"�i���p̼��-�;�m5B=��n�Pj��6���|�	���&@�$I��x�Qs4fK��J �K��E�K��\�=�h��{ߪ9΂c@H^�.F~&I�2u(d��/1���" K����D�[��~��X-ɢ>�
�2�]Z�cU�"���8^��T�~�y�ʕ��?[U����Z��x��֌�+@z<�`�< C<��5YP���>+(k��L/�c�6v'p9F�n)�0F�I"�5���iY��d���t"ƓI�7#K�p�Z�Y���S�nF�R��U�<"70d�%�V��|n[[�7��I�@�̌��}�?����M�eNV�![z����3)�*����H����߸
*&���2�i��c�����|#Ϭ�3����$P��rC!���E�� ��K.N���B�-Q�Wh�K��v0ۜ�u��4�NyD����0� �c��#�7�����PY}��Q��B���(� ��qL�r�5_B�32qFv�E\O��ȶ:�)�0�"A���U'���`���iRY�aTeSj�TL�Xf�~QM���D'�%����&D���$�������Ғ�m�d	w�}��V|v|��g�(7��~,��o��s_;�(+%�r��c����[�R2���'^��[����q�\%���d�KT�E����f&��o	�ʸ*Y7�lK��G�L�/���ɯ�ˏ��i�ֵ�H1!�L2˝�t�U��z����/mn<�'����Y��5.��!���9Ů��m��v�:��A�;���Is6�2�/Y1�Z8MsR�g�t�Zq�{_�l�a=��;�}v��t�_�D5��ܟ>w#�޺g�?�1�.mt��� ^^U1��������ا���W���߹Q^Ȅ�UgB!�V�� ��3�X�=�R4J�i&h/� +#]�HvX8
��_K;�w�u�׼8i�S	�!��i~>�kGe�k�8��n��S�'�v�i9(�l���%k4�ܴ������X�����vv>�������W�g�xy`���,rz�~��"6�w�t��_�NvbA�����kk�mΘ�&�Z
�|����ܸ���q�(:�S��Fq�g�O?�/o_��[��J��t�²�0�e�1�E������1~�i;ׯ�>��x����'�%�:�>�����d$TH�	$X��!��zP(�F�N�
Xԅ,hѲ�)iI��in���s�	��q���}�<GJ����oX68s��_/�ʼL��U=��;ӽ�?�7��ջ���^��yȄ2�W��[���S��y������{_GE����w������<��T���ǐJ_��Bp_ �jN~t<&i��w% �b����[���4�v㻇�H�{<�𽧶���{T~����o~�����7�b4�L�����sT�������?~����J��$zG,Ϟ�q�a�۳�k�J��R�~K�_nK�>`�k���½�`���M�m�A�lߏXF���Y��=Jhm����۞p(h)�%�>������:+�e�va���^{����{�{﻿�T�C,�ܿ,gu�gQ�������ϫ�7������ɩ�[wd��r�)S��S�U�daǛ�8��ET2/�^�]i!Xu+i+�e,�����$-:��%S[g����>�;��G>�����m8.ϰ2��	u-ǿ�m9T��w�1��/5�wn�f�q�;��~��`���*�v��;���� ��#+�o*
V���ƀhʝD�C�S�pw@N���w�Ue�MM����!��k7 \"8�'�8��a�#�!����o/YyU C���H['�p,E���3R�R��`j�q6���r��_۽�Dy��co�ܺ�]��I��KD�7�V�������>��>�;��yj��7Pߓ���2�8��}�&/��* ���!~s�&�Xf��!K�~�����)���~�4Qi��.5F��#���-8]��}�aw3�K%�M��)�r�nb��,��H=���G��7>���c/?����On���̄���Z���U�p���w����=����u�;k��὿^q�����\i�"�0v���d��8��q��C#��4��p0j2�)>p>ǚ����p�ui��B�L�/�bђ�7)�G�,���YhRK�TO��53�������������g�u|�ƫ��(E�	Ne@�)�2�W��Q�x��]�;�r���`3�K�_���9���3���R��=ԁ�w�5�RP�,ZB]�pKkB)�����TOX S�@�L9��-����qXV��x�_�^�YUp�gN�躈���N�u�o��ON����e�Ϟ��={���B��YCc|�����9;	<��>h��e:�����x��_��?�����ɯ������=���[�:����cg����2�3�r�8�P-��� �e�� �R�0�,���	>5���c� �&�����^
S0 ����6(�0�1�G��ّ-�5~>����}��NX��L�ܯ�.G#6~y8~�����+G׾��ɍg.ƻg����V/$3�~e̦7���y�ޕ�*�_\/��&޼돢d�L'ꤑ]��� @����Q_i�.����@����Y9!y� C��]Ƒ,�i�	]ݐFƀ�	b$�淄m��jx�1	�OÒ>;�=���pPZ�����]m�b qw^M������'�b����:��O|o��o.&�,���M����P���ݽ��"7������������Dot؛x�;3Ͳ^/Is���q��X'���~R��8AK`R: e����r(u�4X���zdi
.�\Hd��q���9SP�c��1 m��Ŀ]mz{�1p2�YR�I��!�n����;X�T�gh�߾G�����<=��̧';O�oo���/�#�ܻy����O	 ��^5���m�v�F�}��}+�i>�W�wџo�ѝi$�U5.�/i5�vX1@���##W�qP�Ȉe���ڗ�j�IҐ��,Z���q���~2c�JKc���+������.��y]���o���yV<*�L
n��lzs;7��Ve�W�껮���M���s�"]-���j;��D��⽇q����,�	�Q1��5�j���7޼>������_���_t���qF�n�Nb����Hg�;F��V1��$�V9WI�e�U�	�G�JW�LI�2��j�Dne��అ��(��,xa�n�n'���NQ��"KLj�Op?e�B�O����������C'�s��O�Ԉ�0]^*ˣ�d|������>�~�o�{W^����`/SZ��v�v��5�<��r|�o���a��Ȭs�C ��=���`ŕJ�c|�ki��:��\g�=a��ʥ�IX����"U��h��9ed�*��Ov+��-��G�E^�5l�Q	��rd�_�uj���h���-S3�}�M�x(F�2�ݾ��S��M6��]���sB�AtH3�j�_�u�o����c�K��4�����譟�XF
 �m����R�*/!(PGѹ���2J���

�)��^
���e����b
j���R��hb@���Tl�a	~JX�ܛ�cW��Η®���j@+���@�@����Z��p�b�d��]@u��9+����O]�z��{�S�w��G���o}�0U�F���ߎ9Y��׊��BlM��o��<V�ݵ��:iGUe��1C,.�L�n���O����[�{��o��{Rc��g����s2�����z?;����?7��V����mWt�krw�n,u���-���U��1���Mc^��ED�������z%�{~sZ���$x8�l���%JR��p\7T5�:��>�=��-�����ɩ�;Ig:H����b^�Z5�����]n�HX`T�P0���e"�7�6�"*�"� \X�5����p�!9Y܁cϷ�$2����T�Y#� 'ŝ?	��n��<�'�WLF7�G;����]M C���0�c��ɷ�{������������׭�]������*���%���ّc���� �z��md�(0#�����ѷ r�\O��sJ���G@�?�k��.KS}��1fd��ȏ�`���.����Z���U�1��{����b��v6�X�r+�@C>e�R>>3|�K#��y]We��5��7yu=*nU��'���	Ulr�%���[4��]�v���X���m�����rq��Ue���#��T�=O5h�BƦ�����YF�Q`�]��GU���^v���o)WvA�t�G��P�;v@�=�3K�Ͷ�"����_���^����������;�u�;@BX*Um\~���ˇ���N%�g����n��� ��B��@{��:G�F9�%|�a9����>1 ������!�����m�%9 \-M09��U�0O��h �F�D>u�<���\d�,{3i%\���s-��ɲ��N_9�촑�Ğ6��_Z��d�NW���Q����äxm��_���{[zwo#ۿ�@&��Dv�-%ЋE�@�2(�o�J�Z�Ю	Gg�E�K�ƨ��o�~.f�Ep���m��E�k����9j��qnU��X��T�8K�1Z�8R����c�)�7%k\�yC���K���;wO��|��72[�.6)d���`Xä��l�@F���%��\��>UY���>r��2jt�����-h�`Qq�Q�u��@����}Ȯ���;>�HO��C��ɨ�v�N�9ƺ8�  ��*`��/?���V���k�t����ɫ&ן���N�66J�[��t�Qh��f׼��SeW<)-��Aħ�Lj��v�"� ��K|`��,��M�If�=�dǱq���م�K^�	W,Voۿ������ ��1o>$;a�쌳����[ݽ������sI��&�R	�2�-	���/�6ѭ�<����;�������^�j2|	�D�ۑC��D, &s�*��tdf�Gr�ͯ�hf�ǡ�	m���M�����������X.4�
��Qj%���� �AJN�!s�h�6y�����]��l�M	�J��+<ͽ?s�`�Q,+�u(�̐�h*ˋ�5:�|�OfHR�[w����.ز޶�k_��Ο��^�I�et�4ÉT(U��io�6.~�Z��{)6+\Mؖ7�sq��T=vV��(������D����Vz���̅����� �0����cV�DP �yd�)���R��)s>��|g:�q��u��)a��&XJZiJ�c���*u�]M�p(Ԅ�zE*Gר��%�������ӹ�E��_��C�2�?����]�]�s�/T�R��bM��w*���kB�#���RU�U�q���.���`8�\���WI�2���z�E��{�SK�^ p����ȍ$�!�'C�q3�{�x���H%���k�dT�X�T�C{ul���� ����h
luy��V:��3���\o�]�6x����Mk۾�,9�������Ls�5 |�������9�� J
n��Vơ��9�q�x`Kf�:1�u���W�jG�����J7���Z��y�Y�{{��pǔ[8	��&�=)�(8��̷��j�R��8��K��Or����<�t��*2#�?M+����}�GT��������/>�搋nR�ۯg/���K)���������V�ԉ��C쟗�����W:���5at���ں-g,�a�|�5+���=F�S�/�XM��v��k(��dQ���E`v�I�w@m������!�b��zz��Ŋ�~�����Q}|5�ٶ�a��X#`�6qԩ��@�-7v8��ߎ�����E����S༌�]P��m��qh{A��ޚ�TKn (�ޅmF�z��q���5�&�mp� �͜�PK�E�*�������L�P���K��J��"��~�GL�-V�{Ԓ���L�4��گĆ�rc:���)9s���1����dNtnL;3��s�)����l��z����?^���_ږbѬ\M���_�J�����3����v�6�֊�6�y}^Ô���q�l�Qu��/1��O�~/�$���Ф�Κ�����> ��,�5ˣp΅��`��R��ڊ���hR�s�E�h�1��%�︈ ��^������WW���I�+�]���9z��3v�im���yn�"Z�_ʦj��aS�Ԓ�T�~3������������ʆD�P��6W��3O�H���&u4s�|�J��B�͛��x�<ޭXKj�c�ca� ^�h�hj<�>��r��n�~�`.x��2wi���`�+�������~����>`�u��W�v�5C��Rf`6�6l�6We�c�$H.}ۿ��QtZRoI�l�z4*����,M��h�=.�y1�틷a�E���D`�����������=�4q�(��v�:_J��7��Ŭ-�O�&[�>��ŋ���R�0LRJ	�V��K�l�aS��+P�)�I����
t.�M�r��H[l�S��]�7os�ǁ�$��<aY�+�}��I�����/M4F�o.T��<:�z:)/f�Ӛ�%��t�1o4�u;K���Ͼ�+�ijn�������$��̜��c��qN�c4��iOd��1d���[̚�׸R�s%�U���I`�8	��(mfP��w��vЄ�{���l�HګlkiG��mٴ�7�]p�~w�6]m6��^���Dp�j��U���L3bZB��?����U}�o�-�]��͎�a^��L;AͿ�:pn��m�gP�7��`���,�_��@�QQ����.2���ϫ�JZ'{xiOG/o����ےLV�����8M�L1�J^z��cZ��+�6NT�%Bt4�l�c~b����h��a�md���cl֫�C���?��S9\͑��0��dyB�Hd���sX&��v�D���` s��p��j3���U���j>�[��"�3��Ϩ�Qp-��PjZEI`U�͚��L�����$r����8����V̕�@9�%6���+?�bF��ʝ������!( W�M�L�e�N�»q�����^��Bu8��2�/��k�*�xX�/	&�Q\����6)�K����D4i�hp����l�FRu�%�%2?i9}v, -]J'2w�T� ��br�Z?tQ�Vx�9��7g�	~�0�c�G]u�Ā��b�����h�`M�{@�V�X�	�n4h{�*v��g�,�`�!�X��p+�չ� ���x[���s��a�R=C"iv`��8�Zj�QǷ����yƙ,}]6&������P�2��L@�*:����҄]����p%���+mu��F#b3�����`Yɰ/�]��ӅJ37�h%�\i
�wz����1����������٬Fۼ��;��*'q���ڍkw��!�3�4��cJ���O��k�ّ�}�8��*����}�1I���QR�qD�ؑ 9.4�}��OK�^�����ĸ���@�L��n��T�̓;>'='���xC���-x�֍^��� id`�AX)\pJX6���,} }Ɂ�bEMx��+�Ry�T���q�P~�]��v}=!B\���ߕ�m�E��q� NQt��m{�p@�h��ɾl
�}+��� ����%�0, �T�>!d����ax�[ ���a�2X�lF���9��ӣ ��'x\0aHF�5@Z���7��n�S	D^斸F~�Ȋ<�_22*N&^�d �]����&�uw,�V[L]�g��ǑL�Jeff����`��s̉0��v�[����k1���2�+T�, �.H���~�,��K�V~H�}a�T"�TFeb'i�dbc#�i)J$X�.0���	Iw��l��'.��r�$+��)L_XW"7A��d^��h,�F�q�nBp֕�>�X
�@��"��#�Q��I�� �;�b�$xi
�(B�Bt��*�����1y��h��ҕ§��U�]B,��*�c�n?ﭟy����tw�̍~om�U �¥%1hyV�1��	��:�*ƪi�rL"�0��\D��4��@��� WҎ�������iP�K��b�.���)�8`�*) O�,BWX5�I����y=��} �� �B$V��%�;�@S���t|�x|�|1ھ���M ��r��Zk��;�e!-�Z��[_��&iw?�:���>@Ņ}Z���B���%�4��Y�
@�C�%�#�/�ێ��D;�h}�$/V��J#pT��U�����{h)�8H���X0�gx� K ����{�Z@4�v���:$�2��˫�R��RFì����t5�u��^2��_i�gn9��3����%��A�~�LGE���F����.y���$i����̃��I�o���f�s*�N+�����ΰL�p_�G[��dL��Qv����J`�Ofui>�Po
�xZ�`\�2q�@r�X� ���WY1�����EҸ���>�
,N��X�#p_s��̦��$y�ߋ�܏�m��'�b2� ��R�GQ%,����Y sՀ�%$�>%&�5ʩ��DeS� ��-��B>)��������(��(zX��2v*`U��P�
,��eZ` =ގC��؋R@9 �6���'��[�J�F��|zz�ͥa��T�;���p�~̚�X��,��Jk�*6�UnDU .E��.p�8Iʤ{������8w߇ַ.������g���0ʳ(1�4 �I�M�2�;MJ.
�QՉ�+�K2zh�����f�0�;
0�',�q�[�cY��NR�	B�}up\���$��%"�+�O��U�!��L���磊����}�����ߖ�]�66���x*�Y�x@�D�Z�(���/�S�h��_�=�h�� �Σ��sX�k%NxN��i�dub�]8�9<}��o���s�)��߳��4��*��$��J��O�JL���o+�ш��,���G{[�;�|]���w�����j���[af[ݸ����V�*3�^�u�s�w�sBv���mM�(�% �2,s��J�:`Y�� )�~pwGԖ��ci�!�� ��b�Y#Μ� ���3ueA�ߖ!<S���a�FA�)��:�(��jڂf�%�` �%������xxi�}�5��ƃ���T��J�U�'T%�F�#�f���H^9�v>u>��ʖ�zlڑv�X���&��{ �\z���`?���}��Km�ۤuN��=bwn�Ι�������y}��W���ox֋{7'٫o��ﻮ�����V���պ�����
����f��s44�&�w�җN�{�{{����w��z�;}�
���jr	����{d��u�r*1�`���N�&�8Zg�q �RQpVRw�m���!�^�uu/�y0]$b��]WH�`�C���o����+��5n�\A��p٨�����O��n��U8���G,Eb�8
����
2w�'�����78�U�>s��O.�E����q�����'ա��tQ�L�ż�!��N�P9�r�2!���B��裾N�jy��� ����!����R�߸��ذ�ъ�:U��br�J������=2�]S���L�O�����ow=D8b�2�]���_�����~��y���rP�#�E��q����e�7��L��C'��9`����9ǵ=�V�j�M��
���`����[1�X��ļ_Q�n'�;�W���Ͽv��?��<��*�;e����~�r؎�^�R�J�I��^L��?���蝛������{��3ᕌ��ꈠ�źD�ͦQ�"f
Г\�~&��
H����O�P�d"T�"qK)ٲ���7/�Ǻ[����`H4+Dr=���7��O/��:��'�8�A+3��4�i�Nja*H����_T<���~�N����0޺������ō�_��s|g�s����g%�Hi(�!M�}��&�� !�7��Z���/:�k���$h��Bf}��q�E���֮6$|v+��t�P?D�,��邂��$�����1�7P�m ����-����4��/�;�r|��Ӭq7�T)xrZ�t�Ι���̥�}����p�{�e�ԝͷ�\� �,��)�`��cVIڷ�[WM��vщa���x:/P������1��|�ܡ���>��;��F4�Zz�ڥ��hlJ�3垨���N�������LR���W�b�[XQ����	��n9Fg�������������k���5�w����/�{kq�*J����L/,��Dc��^���� �'�
���+`l0Z�`*��
������V�3V�3���19�`1�-��
�V�~�P'��҉�-Â7�J�X�`��[A����oa�@�ف�9"������go~z�y�c��ͫ7��6�7���j�ׁ��kc�s6��t���������I�����+�;����J$\�����-J���\�_�	�� �8r\�sĎGӔ ��6�jΖ��^{_P��v'^�0����lqh�
B������&Y�I�Ci�ܹ����X�{����˽���x���B���8��9���x�%YWo'�d��p�1�e�?g��O�_��C�g�u���w�GG���M���C�De�yn������Vz�:��@�9OY�H���w��1A�T���t�Đ�����{���pQ�G�Je�`$4��"��~�X�U�Ir_z�{�i��ộ�~tR�6�Fof�tv�ы���g����ŗ�Ʌ���q�փ;d_�g��J䖃FNP��)��M�F+U���eV:Q3q�[(2n�IW�s9�������v�GZz�+���:s+8�ОR5!�Y�o)�L7�}u�./u���3�۟P���SN�����5,7A�2�����,�S?�=������S�����N��i���>�l�
,�a��e�n^�X'����#1��S�6���¹f�D�'��$���9^�q��؀���4��S{�elvp�2(^.
}�쩩лwO��=�������G��U6}��t���y]du���������%��w�����;���%��k%�������E��	3hŊ���@�A��*�#W͜@�������6�;�����P�I�٧����v�-��v�Z��K�6�%�~����m~�������T���Qg�*��C[K�?���Ҏe�E�P�d�?V�&!�w�N��>�����}v����s?zK��v��i�%�A�8g�q`����IaD�^Ϻ���'ƣ�C��n��R g{_�!Z�[lE�[8�̸�*�Y'�U�ޭs���x��������]}o�w�>�".1��H�vi�?�nl�n��]�޹�~�쬿��T�ߵ|�	�+�xb�0
G;�����˹s���rr��;���]7gۺ���V���7�q���T�Cۿ�H&�r�u�N��o��3�t����rp�M�p��&/�(0�4�K�h��#kg���":w�k�7.<��;f�f)Zϊ������s����Lt�7+�ߓn�M���n�c��uo=�x˩S�F4�gk�w��h��Χ�ʽ��( �II�#�@���t}-~�z®����O�����7��ߘ��1XZ@��n�˨ <>�sJ�s��5-��IPrl�;.I�_��>�yf�U��� �v��=}ǫ~��ީO=/�<���:���N��sAx���8��J�3���J���B���M��(���`��=���?�3�'��}[.ߠ�����7b�X�` w|'�
�t�i��^;�}�x[q�m(z-�([(qw#6���*b�M��y��o}���O��������v���K�������%CF7Ez�s:9}���x�\n^ء�̹���m�Q1�|p�e�u��勼=&��5,,�V���N��l}���K�����}����Gw�<;�/��^�����d��m~�'�������C�G�~��[�*M�]�Ե~�*Y9+�����������Nf���[��g����1�v|�L�~o��O�����_~�ՖF��d�CƛW`ø�|�5�sݎ�t����ѯ���}{4�Վz�TIPfuhRv�����.j�ΟI����	.���!;s�@L��ؼx�m?�w�������W��o쌷�E�ƛ��L���n�V[ߎ����b3]�Lְ<Xx�������Q/br-�ܜ�A��=��&	�c�Uc��Ɖe���	!b={����(�3o�(<�֗0��m�}0��Ip%H�X϶zk,��ŧ�c-qR����q� �#Ђ��QZuz��h�v)�C�)H���JӨjPS�B��aq�t;��q�o�o_n=��+[�Ž^�CPK2:�y����.p*�q��8�f�������2S%/b�zeG8&xH�C]������Ë�Kͤ���J��B��ٍ��m
��p�������G>����ᶩi�chD�M)�-�
��*�S�%�T[	��*�GA�eD���bn�y��n_|��hg8��g��O�,��,�*�Ԕ1p0��XZ����*��R~�T4�D�$7;7��&k�nn��κر��L-񠜱���?/}DF̬��v�k����CR�|�a[��cN��j�lSJ+u�����	�|$F�um=����ed'[_r�ƪ��%�B3�R	��:B!�z��ǥ?�It�"�2�}�W�ؓ�b.h8]��Kjɓ�W�7��M����ynoz��v���*r0��4�K�s�39�Do���
�m��.�&fE�X����ݳwt�CX$�J*t�n�d���Zzƪ4l�7!���%��<5��������5n0��[|��o-?�}m����:�a�{P�f���MUMY�M��Ǎ{w�������O��;�}.�q�7���N������`A��p�L(�F�n"��*d��I��!�q*�T�V�{�yԭ}���-T��$+�z��.��N�s���w����K➝r����|���&�'XS�����]���X�Y��mF�ch�#�����Dk�pu�nʐ{+���\l�����`�jR�R]0+0a�Tl�e�;��^>l�7��_Y��tgW���D�[v�rx����ɞ��� u��^�����X��p�a�"���n�݈�1��2�0T�.6�1&�	��uȠV�����v�A�����{����;�Ȣ�e��M!�ft���\��5�VhKႻ+��
����?���LT34��M�PZJ-�2�%3���9
���>�c���_I�ո�w줖E'	�N&�o��$���6��(^C�D�91�?.tT�
���P�A9����_��6/�>l@����e���~�!#dW�1wឫ	��-��O��������N�>,���i��dx�1�Jn0��H\eS���u�xuIi
���˙������W����d׾x!�mTv����;:	��pIg3c/�l=�]庪�{r~�吲R0~c8�ɄO��Dv���p
���U�9,h��8���x�C����a�OY�����33�x���|d9|g0�U�{���W�Cv�ry ~* ��.��vbM�'[G����N
 viIf^m� o�N����/+�
�ۅI�L�H��P��(��� J��y9�����E#�%���F�c��K9�̑��&	��
����}��:�� W�1
3�k���"b��w���^T�̛X��$� ���.�	b\$�K,��=k9�$�eʎ�ӌXgX�8��hj�"?�Q� <p��P�4�Շg�QX�!r6������H�U.��/�,���B�8&ή�M'Muw��յ]B��5G��r~ !������
~�r�tp:��Pr�/ [�={��)r�ׄ������,�z��]$҄$M+�2�~��2A�f��"-j��Q��f6R��n!�&tS��Q����S�4g��}�$MYiU�IY���h��)Kӎ)ƙF(� @:����f�Vi�T��
���{�1�𽠁�:��f�T��RߥKD�8^N�����"��]Ӟי�L���8tN��V�s�f�-y}#i�J�R*{nfŨo����Ys;�"#u�_[�T��;��ʡ1 F�;v���i7����2��_�y�d��3��7�����&�f15�J2j���\��=�Me�1[f��Q��A��l}����1e�����i��b;~
��ϪV���7K8!�Aڟrq�,H6
��AcȤ�.��F?_�<�;e��^���Q3'�4���ف�fˇ@��Ȳ�)QQ5w��'�V�r���-�QIBB�3�z�i��X`h�l_n���NV��������۫O��[㐦L��1+5��N�>d��&,�^��G�;g�E;�Gq���0���y-�ڿsI����cn,���PV�B�=��
��T�G��?�7
���Al���>��H��j'%�Ѓ.�##�V.��cZ�!̈K�
*�^2F�ɩ��
�8�2�����%�qZW��C��..޾,D����t��~P�.�7��
�-)KĽ(gC����b�n}���p\T@���|�����4uH?�B!R�r
��DK	I&����H��W�l�fjRK�gR;�
 j�{�_��d�`+v�0t���`3�����x�!8��lXZ]9�g
٭K�#�4���ZѬ���"e,��ː/	,b�>�tcD*?��(�bͲ)1Q�Kz�g�}��i��^���H"���E���Aj�����4� �J�R�D�X�쀳��&�=��}�0ў[]�Q��\�(	T�xS�1r٣9x>M�n��� "53�;�� o@`�j�p%���Z@cNAj;K]h�pn��n yUs���OI]K�����`� ���$�R��K�&�J;N0�n��:��M�8L>��:0�g'���ۂ�w_�Z��L[��NڬQ8�X�t��gV
���j #�[F&":W�[�$�h�m�,J��
@� z��$\Dv�D��Qܲvc���+�u*AO��@8	�b��d'G���(�17�SM�:c�%��k�obF�M��L-�t��
s�Qh�]�OՋ �cDG-���E��6�	���]��]�{�%i0q��n��?b&/���3�I˔Q,����	�|���B��@?�Ru���R����ODc�1M�u����0��;3"�i�K�P�r"@@���*"S�(:�>|n�>.���Z-�W�@��n�sc-ʬ�F�#�jɝ 8R��*"L�Uk�uӍ)
�QL�)�f56ߖ�[��&��akFC�t_�d�7S�07�Nx�H�}�������x�5蹤`V n��p�S@<u�u� �	�>�:ު2ch<��\��|<�Z��{Ɍ=����Ў{���S�M�lÇ�[Z��l�0$\Q
������3�C8)�b���%JE�& 0T�g2|��]�Y��Cm��0F�hN�B,��^6�#���fuT�Y����[f�B�!@�OC?�Ԅ�*�*;&4�^��d~ X4-9����"�p,�u[L?�q j�	Ҽ|��B���j����{zs������ǿh�45�X�n�@�������7Yе$��ud��T5~ �0�
���an��.������Ba�v�f6�@�TV����V,~TMV��7O��G6�� ���h���<3�L�c�}�ɕ�\It�Y���C:�]iK3��ݰu���Y�a}�h@���$�TWh�0x�3���� U0��g����Q�툿�g��I�$�I�d�	�k�V��42n��rNR��<�^;ڬm%�R+��q��KK<��o�zh1w����g�i���.kA> �R_��ރ���m�&�fhv�P�߈eb���-b	��,����̊�Wv!��|��K�UXL
�P�]2? �kd��צW���4�X/�О=�Ƕ�v�?���n~��e����2)�@Y��i��"����Ooc$jkG�����3S G7`���_�8������^�w\�Ѽ�����^�M#�>:4�!�h� l�"�w���P�2�"]�Ǜ�Ȝ��u8<&Qm�#a�d6L�e����/ms���s�mf������ۯ�,�֭���A�"o?��A�KB È��9a��Y�v#�G���9�j2��R�FNG�LӯI���C�p��`%P�$8v�i���#�f���I��iS3h\�d�a_y(ܞS^�u� FӬ�:G�E�q������^`Z��A6eD�M jU���X�#�m���ld+O���G�����¾d��Ċ���>3���?��J�b���<ʨ�h��3�ܳ�"�1Fy�@�L�4���ߕ��юn�ԇ����"�ń��Tm��Z�Z���J/��EN�q2��o��	�塺2ǐH����
�DW2�P�C�!���jT��E[�bb��߀�M�E�P���7E��E�7�	�V�z5|	�^�v(�wIJ��PV&�:=|1h�R��S.��]�른�W@S3wR�U %�<
.��G��JpQ�Ā!w�ez	^ �U�W8s��a�>�-z�P�%�����A��Өw,�f&��*^�n>$������8q�!H����nL7��MX��XR:���oP��u�5�9X�_Z~��/�J�y>�Etl;�7�1+s� ���>�2?��i���>�+#IZ)�2�eG�(�p����O�
�)m�|9d��I��]��<r6�X�V�8�1������NmX��ξG�h�cS�F�y�&��l��V��+�Z)N�.��uM6�0hϰ*J��#�fS�����J#��� �#�#�C.�"d͖Tt]Y@^�=8Q�"��9�X�0�5TO^��W.��J�<�������_��V�j<��&�A�ڪ����Fb�x}�B���k¨�jx�#(���q�%	�0TR� :�R �-�Hs(�gxf�_�[�L�y�����ݽy���`i���pQ��ś�ڦ�yM9�o%�$
��wR �� ��[F޷�8���MF9���J�.DXZ�A�Wt���&��AlT���4����1��T��%X7M�R0������ߚW胦0�\���3��"Lp�1��ߨV�	 p�d�pyV1
`w'���MX�&�?<4K�4�Ө_�&���ȏ0�	y������d�WQd�E�3�K;u�W��� ~Tʪ\d0c�RV[JzL��%���Q��T�Ci	���qU���`�8[&�	�<�4X��ʹ�x6x��<���{������:`c�v�v5 �	8� �AȤ/>A6rm"ɟLS�#�r�r��>�'
+��	�kj�rQ�ɷf��v!PV\OT�c�1[�TJ�^S�]e�حe~l3�Wm|��m�hK_J{x!�v��Ϗ0x�V�_�Oof��в�b���k��?b��gtU޴bRE:�*y��:_�Xt)V�R��(���cNR��g.�ѽ�*�k������"O��	ǒC���@ܺ�$B����şs��5�(��F�ƨ/��NL(&�G!��P��-	��ZL�@sc��Ǣ2�%�VL4�����;�Ì�5MGm�J3�n	|��z��Ih����
"p'`�7-���C@=j#�M-SB�ZD	l���:=��~�����l�w*}B��c�ǖ���?so&�Q݉����V{w�I�$!	$��4�j`<#c<l��a��6�3����1�ޛ�g�x,l���f��f� 	���꽫k����✈�y3+�*���ԕU�7�7��9�s��`mem��J�F��[�f�<G�[��OʼS�V�u��.<eMPQov2v�S�6��{�Cq�V,�m�z����"!�g���q�(㴅s���,���bY1X�����zU1��z���z�殒n�9�U���,p� �FE[��dX�XQ7������DN���r��+�J �-�-�0����f�(!^`Ǵ|V���Z�S�%(�Ѓ�$,�;ƹ�>�U�۰ТRjN�r�S�AbÊ\��*.W5����J o�=�_2���a�
]-����ߺ����te�����T>��Z��۫��NL�@^�Qs�ĽP�j��1��x����)����g��:��_��4e�V�3�-�Iw�Q?4�8��+�,&_X��q�)+.�q���S�y�Z�#�N{��?���v=��~��Dg)�r���$w�3O4�+$���dճ�W�V-�z�V�9e��S"�z�%�c�6��>��_����!��A6ؾ�8Lj�N�c4,����a�d��z�WM�Q�EE6d��#=�[��+�9�l����w���W\������5{~9S�JC�����^�C;�.?:��������:Lj׆\��/�V����/	��ۻ���[�h0�Q�J�1(�:����$����C�jWi�|���>D3t]+�PCʭ9��!��#Ͼl�[�y9��i��7)��Å��˒$'ҳL�0�p،p��:5c�����$�;�8�
ʏ�7�S�є�*�p�&^�p��+ִ����%����ҏ>��3�m
���= ޽�jBg��k�5���Ϳ����W�[���/���k�̛�L^ZeU���:�<���i����q�	�tc�Q�
����
�a�N-ՙ��������(�Wz)a��U�!S���r�9T}'��ُ���v��}�E/��@wVT��s!�X��A�œ����;�L^�$��e!�ћ�d�U��L���N�bhy����l�T(9���\P��Ȅ�e���g�Vù`�� �)�XBrE�7��-�x��@^��+��oǳ�<
[j����Mv��n#�/�1�}��{�w��]L�-	T\M����Sm����g�~v�8�ּ�x7���q�s0�z�!����h��[�K��9���G���(��:�D=���5�$���)�	���jv�7�K+MO����"��Y@�Y��b-}�#����W��#D/�r��;�߅A]"ӏ*�@��/[G�~s*pDM%?zڙ��=��m߿�R���5��7�?��Q{�:�5�@T�D����Yu�������#^���w�S���̫^���˔�K�WE�4zOnt��x��rH��X�T��rvh����4M��� ��Ԗ,{aJ��#"|_T����h<�B�5��>K�f��߿����o���΅\o��,�����Q ^ԅc��C7?o��w��n�����[g���Zɝ�&�����a����6�M!��~e���c�h����Ms�Mp+G2Zt�	hU`�L�ϟ0h����qn��+����+����W/3v�P7]����s����_4s��߹��&�p~�T#ϥ���+��l?|�G�9y�\8z��I�%�Ʉ��f���7�.I�i��dC�mE��%v�[�p�FmP���#�NVz�h-��$)��gR]}�pZ_�hA[�R�����,t\M�<�g"�"m..�Z�s��鼪%с��S~����T��ɩ9�xW�������������k<c�cN/��M*q Y���;�N�c�ݺ{��P��t�r�p�������vi��D��I����������¼�7�g�o}YX9�+?z����Vr��x5�9�p�����\O@,�0۹.�kuH�r��{'��[�����o��`|Y��q��ņS�a��m�WJ����7_������/��\va�7}����sj�{!?7Ϣj���t��ٗ�#���9p�%���������	��֛)�#�7��q�(�����D��ֹ�#�a�z�8W��8����S�[Q��b��R�M�S^BMO���:�xϹ�?��s�c�^���o|����{����?zͥ���}��Y��C}K�5珪���Je"�Ƀ��֭�ǿ�?z:����k�,�b�|�Z� O��B����"������c���V �C���_��p$�Gő`hPʉB#ORR
�C���tg����YB)}4���"y	[��yʑG��%6�r�|ު��?�[T�/����o�Y�����G��
�"���lԊ(��i����}��T ��k3W{}��*r�Lm9���/�Ŝ x���n�wް��Wwb/@��B�Uu�7x^�}�gO<��u[��Vȗ��+U�S���m}=,2�kPe!����=����i�? $�[FS�]�[+����EY��+sJJ��4�ey��^����Ι�G����W+�ޑ˭o�Sw6m)��
�#��2x�ʛ���Cp�zq�[rA�S�.���<܀I(:�pMR�����ԐFQD�˓��;�u?�
��^�jqJ���$;o�C�dvög=�sn�1U7��}�����3U��J�:��Q3���YT��=�3S��#s�3�[�rר�<w:��w��Y�P�3«2��i�Qe-21�{�0ӧ�m����W��w�F��4k)�5E<�&Cf�B`d�,OtF�)d|k	��� �$|nrZ
cFb$��XL�!��(~drv�Gx̍����zv�O��K+T���Ua1b��ܻ�~��Z���0r�G�:YǄ������l@/O����X����O���ު����5+���VT%X�=���z!,tV�z΄�DF٧�W�{���۫�3�f�� F�;7�u��_�eCz�;z�#�`���C{3�R8��ң u�<k�r��6�b�h!�(2�q�I�Z�<o�o��M7<�})�~;8�ߍe8st9��W�A��;��.��U~�u�v��|����}L}��n~�V���fr %:W9�	�M�,��:�j5�r,�C�������p
���P3�Z�*���ϻ��[Ͽ����|s���u?���]�C������h�l�n�Ѓ�'�Ԋ[{%b��S��i��O1��L�ku�\�S�y��BDq�ڪC��=�M��n�ƈ�3ZT?����/P�"�Fh������;6z�����%̘ΆV�S蕰Q��퐭�尌�*u������'.=��&5����Oj{BVݒ�s��Vsc��R$�Z��W.��Ȗ���1x��Fq��So��b�)6E���H�#�,���;9�4h��2��D\Sd�>杨���v!+�Q��j0�D��9�� �ia�=�%r��'��3���%��N
a�C]���{2�h�s�p���q�Bm�F�8��3���~Q���A����Q`�깷z+��Rz�D���zB�a~ܯF��JX9�9U}��NE㍭ę9�D��*�����w�9\���v^�W&��Λ���:����mt+���]؍�������M� �{�c1�1�l��)4���!��"��a4�"�LT��D�c�j_y�-�4�!���?�ug���D��k�����\��^C<���X[�&l�HD���G�`�ޚ� �$$B? Wk'�r6�QN�Ą�D%��B4����S�F8fFj�|H��-t�J�.@j|����n4q�2�N*��i���h�To�r׃'꾳����4L.��g&�rQ+J�	/ ,�Q��pF���MQ[W�k��U���uU ���H�R�X%�W)�=o�m�8���%-w����)����K���k�a �� E���+z��q	��"���@vS�^ �I`���?5ÐW��u��4(-X[S�8F�zÀt�Q"`�^���.RX<沴��չ��.BJ�L댡Ǥ�2�v2$��Y�¹o6Q�������.gT40�Iϡ�Rq}�3�>���?~,>���5�3ډo��\ox���rÍ�Έ�ҝ'/mu�<����}׿�5��'�J��;��=�5~�&��������*�g��1���{J<�L�w%Q`�:V%���V��9��=�	X��[�[~������WM-�kpbJ�R�AR"�NI�S�e�Խښ60#2U�J�H�ZZ�W���F������d-b��جYW�-=\����)���S��c
+-2�e�)zH~)$�
U)�q�I�4���U)����9=C����֭��6��L�oMw����4���c���}P*�ӏ�N�)�Y��m5�)���8��8��Z J+f���p���X׸Fł�kVǄ�Ђ����ʇ�0�$~h�F����@�P��"'���nI����I�j%q�&�Ҟ��>��'��C3��kH���@g�s�>�i�V7�7���_[�ɱVC3׵�׶6G�k1nDC��1�nsu�����ݭn�A)��,�'XP�d�Ҽ23FHG��I|�B4P�vL�=.	e��^A]�=���rϨ��M9���q���m��}�bW�d�.������ʑ�_k�zbi!"r&�7v�~쑃uݧ�������bŅL+!U����˟�/�˖d]�)��|�R� i)�5�a�*��u����y N^�W���!�_@����w�Xo|���W��|�6�K���]u��G>�q�u��qy~�������:��ڦ��1--���l��d9m�p/x�8erR�p~��+�?T���o��<cYO����FĿ�S���f�~��b��j�a������D�n~�OV���_۽�_�)�g�<g��j�T�F�B!�"�tyTfb(膍ö�4����Xx��=n	�T{I�ƫR�!]�
E���T���T��C��W�z�:�«Xv�_￷�w:��O�Gn�T`�6}�rҒ�(��{2��p�K_Ã�0�Lݗ���*�@�%(@Cǃ4?]VB;�0�a��{I��Ӛ�R���������I�ř�[i���b|�G��[���Ji���i�H�����ɚ�h]{k��G��մ��g��אfA�EKm��l\��f���fn8��9��[�Ԕ�B��>��3�f�(˱?��sSk��ԍ0����r�)Y��1x�$@mb0��dlx��	���Ӹ=T�uƣ�����{��w|�Cg�J�K�+'��/����G�~J��ub���BNC��&2��l6��Tۘ|7k}���b�G5�@SS���X�T�����Xr�{�L`۫2ᝁd��c�Z�����V/���Q<5�;IK���0D٣z�8��^�&��<�ӡj�}�1���O����u����?������G�/��L0[��َ�\KoeA^9;ybW0��a�?���g=�Kר�?��嶜|�V�&��bZ3��}B4%���뵊�����zpr�&��#X�g#��fm-z�`ײַSl�PX`��)�M���k��(@FH!�+��ubDWP�2�R�����v�Ԣ�h�N��=0a˶��ܹ�Q\�kB|�D���A��y��e�vT���� ����:ʘ�!�*�����dc8�|��7�2	�6y�-���u��׼�%�ٟy�[k5�͔�<3z�����U��O!��)4�i��:�YШ�9�ג�g��Y��,��gȰa}����hC?�!�:�&)��z}ʺ��ﬦ_:���������%ݎzI�˪��[�W��`U&a��,me3��j���y1�O솢f�Z?�앨�P)�)	0���Ѯ���������_U�����?P���vs�R{ǴWw��ܹS��>tn�9�}���z�W��&n����޶?lv�KN�,Xܚ���hz�#7�!��#�|�_ 1�*�>�U�O'+;��I������&�q��)��12����q�0�9��;�$���X��;��~������9b�ښ�'[�sL�2�I5�	�2��G ��\w��������SE���&�y���↓�Fə����w:�u�`�1��#�9.l��,8�q)�$�b�Ϥ��,�4��󻇟ܙi;�Ӄ�u���0�SjTv�����T9`ڦ�InF���I5n�Z����Q����u���/���gL��*���?W/�<���L�;�H5(��k�����V`t�1����B�W^���u�����X�Ϝ�W��DD���z&q���D(�+�:w�S{]�x��{���<r%,�۪�������ؙp/�:'�=��3o������aU�ʗ�&�~>V�ǉ��\`aHk������ӌ���{�M�@G.�/j^��p_ᵑ� ���(��ڧX��@֭�O�Ց*8�O�:��rN����'2ӆHSZ�O�Z���Ϛ�+a��ĂXt\��x9�B��W�D�N��0F��l������N��Թq�S��JB�P?���2�P�d�{4�Z�-�`g�9�(�s�]bz
d;�8�������j���3�����m8%�ez�^�.΍X�p���r��9��Hմ�8ok��]3@��fw6�̼L�SL�5&7�e9�O����3�x���X]_*�K)ʸR�X8t7LSW`˥p��R
�� �Bk�RL�@�G�-��J�����������ᷮ|��ߜ���W�C-���σ���O�����6w�������~�8Zeu(�ue̾Dfa�N�$���C��־��n@�(&j��S^y�'k��b[�"� h�?gG	
Л��|�#���e����V�� b/n��V��A�Q���$�@�Թ��_��<�كh] ��D�iÂ���n �(&z��[����φ�4��Z��`�'�~R�A���׈,�`E�փ�!�:ڌ�hE>�+ޅi���<�z��# Sm"#�5�������y0�X������9	���8�a��Sq0�5"(ϻ�g�ڲi}���c��Z��Κ���3Y�	=�����6\���<�I�����b��{A��\QFȮ�5�C@�z�EG��RgG�̈l��fq�'��3'�*0�7}� �	��ʃ@�7廰Җ�4`2N�=���[�^��>��{���>�Jq��������3����~y��5�h���"@I<�VC���A|� !9��\��xP	B�^t����P�LV��8n-���fT4h���C]I.*��y)gO����{Xݽx>���/�9AV}M#��d�ذ�����iŉ�ɩ�O�h�/���k�
�i4�`e�ďW��d|�c��:EA9�@]O�,V���$�'b�+�M��n�.�	���JXB7�<O��5`+���"�)7%U�lV���W��Kt�Q�M,����2*ȡT���8m�f2��N-3>�NC������������J�^ν�$��-xaʁa�"I�G������Y�4���������dier�d�#��U�q�V�D��W�ЊQ��萨5��o�i��X������cU�m�g��s��e��������n�W���lk�5�X
��
f2
���� N�!k$�<X�d0ʹ��=��Ǒ��u�u@��T��8��e��eq	2tT��ZU��l�ęq��YZI��^���M�����D�����VT飥���I�*�l�*��3�~�߼�p�U�7 }�fܮ�rKP(�Qɹ��&7jŞf &�?�4S
8�1V�qc�LMV�����ȚtC�V*��E�ɀ�V�$�.�r�٧�a�:���P���0z�N);�w����SPL���h�#5���}*eH�h�"��\�J�R��5�5���n0�]�X�>]�lw��o{	��M�7��'g8��,��(ܕq�k��^C�8�S��
��X�*����䆪5˴�"�8�}-;SˊSA�:�Y��x�=�п��'`�}�T���{2�7�Z��gn��7�3��ϟ��c�7e�Rt�o�H��E�����u�W�����ŝ��W	��`[M�R[�n.(�l�ױ��H�J�f��L������9�����u�W�A���X��(�H%��=.�!k���I���$q�<�������FY��_:t�J{;c�u7<��ZP}��<{|��=o.�4�O���}��}鉣p�G���νy����<��]�,<��1?��epMk����|/ƲO�fj��{��hF�VC�a�uDfL�Jt��̎O���oj&��3��<K�Z�;um�Pp?�+rhB!�~�����H0��j������r-�G�,y�������5��>�	m�GL�tJYRE2gl�mj��#��S&�B�e{�2�^��^1w36���V5��+�8������>���"��w�8���7��R�{Y{/4�'�����^v��je|>s̆���ס�<ד1E�J��y|�6�_�������o��>�������p?{[^����+�3��]�m�u��c_��x���O�������^|W�`��;j�o�Z�Ǻ���Z)Q�z�A�Y�oZ����V��et��f����\Vg����J�����)�HM��o�.rz=`��n��K���3����u�v"��u��~,�鸺�@�z�>�����\�s�,H����_7���?���?��W�������E��Q~�EQ��M1oG뼉�y�O��ڷY�k,�Z��͌p�n<&�/EU��C4'�i$���p�Z�<�x�fSΧ!H�b�V��l��Ԋ�d����"���6�ߴ0IDW��$On�G���Ic��^�`�u�8zb��ʗ����ڏά���݄Ƌ:�������:\F�8��P����a!_�.�WDi�T�{\�t����B�E3��X,�~|��$H�?��ON�+7��ֹ��������ಇ��l��k�:�0�������C��<3����1�ڛ���０꽿>{�?ߤn||)��]�ϺQt�̡�8e� �6���L� �;�ւޫ5ؓ�`��D-���F�%��Ϊ|�d�ĐRdw��Np�-ED�i�&�����f�ǥ/U��}��&���^qs�3uh�68m�_}���({�Tu��s�9��G?�/>~"­�$�
WA���P[*Jn�-G�I9���7�Xz�V��I6�U2#h��m#�B��Z��4������d��6%Չ_������|{S��N�)0|Z�ӱ��S
�+��,��4%T�MӁ��\7{ �t��6v���DS���LM|��w~���^����'�d�ܥKq�Zj�z���s��1��5��Zq��&�4���f�a(���5��X�q�(�d�"ʆ+i�j��5�W�����߯-�������+��3=4 ng0]�CG%0��I�֟�:r���˷*u�������Nt�\�超���U��E)�����}�$���X�xiC� �Sa�R���p��}���p�AI���!�����U� ��I��_�������,�����+�h�Iܖ�;����q�]ڎ��4mo�{G�c�f՟~�G�RsnG��k}O�iD.��Z����Rt����>/p�Z��t�<���d��(77�i߮�:qֹ~BD<k��<ם�%�#�Y[%O*��+�:!B�պH�����ɽ�甒�4��xm~Î�d�⣠
^+ԯ�������9ʓo�k�<��cz�*
ȳ�������w��� ���v����;�J�c��;t����*I�6	�(�Q�Pq=�լ���K��%�ɕ2���V��i�GFьRΰ��5`�M���l�K���IX����m����<ڽz���Ci:��G6�7���a��E�������~�D��9�yI�����Zvx����rt��_���"L��� �3����B�f��{�y�aE'�=���(DW?�D��=�^�Z/I��&n5x
��VMa��Jh~��Cd(4�`1�v%qk��-�t��.x��Я�6L4c9�S�$Q��o]���'7�����c&M�ێ09��K��(�</�C$͛��;6��H� )!x�'��\���^��5�c����C���f�P��g8�O�3v.9GW��c'�ᅐ�c�Ej��{B��F�5h���n]��b�'�A�Y挈����,k���F}o�+z��ߟ᝻�Rї�������v�3�'AR ��vq^$�=�0/[k���� $�:5����a�lxF)|�I�`-��CM���)[h[aZ����M�a�nb|W�p����l���-W����'���S�k�|YZN�M�5@�E�����+���s�i/�W:���,���iiE,H3��~���H��4����(��Hb~\�0�-W���$Y7���d�Ś���r�q�7�a�Q�
g�)�B�BV9)褓\�b��&���h��y3�:���	L֧��G��h����sb���pq�s"sr1��ć9=֘�9
��;�?j33Zg�fj�����$�\�U��w��tT��.�2v�\7$x��(���}wm�}\���v�Q�/I�!��1��L���?�f�iT�O�7!Oi^��C46�iS�o=Yo�T���l,n����ST��C�[	}�ٷ_w�c�c@�4��N>���m��O0�OaD���L@Y����d���n�^��wb#*䁿�'ʵ0.lE�u|��f��p�ʩHy��Q�7UӃY�Z�%UR�a)�*�wj�Z��w�rR�9��3:q��g�,cq��0�eQk��f�{Gs7�E
�־*�~c��Ϡ�d��^L��L�S���q�7���N�Db�l.�U�1��ؕ�
���������`E���e�0\�*�|Ki!���(�ZX��hS�\��:9�A}�I&�����v�I��zQ\cg�ɀ��\���o��zr̈́�����y`�Qi�IOtƓ���JX�����;z2f�p�K����z��}٧�\q���7W�z[�'C
��@�B�w�0����o�<Ŧ�MB�0�q�
9����E�l�l,Y&�@#55KG�MЬi9��ɢ�4X����w��$��Z栊�P��֙0�!y�ݺ�}���r?pÓ��r�:Դ2H�<��7V8�h�ʳ�^�6޻�`GΖ��RD[��5V�����]_���I�������}'�jA���^P�xr����'��܍�W��'�r�3�:q�'���9]G�\}���F,���%��z*t�b�h3?�RbA=��}8�M��v*���S���$]�-!Z�V���s#�v;Xq�7��Q�d�VޓL��Yp�>Q�Q���"�e�! 6'�XA�o� /a<m�zl��wS�L�Z-xldݓ,�7����U���W���]Ϙ��&mh<פIvn �
^�$P����Y�z�V��Y��[X��j�n�&iMEm�1'㨺S8���Vc:P I����$8KD<�����ep`뭀EO��W�}������u��O5~�]N8
��|��U��$˵(AE�.�0IS�c�`��9�6.�̺>f�(J��dWۨxvR���"FmF܃b�p=7���|��u��P��7���0�5��P�R�!�M��'#���m��v*��t(�*k>��n���?ԋ���m�\��ݩp�~k���z�˔�
�^�)%�gCػ����Q�}k���3�z�<���ӾVΌ��X?ەQ�\G�Oۍ�(�a���f�a:4oa�]���g�Wna��T�p7�i��������[m���cjAð@��?E(tB���ģ���x��l��Ǩ��fQ;������1ގK����􃂤-�����\�G�
y�������տ}�W������Ȓ�¾�麒�¤�yT�Մ=�:Ml�����+�;	�v�t��&Kum��L@1�lAǧf6�j���IfB�:�f=��9h�v�0w��]7� R ��+Sf0%X)�jc������.PE\�E�
�X��	�0���M�ip��q�d����.8S
RQX.�<:Q���[���>9����_���޷��<�U�ʖ��ɞ��L������!Vi�z����x���@N��.F�!U�^�ZWR�7^�1�>!�{�BX��n�ڼJ��_|���>�L֧FB��GI:!�,W��y��(.�J�)YqA)�O��G���\�֪��9w�����˗�|�� �N�Y_��#[�$�L���i0�e'��UkC��ɭ'Y��;	�ɠ#�jj���~�a��澥�*�:���=/\��*�}��!ù{P�b���}��G*BZ�斳�j���-���'s��C��i���0��]����wk����Lܣ��A��������毪U&�I3=&��C_3֠o�B%�n�:Y��5��f'���b�F0�9&b��wO:��{Lo>:C�N�*��YL����o��Ȟ ���ز���E�0%��D���K-x�\:zfZ̈́���@�F>]C��1�޾{���;�A��V�>��ʕK�se&�,-��pn�,W���m�/�gZ���Æ��!�X��Ұ�bt+Ld��
b,�0~�����r����=�yD�y��_���_���3��1}�ܫ��ҭ�C�p!���"��H�����z� }3�q�<ulsu�B^�	�=T��MH����P�~��7�����8S�ȥ�.�1����������dP}x�gh{U��g+8�.�B3�����7���R����c*[ɪS��g?�����5�7���W�~E7R."hh6�pd��\*�K��3�Hn�<�	����)������lx�J�����-�P��hJ�]�Xt[��Yo�Z�ƹ�\�a:�?���s�7�h�ֹ��w�I�\�-~3����N��4҂�^�Մ��	��]�z��P9r�Rξ����Ƶ���_A�ƭ�舅To�>J�Q�Q�v#�?ki��֭5p�����Tp]�{����Ӻ�����p�@�Tn�|�`�Q�=�kEj[-E��m$��:������U��l�����s۽�fj�K�U�o�������2]�gKmV�|Q0�n��ya�J`��Ǹ�b0ny<��3�s��	�dc��(5�����-z2mܭd;��\���n��z���dW]�ܿw�}�o���<��ęW�Ի�^��R�����<_�ǫ�1�U"@K�r��d7ku�yHovAR�E^�Hh�B�G���������Nc�L+s��u��A��T���+��Z�I0��]�����.�=���[P=��<�rE��ޘ�
Ț[]r�n;/8�����0���/lu�����������fX��Fέ�T�I�����w<�#���h��|Gb3s�V�xs �@���]0]y��BM:�m$��.���eB���Wv���z34���W��U�����#\��2��F��<ޒ>}/��Y�fn�嫼�ܵē_��ͮ��RQ}V��;�A��v�C��r�������gU�	�D�6�4'>x�^xJ폒�C^}=ҕ�c��?���3vf�7�On�{�7~z������L�����]ԼD�l)t��w��tny�v=��-��_���o��᫓�A
t���{TeAD�~?׿���I�r<�!.A�H5�X�1Z�:�`�0+��D��?�^o�g>���ﳷ�ySݺ��#����?���<9{��8�%����V�:��)���ss��,�Gx��d�w���.!�����x5�;#���������xٍ�m�I���ձ*Lr������}Z�:�#�P5��rG�j�'YRX�_0c�m �_Y>�����E�"�U��ƹWI����ո�7�@y_����d�+	�Q���v/���1�L9��h�4_!�N��YZ(���|��(%��l}wq6�/7�0=��zcՏ��(�#fj�j��?�z�Y[�7~����{�z�zƚZ+���<q�J�_��NzA-H�V~���78���l{�Z<��r����fGl�'R��e\'�S(������P��rx_W�ň�n��&"�76��lC	��J�~����D��Z�,�����sm����Q0��Qw��D��3����Vs���m2f\\�PO�o��{����.�����v��8������8q��X)z��8��4߇۩�cW\F���8o��&��^)#�O����1+�Ђ$�//Խ�������O6��u߄=�Z��B�L�'nݳ��y!��;w����l�󮑰��}���/�VVR?Ͱ�&�n�eT�+��DŁ�\m�M0^C<�肉%pL����s���;�N��OEE�{n˜z����}�@\q�A�W�	'�`�3r���gP��ib���(�
���C��d�R�|����G��Ӽ���I�^���s�Vvr,zl�4Dg�sFe+��V�M�����Z��&fȖ
�_n�wƢ*P�#��b�����v�Ǡ��,�^:V᝙��\8�oϫԺ�~�؇�����������������yWI~��O��>��ZoZ��٭8sМJ	��$�� �i�½����Y��n�gz��>v#&T:�j�5�8���q���q8E����sn#��A��j��\�/� ǵ�Q���bi��e������y�T�mWN�o� �Q��=^��r�Q���c����A>�>Fr�Ø�Ƨ��'�Q��ܰI&�u[�tPWQ?Y^A�"W]��(�=�:9t?�pU�j%�?=v|�c�y�W���ˎ��_��޽��g<}��ҽ+v��g�|ڔL�)Օf�`yJ�^m��N��k���1CA+���q���$><�@��s[�MR--.�Gn�d�
�ÂEV" >�14�i��?�n��E��D�mv.���� ׅ<A>b8�L�����<U��	�B$�r�#jTX[fZ�w,��zPP96���֎�8�ĵq�Z٠ؾw�b��.^ �&��QfN��Q_��	8��dۂ���G���6/�ҽ�s߹�-Xy�����x�J�ǐ����4o0ǭ�V��K9{];�ˣj)��A�P�(GA��ˡeXJ�q}07%T}�$<��6��7ެ~������J��vKw2�8lD*mQk���e�ѤC��9==7�ٕ��UWT^v%<� \�F�����c�����:���=ߥ��,ޝzm���Ǜ�$�a�G�^A�Z�k���߇d��k�T��!k�I���u�}�*լ�!Uh�\b� gѡ'k���k��.J���f�����?x�.��D���&Rf~��W,[I*�ϼo����>��Y7]yf:��"󣧳,q�Ж��d�S!�=�)��a30�������/{��JM�bϋ�'�X���me���*�{�/	Y^J�Cឣp��uXZ�4��z�h�pQ����n��ԪQ�{��ZiT�貄F��v��;ƥ�z���0ZZ��@���c����/�%��|C� Q��7�u��'�l��bH��^��%�|;XV'5�B7W����ѥ��	��V'ySXq�Ћ�&�rLj=��u�k�>ю=|�~��i���)�G-^/ެ�`
���g�';a�|�����ӛw�M=��L����I�Z��ŵ�� �H'� ���$ve���m7�� 1O�
D.��e�vg���� {��D~�B~5OT$����l��s�أr~~���r׊N;ћ�k*I�%28�^�p|9#a��|@í�f���&+B4�4,�F�/���q���T0��\�r0��{Dw ��L�/!���͟���Y���/��._�s�E���ܵe���6�V<��I�mI�٨:��4Je�Q�02YY��.H�6�LD�値:��ı�������e�c���)�����c��,�su�׋���+�}��L{Z4f��j0at�&�_�����)jY�m�՚	Դ�2U�t��C�]{]vVz�pl)��3c���k���]g��~�0����hq����iP&%U�6�Ʊ��$�qB/�Q�L1(��i��A��̥��Sށ�}]-���O$�fe�Gj�'��8Rq�{=�(\�U�Pc���,����Z������޿�r�/�:�\�c�Qez��*�;�{��a����O>�A_�����^�x`�=���K47}��V�t"d�R�BuK2G�K��"�ß�Z�В;Mb%�̵� �V*|!�@��L�_H��0��E\r�����\�R�-�%9�wk-�^V8�n���D�����o��8
�4V�D�>D#l|W�� }*o��NP4ky�eX0��'�jM^�5&�s_zr��S�DC3�t|'@�딉.b\ E��pL���i
<��,%S'�u�{Da���ic�tR>�N1�m�=��=59�^��Տ�<��N�lH�5��+aqk�@p�9VX�M1ʔ*��E���Ot�s�\�Q���a�9�TE!���2���|W���k�����W��aq�I� ?nT�F��9ԡ��'�*����pݙ��7��Eo������I�ꑤ�J$ԉ�E�g��7�܎��i%�G:�D��k���G'�����O#lP0����Q_��?*)�W�h��B@k�N93�[���{��C>�A��+�(�8B��j&�V!	��Z�6i2}�����Jl�׏�31tf�U�p��U��(��_�N|��R�&X���wQ}��n)}��f1xu�!�J 
kɌԕVA_����5�C����@l�l�2s	�+��'77�(f��Ѓ��	y2�'lY`�j_
��6?~#�t L�E��f���S���3�?��.z�]���~q�`R�`��(ݙ�{�*��(.��>̔�S�7
sSCJ�?d�	kP�o	8��\;��6Nr�$N{E�Pf�0R��P�pJi�1�if4}�4ﰄ�jV��H�c���FJK�/�C�������V
�2J8{U�2C)�Yh��p��� Đ��Fc��Fʍ6>��FJ�Mr(h���Y϶d&��v)+5�^�YGXh;K��OA�^L��R[`�"����P��&�
)��5�g7ܾoat��������Z�?��l�@I'炳S�A*�)�ʙۘx�[;Łt�I-�֏�A;=�������0S6S��v;AYTq��t}d�f��X��̊Nk]p-	GG�Ղ�|�6��v3����s���L�"�a�`2���E���5��ױ�����fpr�,�k�~�`4s@v�B�^�gDqS�&�`�O�7��g}g ��%��f|�]�D�2�m\8*���9Z3���L	ʰ�&C8
5����V� ����:/�6!_�ܕ���)V��&����ќ�V�0��`�D�2�~���eV�
��r-59=G�۸ܺ`�4K�c��bE�\�F��"������N���޹���Ǉ����cF�f޶�(�e��fi�3!#���bl(F�G.x��J<�x������5�t#��q_�Ǐ��$h��`���6�h�k�F�C��X$��y�r�&s��PX���T	�itۤ8xR+�a̘�C'���Ǹ;w���B:],����X�	�c�+���%�������{	����f��J���B�dFh&���q3�# 6Bɋ�β�ԏ�<���:�3Hq�N�_8���CuxnW,LC14��m�D����db�	�ݫ@N{}n�4����?Y?Kx�.���Q���:��jT�U�.��+tP��,˳uǄ�J�L ��/ZE���^Xh4��U.��!��wH�%�8_R����itR�j�Ib�#�l��V����c�������4r��ٹ��c6r+w-灱Y����:���5�N�
5#P��`qq��~�b���cu2�������ZB�Ht�-�����\$�D�����)j���q�����C�c�pQ�B�]M@�V#x��1�NK���P)2
3}rw͉8r���+i��j�F���S��e6��5����(UhS%[h^����5^�D�P�eztm3�g_P��%n�eM�ߋH�w� |�{4���#c�2^9c�%���#��WC�$0Ug̯�p���a�ōXP	��(�*0k��2�l7�
g���,Bg�'�P�Ex�^�/rJ���"{���E��Eu�ЌC�܂�l���m�������[��_�a�0��8�K���`�:ɚ��V��̐F��&B.�����8E�(_��uprZ�(l�
(��y���2��f�؈��u�z �\O����*~f\4#O�,/���j��2) �r�Ox����$1^��މaD���^�d��1�Òxa�aq�<�,64Р�ED�_�Y-'�X� ����'�۰0��Rք6� ����i��jHQ@����]TX+[��(��A��Jh�(��	bή݈cn�U
Ņg�!²��4��1.�V;U�k�˼)�5���������x���S���q��X�~=ԉ.e�۔}�d|ƎpKɊQ}b<��`&��YI$���WɌ��5��kT٠ [�x(r
�o�%�3d�Iș�k=b,�z��d��q��ߥ�F���:9�f�ta����������o�HB[X-_i���hpS��,�P��}Dh�p�ͧ�k�)�h�jO)���h�?73�^��G"�y��4�i���Z��0Ho�s��&�a^F7�͘R���
���R�1�J����]v���v�b�� �_��5k��C��9
�!�8z"�]ţ08}���2h�Qmd%��$]��Wh
K�3a8>h�I����)*H����f��c�0��;땩+��bGȥ���OO�򁍮��7� 6B G)�La� �L�^�-*��%��&T���Z`a�.(t�T2������ȁL�n��(v}&��MHr�{�F�7�F���G��ƃ_R6��G��y_5V�uB���u���/���c���Ɨ�!�Pf��UJts�0�<���;M�9C��M�����`'��0�;&y�BC3�`���`� ���B��|�}��`�'C�������ǭ*Ō,��
C]��+�����+ث���8�]��o'v!cze�}��Ӡ6�߸I��\��3��h����44_1P]qW*�NԴ;+61sS�j��C_\��Q����&�	��[,�0����qq2$%Ja�V1�VA�B2�B+���"W�)�f�)"QF��Hi���1�]����a�o��_%hJy�G�I�NЌ�����s�� ��]����#�Y��NqbbM)T��ꑇ����D0
a�^h#X���;YKd<�Γ���$S}�ص�O��V?R��Jڶdo��V߿7��u:{�ae{����܅	�
N����ٻ1��Np���q���SO
fh~���O�r�����Go����BE E	Uz���$�h�9��9��	���&d�Z1o����d�}��9��f��6���
�]tς��։(��`�Pu]hR2��HD�j(�b-�ur�Q­'�m�&I���i�0��������*���s2�x;"��^�;���K8$*���B���`�'����{�%�C�^������z���כ�SH��h!��1Lb�:d�j�����,K]w<ѽ)Q4k��fP�|�$��+��-�����q��8�^�mP�s�%m���]a��G��$�Кz��4&2@?��T��[�u�rYi�g�����`4h�8�סSr6(�XzJ����� ��L�X��	|Z]F71�Wc����\�2�S%q��(ܙ��s'}��~��prH�v����0V�wj4SX���m��npLI�۝cȋb.���iv�\�V�k�o��<���X���]�p���Z
�"�0��!��?�!�v���H�,� �`�w��R���@�OSa�b��B-ܼR�����X���1�c�}�`�����Ƿ��VN�a��/a���M�2��{@%��|�+uu#IZQV<?ZM��X7;����˵ʐ�L��K�����Q ���/E7�a�*���l�*J[D���q�Q�����*��𫰖���~Ͱ�����aԷ6ר)���87�Q�QH����������m��oV�$f���N�"�j��N����*���<KPaW�$eBkd�;�+���>i3	�r)�(��i���p�BiѬ�T�S��HOf��c�o�5�J�V�ҫM��������_l6��ŌQ�C��
Z��ZXc��y�*7a^6��ݷlq ���$u�YαD�2B�K;���&��;���i	(&���^o6Dh�7�{�{.�_GC�h9����h<�ck[�Do�� !��D< � �n�ޑY2����r�m�L�T%q�U� lx�S[O�G�-?��+*�vA0S��[%e%H�U��3i�ނ[����JYk��G��V@�ՇN�5
�����ds��ۆB2�S&�;�7/�t��T
-d�ēyZreq�E0�OC�,�f�U�X#5&M����A� �ۈ���Y��s�[|��@���+szUH E�;`�l��ǟ�+� ����4���'X۽��Ud'W�G$���HZ*,�{�'Q����f������K�,M&R獿����O<�J⎨�j.N#���Pi�N�8�>�!f�!z���ͫ�vn%r�1I%�9"|빂{�Č�Ҁ�/j?���K���~�|��~���i�ję�����%�z���/����av���T��n�D�N�E1�Z䘼
����$���$�ঈQ/�]����<��z�r@Д�sJfey#�Ÿ��{�}����E���}$ux)��ӌ�n�3\P�L��UCu
���D�\9L{t3�d��!g�5m5xya��Tk��$�	i̼bo`f$QY��l����<jf��Ɂ�,���08 �P��}A>>�ʔ�����q�)���oL�����w�x����+�t�EW��wb�1\�����|s�8�1tSIG�hEUŎHT�ˌ�/�y%�,�s0���Y�l���"!^�4�2� V��+�Ŋ6�׆��,5��?n�������lt��!�b�8̑��D.�	�s�yZ�D���҆�j'�9ց�%�iSŝ��`%�p��4mW����чf���^mvYF�l慬�9�K�j5���O��!z�Ņ��5[��j���K��!�T/�vT+��"Zt�)H�uCb�)�+�<kr"vm��
�2c$�zUH�F3VK�,;~�}wE�'�+��WD���P/d*ٚN���q�|TI�"��h��	�|eF�$-�Ȝ��X�~ٓ�xmي�j�I\0|����b3�A���C!���
��C9�	Gq�c�[�{�z��N�Ͳ��?�Q���#�Ja�v����2���.PM�w���D�P�V<��<��
*c�hM����Ke���Ŀ�6ә����X��x�_�_OL(0�Wq���JZ~/z���Q�L*)IF��!��p>S,^K���\�͏/˒N&�S~���Ź�J�R!j��E����Ó>o9[���՗5���b��6q��C&g�:�`�q0OozI9�0���m<Y>_�M�������?��z����$��L���*�A�B�W'Z�-��m����j��s
y'��ɥ�Ƿ��_��|�ܱ%8��U�K3�!���:dI�Qa4X�͢\k��'�%sl\-:��ȔѢ��"/=�Dɞ�o�=��%��\��Zl�����a�j�,��ð��F���P��	����Vk�_���l�O~z�̓:�'�l�$�D6��ڻ���X��L<S������\/DՋ�P��\WfRb�R�UϜ��串0AZ(6��R�Bq|�I[j�4�������(}�7���yQޛ�"�5��#��a�f��T��}�����关�V�2������K����^x�{����C�E,XVA�>9��IR�*�ʬE��e"��� ���&�`������PJ�1_83�����U�b�����d�}ֻN�y�<�8^DȬW?�����s55��+�Ç��r��ݓiOA1���L��\��,=+K�{O���α�%���3��F�jtV�g�O��rO,ĥ���J�QMm�~�D�u�dx�,�uZ�1[���[�=/zpS}/YcJ����Y��׾������vw��.����z��1�h��q��4~䛶�����4kć��;���ŕ�/9�����/�t���+&XB8'������.���g9a�Y��L5�i ��	�W��q�"
�C�F��`h��	��R�s��[�;'�jY,%�l!��l�c�بU��EG�!_�V޲����>�����a|�:�f��'v�'�m]�?����t��+op8LyH-`&���s��dڣA���s�����Z1��7�����-�h��$����ݬ��a�c�k�����������n&�<9�F�>�t����}o�//-/>Gk�U��Z�H���Y>�S���\f���~�ox�Y啰�!d���Z������u8�<��V�b���-Z5���|�W"J̬:��J9���%�� 8,[c����8��s���L:It�y�i�>x���h��5XZEG���"���(zU3��<����o�s[���غͫL�\���v���*r���8hH��3p�	묓χ�%�6m�+�����R�������M�m;�:ѯj�{8�cn�KF�` A@@�&@@��T��F���sx�_ԟ-<�)<@p@�A�	*2xA0�l�@�D�{s���XU����Z{�}���E���u��k��U����K3�}w���1 V��zq���w�����`�۬߼��Yn��r��Ӳ����l�0�v�mu`�N����Z�"T����G����>y��;][|d!�3�^V��~J��5g�6W�J+�+�Sx�v��&��]t�����l��b�[G��9�.��ۘv�e\߿���1^|FL��|m���6n4Ҋ�PJ�Y��B�&�9T�"Z���'E�����{���t��v����l���T��g?z���#�Y�Yx~�ѻ��Z�߬��'��{��^>��/��&��Y���La[�h��	]�B3ơ��_��
��Ic��fb�L#WK�=B�� #\e]"'�+QQښ��e�~%�.l���i���/];{���N�*�j�wI�!��x��_�Ǐ=��%W��?�v_�)��5��Lv�B>�L5D�]Ͱ30�%�/���(LQ���.��[�i�(����g[]_��1W`Џ��"kwW+�i'k'�g�r�����|����fQ�J*ƙ YL9�D�<
n+͞u�������3S���3��O�~.��[8��
�$��b)R[�;��eI�dB�u^�@!��	�|B��r���O{T�U�8�x����i.�\ڎ�b�9'cF�tqɧFD4�hh��ȓ%��di���Ҕ�u���0����_�����?�����r��<T��}��TU�1�Bt۾1���H����2�#e�sFC�4�D�:���G����"\����w}6��͓��TY��=�q��sζ(�+�7�2*!V�pAF�i3y��"!�ܹ�Ӫ=��˲�^\L�]g�P	����kl��ʄO��ޖv�Z��t�A�@�ư�?���
{�T�r�_^z�w�K�+g���/_x��υ^k��T�T�b�'���kC���ڧ�?9�+J�)��sl�ĭVR�	�����!�%a�JS<��"e�q��x���l�*�C� �Nr3i�<e��b(>+�R�y
��j�&���as���҄">ux^��p����+z�j���rZ�i�m%��읹�U���T�{��%RSع�^*�+�ً��G�e�y��������w���;{�����ǽz�	�N
m&s�h��%�ޔ�m9dfs]�h;������㍝Ʃ�3<#�Q��h
�[�Yr���y��]�G ���G)L�� ����3���8�K�ΥT�&���E
5��\!��b��2t�S�6��q\陸�|Gw��/�O�s�w���㿴�w
^�H�M-��]��Zx�V3&�+��'��CO���'.}�͟��W������P�P��:�)�1��J�jڴ'U����ʗ��"���I��\�7+�^�� hc)q��|�2�����ڪ�=4�O�U��!�G~�L��1F�Ŧ�2�]+ȣ�tȦzs�ME��Eh;��J�����T�ݻ޹~1J���*��]1[u��+�em4�W!��i�9�->۵����=pS�L�*ry<���|�UGO>��N��������<�Ԝ���SQ�5K��\�|��^7|/:f����5�\/�5��|��O6����`IO���{�[�m������kfd�i��q/y��������:�O��%�X2|a{���dw�$�Ė���5�X����Ie�d��3W�}2X=�����~7Da��,�5�6e��+l�����}�r{�=2�����=���]�=�^�����QD=Gky?�7;>=t��x��a�1�`��}ᓟv�������y�+��ҏ@֟���d���W�f-�DG�����Ϻ����k~�ƹC�~%\����yG?�ڮ�YAlS�`�'�2H/�"���P�l�T�L�ܶ����B�l"�СH�2`��*��/-�H�-i���T6����U�c\u� ��¤�1��5�#R�)i�t��iۄe[=W����bmL��:ʲ��R�����tN,N�a&�=���dey=�,����k���ޫ:K�µ��a�0b�7�cp��2��_z�G?q�$|�����z�K��#ߡ��g+׬�Y$��|7�o[��\��� ��}��^�p{�g�����~|��!�j�w)�v0�u����MV .=�RJ�#�Z/C��� �~왻o?��'����sw��E�
W�o����f]..,p��d��	R�5a,y(�F�1����m�xs��"��*B�<��K�+���J�O�[L�չF��O,�yqg�� 9�eOg/�Y~���wY�&�#-�w�m��7�P������C����z�A�>a�(��(��R�2����l�����蒸�z�K���L��%�O[���H�c�z�Ep	C�G�Aj��v'�P��R���i�25J�_��f*�8=�/s՘�N(�$�ѵ���h�	��$1����k5��7���D�`-ɑl����@GR�m�����W[�A_��p�)�S��qQ{J��7���0���y�ŧ��U���[揟��dy����#��-w��,��.�,B�Q�K��rp���&�W�t���2������7q����>�˳�w�*EI��!gR��~I�O�y9���Ga	�y�1f 2Ҍ�(T2#ܻ��}Of���+�ж=0.g�ձ�~Y?:�m->����{�g�/�+�(�\�M6��߬�����+��G�!��7�Ο���;��ZM%I���͛�%"J�az��d��
ԋF3�L��,|� ˆ��\O.�W%g�/ί\���4)PT(���L��=f5��������S[\�'E.���A �ߢ���d�YՎ[�h���&�P���4��)<���ʕ���j���2�,���C8�3,][ӖY'�i$ʌ2� YE;��S���W>R{��	�cPx���y�bM�R�����\��f��%(����cD���㨨ߧ�ST�(�I[���5C�BB�P5	p�:n��k�)��γ���yډ�	Z�{���y�Z;�W?-�.ga��X�d2��VB�W,���Y:H����藱/�2���凬�ke��;uP�Q@���1���c�l �9�5�����}$	l%�>R��dQ0㳐'|VU�P�M�v�&�<j5����£�4ff���@|l�F�+�D��2��[�xS�sf&��D��Grh��"�D���^&���9��ɺ�Aq��dZ�Q�miӈ���/x�����pT�j�f�YSv~����S��1�Iru~�b~GSI�5'��4h�%�!�>���#���l=�g��>cmq�ɍ�����P��#S&�2���(6^�$1��lx�6y����w�E��xO�R����� ��Ā~T�&|��$ΜH)W��r��	��H�pV��)�4fmK�i;bzb�''�=q���s�>ng+�/L8� ��NTq�������u��
��Ҷ'/��uO��(��iOH��*o���[�"֊��Mw��n��	O�felpUhQ�\t�������@(qH	��CG0�OQI�6ٙ3��)$��F�j2\=c��o���I�4�l`2���-��6��421HB���$2���ڲ�_o���Һ�����+b�M���j0�b�*C�y�m����\��v[g�<�	�tG)��HuʃFM(��T��ybF�a^f!RTgmt�}#�U����ɛ�Bp�2������s3����9���k��Hr��(펆��a����٠7��l#
����%��s1S�rA��#����fO�j��wS���Κj[ۮ}_m�Zv�*��O�2���b��q�DsbG7��2���9���ϵ MⲘƠ8�]:~�V����W�pvwd��+����>゗�FȑD�(�to��sQ�MQlJS	A��,���c��4�2	�:��� I�b���Y��7f��W��h��թm�������/�ķk�c� Y�ة�ù$�KiF�����~hʡp�<��<�A�뫀���!i���/!N"�d��4�?/�E�����6� ���<��i8�lOm�G�uԘs 6(h�J�#�U�`����'ay/Z�Q��j����\��ܼi����.�7���Yl�����rS-���DkPL���zYn}`�4T�p��b���
.X}L&����򈘚"2�L��#�N��D���kt�P3 ����P. Z���h"�qR�	���|����+U�*(��/=Mӊ�������κU�A�OD��.@��^>��F�&�r�.h��aj��-.�&��Y����9�����=.ϥ8#��_h�zI��N���1f:����4z&i��V��y�ʠ�����b��=��h�%,���.�����C��l�.�՗;h��h�9�R����y�
ށ�� �*Lhon��E�䨱�o��ep_S@�Ti�ݰO��C�n���w�
�R��&?e����23/z�"�-9�|��̅b�w:��z[	ޗpn��2'IR�޸�������x�v���L5,U���Ht� 6�I�r��g����ᐋ��N�,�\3$���E�P}Ʉ�S�X^�|�N^�1lb(�@�\��4DR�W��E��Ѝ��(%�eI�_^�����&6��3���'o�Sb�ށ�%�;-]3S1�����5k熰��f�M����yp�)�8�����h1?�k���`L�ʖ��?̝a�M;�T��!1xf#'�zN�몯fp�&��}_F�g��������aPP�!T���H�[���_� YX��+k�t�ч����&�[�'蔁"�`��[Ǟm4zH�>f�f[-`��[����<e0F�h"G�+aLy/Z��@�ұ3y�X!$H�s�J��%��k㌣���S��2*��9��ȉ��<BX}	��5�كr�2�J_�9�#��=J�0,�W[�A�A�X��]�{Ax�L�+�o]���'oc��4��f���hv��@	����[��z��B�F��.�3�p��]+���%�Q2G�;F:�nԜȳ}���3�M4�\�!*l_CEW\�h�1?I�\���w�3��i�d�F㎶x��[_��Y,"�Kx^q�$��W�kR�*��m��=���~�0�ȳV����gUm�D���912����T��l��TQ�����.5z�|3�����J�r"?ԍы�FU|]�R�*��Z(�y�G׬�?���.�m������3J`��w��������|���}����6�/��h�� 3�{EhS�V[�(W9�y0����d��H�ҙvlw�l-A�5�k���3��JՋ�9�/��ţ��%��<��`Z�Y�j�͏��B)��;.��*���5/�6�l;ά-��F(-������7�2�䐔9��-,�{\΍n�����ͼPŹ�M���;>�۶-�I7��GO�եT�?%�*Ƞd�����ʢ�C��c�<6�G�����E�5�ذf�Vz�m($}�v`p���ӇV[a,�a��Ԉ%�J��D�GGU� F�9�Z�u���FUį~<j�z����p��u���(�`^�J�� U>�<<�bE96�v̭
s|u�K�S�˭
��F��K���o�~�ߏ6U��T��Ԇ�(+Ε��!ݫ�����PU�!�Qh׶q;������Nn^�c�gΔPV�)���EI�[lk������� `������|����k�V��fD���0H�:y��3���&M�*"tٙ��g����|��e��ѣ���>�c�����g\+B�
SW�(Y�Ύ!`�UqN��z������61a쪝C�oA�Md���8;G�
�H6�WH�U&8�h]��т�\�����7�;�{-]ZX�Y%2k�fo�$s��a~G?H��:@�/25K�_iE�@��FlZ*�[���_AAm�e5KU�n�b�#���wQ��r���?f�Ä�J��y��h���丙z�^>8������g��V��7n�}�2�A_��ɣ�bm<jF[%)���@A�?����<dj�ɩ�fz9��S��X^!���g0��];hI~��8�G�)�mR�U�@�:��=�~z�嵴9S�/�Z��y��b�`B�LEui<Օ��[΄ۮQ��PD�����*�6h�]���I�א�7t_d�K�v0	Vz�Ȇ�b���o�OMnE�}�رG[�S�r�͞������xdW����?���Q�3R���<f-�u�����z#[9��&�%��=����JT�Di["_T�8�g���T!�&���oA%Կ��IcS*V:����B2͙]A�����X�[=�@l����Qqc\'��k��m��xj�Jٸ�ܼ��  ]T�b��lQ:��5-�Hie
�c)�7�|e�y*�@A�G�F��Lb_ w"i�Uf�.!�Q�K����F�����7'қ����񗕋�[�F��Ӟ�nl&.�`H|Pj��$���&!�� #T��[��]��f=U�Yw�}"q�`/�4V�I
�W�V0�Ơt�����#��u;:��'�4�ʀ'1���4�c��7�B8<wP�j(�-`<���\λܶ�&�pe��y��I1�Xu�}�������7���ɺ�&���E3Q����چ� �OM�l��ڪ�t�ɘ��"������W����GF�pP[s!��L����Q�;���,�#<;JXB��G�̲�٣��S;�,;jB�ņ7W�^m5�8X�si˘�����.^�'�S��O���y�%�J��h��d;V�jb��W��swIW��aњ������L�=�+J�c&��������x�c��h)e�ZЏ�]i�4�Z���(F~�@%��}�{����:�y�"��V�׮HZKW�Is*�r�����rU(}��-�B�g�<��O.������G@s2W`-il�f�����LR�UM�0�T�� �G�� �Z�(-[�p:5�XGl�R(��Y��8���W8��+�T������#�4ڌ�߉�T:&�|+LgB��~W�,ȋC�S/B����R�Y�]8Z�}mʵo�s��]����G
e�K9KAP2�ejjX��X��B�,kþ�*�Z�1�:���_�Mӑ�^=I���xln=��%O�q����,�!Ѳ��lf��*Ϩy�%�����%�l����@1_�n�E8t���~z�k<t���i�r����n��,5�61�&s;Ͱ�������_C,����]k��m1͵�U]�S����෤{�����e�	\�W�\�����e�-�%e@/��'׸w�����̜8�7���מa���ǚ
��7>t��{���y��0�v��/��?s5�A�K.W�~��W��M7�V�+�e˛K|;]�������Խ�a��|���S��y��o��3���C��:Rn?֜��d�ܫ\���(vD�vc�>���Q=�T-9�+7S4ѕ�I�o�~m���8�ė�=�x,�rd�>2��{�[���X7��Tlj��D9��;�V���� �)W����Dd#ʈ�sY!$J�c�]�Kӣ}\�������p�5I�"+)���`E���)L�x�s:�V��q���9ϻ�X]đ�U�)��:LE�/haN�f�n��WU,>�u;����i����|��wP�Ztj�Ne��/��Z��8evB�q�ȗ���e:�z��׶^񊸸�9T�n}ޥ�^�*��[�J���L�!��zl#���#AН�c!Iv�RQ�,��~����	UG�*C����Ycl5�M�l�3N��4��}���k�(��F�$Wϓ�?yz�J�O���R-�4�%�ӕ=)m�ۀU�"!���'��4[Y��gf]�{�ķk�O£ݙ�b�6�G�z9�lAPTG�5f�,]�
	�L]���*[U�{7�H5�t:
��]���=���U�jӵ"KKD�m(���w���. �y,�5.zEp%�Yv��ǎ��r�:�ˢ4^]h�����_6�ǋ���~䎟�����9P]��4̿,
��^�4|��q��?u�_��&�/@��Ci��4p{~�O�b"D��Ե�[̓�H�G���O����OeVa�U0���Y��"(����)�A����`��H�S�����r+�qq��R��c}���ܨ��Ư8Չ�i+��*�F�F9�|.k��Y���E5�_ܘ��cj��!K]5	�ad�5S*�"- (']hUH�B�U��8��=�Q"]ݳ���T?,5�q����7ߧbù�1��/<3fV��+[LM�{�f��}뽕:�/�J8�����em�ؠ����
~P�G�$���f<Mcy�e�}���������˾�^$���Qz!	���]--�5	�x^9%�{��������)l�=dH\�2a�="���9r��"�� a/�q���������3"If����ĵ&�Cr�*Jۖ�@m�v>���;�/M]z�c&�\���:����	�>�3�\����+PL�'����ܛ�2�b엛��Pi�-���	�.!B2]���)z�[�x���P�c�ۇ��6���|�����K��JԄ��c�>3;�����f�t��bb��{�I��Y������{u�����lZ�{�ds�z���<�I�V�d!(�#�"u�3�K�p���5������Y�m1���guc�W�)�L}�!W�-4�*�oޕ}�%����l�Ѹ��׻u"l�>
DY�K_�lf\�edo(��2t��bg.��o��woy\�9t�w~uN�/�vJ��9AY#�O�¨�*6).�D�g�Rq���������#���։Fxr{:��>?y���R�C���R��ͶWl�5�����(�Ww������!�A��4p��;lB��=P�����1,�~G��Ԑ4����eƑ��u�.o����t~�--դ�1� ټV�uF�"��3{K��������G��W�t��R�Mޑ���������GKn~?��UI���[���'���o���Ca7��{�l	�1�d	C1�dN��L���C�<���˟���E�	�7SO�5��"�����&�=���%��:�m9�Whĸ4�i�gB��T+_�V���� V�Sп^RTӘC �����ӓ�ə��vӉ�ٛ��W}��� � ^��yZ{�ZO_0���f𹫛S����KK��q��i_��!�Ұ3��t!>S!���� Z��yh�]j�a�H7�XE�t�u�v���V�p\�����g�ob��������z�^Ŵ�5G��a��&���;�S���	���\�E��.k�ğA�+D!UA;������M�L,�G�W�M��7�/�07�����0�����y�M���W��T*�a����Su�U����=-�|��2r��BQY�i���vŕ��7�й.y�68��:�qN5�M[�ʱ��˚�,�����a�n��Q$Z ��5S�m�A��HX6L������H���i9Y�n���G�VJƖ.X�����K�����d�Vd���/� ���V^�&��Y�>�u�>�N͝�iO?e��m�Y��X@�o@H�9����"����u�}9��P����ۢپ�!JD�v����{@uz�UB#��Sa���į�����$P�CKeL������_�Y~�#7��O�}拟ug���H�7�_�r�y$�������Fm�Z�:�Kk���^Z�����ߓT��6���MI�62Sli|��l�B���S�҉8z���vݥ6ԎN�j�������Q��ӳ�}�Oq<)ѾU��)���ϱº��:����Y���Ņ@.,�C�+{HڻY	���H��+��겑�!���l�W�����`Þ���ٜ^�08����b��eެ��_6���'�������ݯ��?~i�ߛ�M�_�/�k<x��#an�lS�RfT���'k����g{�]�?9m�Oʥ�\ ����9�!!�MΩm��f���$��k�u���8�=��f=��c�hӳ��\�J����E�;��gAD�+�XmnS4B�k6O�3�h4.�2����D ���hP�8�;��k}2uY(I�JE [�h��2��Vq����{q]w7�@��I�5�xMv`׶��MtE,
x� �>o2p����;)x\c2�^5s���x�{-�v�r�����N}z� Q�Y��g�7ü�)`O�e�^?a�RWw���:ɵiL�Х؄#�D�2�������W	�VIc���R��0�}{+-h5W�ff�9c�?r(��c�W%��F9�����\�߯�&��3=e�O�H9)�����k
#*QVR3D\���3��Q�:&6�v�o�<�����_�`��P]�Cx�h-/�4}�z��o�i��t��r�l���_��������-�������VM�[ 	�cu�A���W�ʺ��_sY�]éBb�C�lڥ5��H�Z�S����R���q�+T�3�j$�,M�r �+��Ѓ��;�Fݏ�A�.#,�,�a��e�۶��nԆ0.��C�h��KK������q:�ْ�8W!����(�~d�R�!��q�.�6�L�9AU�2L�����u�]eB�[�
m4k3�v?�f��MW!J��y�s�P�s2[��~�"%wz��HP��H]v�`V-��̞v�jQ��{G���v�k�S��kiv�Jzs�92\w�Ⱦ"߀�y�
�2mE������[�����r��W�T�pVB�Q���)D��L��*̝8��'��ϝ��/,=zV��6&��,Dm*���pu��5��L�M��y�����3��)�%Scr��q��!b����XCi��tǌ:��Z�U(��Z�����2v�y2F�G���I�3��=fG"�"��A�W�oW��6o��� l��ύz����}��Z<���Y�8pG��΍���ցyzq��j�����%I�z��zP�����n٪]���l�lY�>*^��ڐ��2�ָ��XU^g����}��Q;c��1����	�ŏxbdn�"I7�k[�!��[�7m�a'3��,�p�5� �4�EFC!}�&�$Λ@���&,;�.�E�U9��:�Ɇ���%��\QE*eC-��ȫrl�� ӟSZ=u��]-]�,s�:���F���N*�Y�"&�e�L|0 �>U&<'@u�,���u�z}��A� ��,�H�2�\��F�G��;��<�֬�r�!�T($;#�����&.6�؟���:xMi�4@��7�8���8����O�3\܉I/f�t����>5���|.։9sѕ�d�|�܄/�A��g�����q<I4m24R��)�%�ϲ���|,�h��AE���wN_��kE	���(d� �+�w*�ȡ�̒����WhW���iJmgB̡9��w�k�´D*�Ą"��ky���"^ދ�ףϒ��^�����ۆ�P�U���>���Ԣ9-8����vi������-��KbZE�ϗ��bqVV��m�e&μ`�1��M��:d�n���Nty{\ $�#���$f�2>�h�<|�b��,� a�ɷ���-7�8���$N?	��S�`�xXRc{��&�C�і���h,����4���}}�A&&�&l8	��5�(�~�ﶕʸ����A��y��P��Q\��D;��83�#�B��h��=���ݶ����0]����y?������Cw�Y�:�#���S���������*��
���̦~�����{Җ%[���j�*S�@�"��Bb��L�5�O)~W�D�N�5�o�{5s�yH���A���p��r��w��C{��R��6�B���t��V�i�T��A�^]m%�������� M4j�}�v��QM�训1r��rm��N�<w6�BZ+T�a�i0 M�I�*%		Y���OdP.��v�S�є��f�"o�����@yN����� a8e�f��L�����ra�,�w��x^�I��U��\��Q|�Y��{L�,�h>�)�����<��ި�� 1LK�>��	�9x�� �°q�**�!������td�!dUi=ϝߔ�I�y�T3Rldio0����//�Ѯ�엁2�W��lC�YFА�F�������玎�OҼ���EF��.a��E�(��B���)�MON�_���a_��_g"I�6ii�;y�-����Qr��fP����[��!�msZ��窱��F	TI��^z�B?��B+5�,�9�P�̡&�8�P�"i�d2P�h�����w  ��IDATUL=��ޑ�T�sJ���t{W�"E�W�yH�*^���u�֯ު�d#�6��e·�j#l}K��Ѧ+�n�-�r
�zr��c_ҚA�`�L��6H$3s`��
����M�.i�I�X�c[��_vٴ3���%U�[[LZ�����Yz�풖ҝxYV���~�k��Q�๞%��$Z&5Y����9;�R��v;(�cQ9[���`�P����NL@��J���Ü��]#��jӌV�rCmD	��B)�XJ�K��9#�E��6;�.�v+H��F�]X�I�/L0���\�g�
_��-�8L��V�e�-@��|q�A�#���w��J���������
�'�c/���g�M���
T��A��GdQ��e��)ej�%��j��
��������:���!�z��z�Y�^��o�:�M�ˆ̎�_�����f,������j�����We��K}���iԲt��������q�`'�K��؁k��J��m�ж�D��e�}�&-�PAe�T<J���u�exJ��䥱S�l�D��mD�u6$���"�_���tG'�SeP�e�Y~�f~|'��!mMȕ����̄��6�P.�@4B�<$�����Z�lg�(�4���ɚmC*�"�����G��v�y���ǫ��~g���;6��9�mȠ�8��/3��<��,�H�j�8�L�?���%�خM��L�{��!w��@�ȞIQC�Q�\q.�S%͋�GO��(V�.�W׾j����H���ER�g:�	*�Kµ5X? ?Zٷ���kC�T���u}fgg�?=	��^�B�8D�ya{� �i�4�U���Bم
=,�Q��V�E�8�s�
��_#�&�e��`��o;]bD`�r���Z��J�j�J5M��Ut�a:J�M���]gj��l�Yb�\I$&���W<]��A��������@�e%��xh�r"ӡ���j�_߽~��|˒?�V�:T��͵3�t���g�L�tkyi���#��K���-3�8�mp]��x�VKB��'l4YQ��)\2�Ȗ�j�l�
!Jv�30�hZ��p
Һ)�Mƕ,�r�V���J��عd|�O��έ�� l�(�s��{����w��	N���' ������칅r�!�*9phq�J	�3����z�k�����`�""|u#Ƙ�5�W �Ho�����!�a�+�m���1�৉��q��H��j�@�q���8݀:0���LK�N��G�'�����H�'������M��E���1���X��	[�zz[��|G���<�^��7o���{/_g7-���P�F\��k���f�{���D��t�)9Y"��%|���I�{�R��%������
!.�auoJom�Wj�6:���M�m�R�]&�����7�P��s�5&�������g�+��{I��\�ձ!�t�)h^JG�RK��(ځ��-����v�xxUz L�6�v��r�"�JU�@��e�������l`�F�"Ş(��U�p(�q�-
�l�)����5��Ŏ$�_�*!Vi��&��w�8W�q|�#S�F�4�?eӚ8�A_͘���`��(��J4c�y�,Ȳ\�c�;o�-n�W�d#T\Vn�I�h���
E�۶Y��Ʀ@z�r��7���ըc`��*�ix]�����w�~���~��E��U� �Ef��ۅ��x��gë�D�s�s̈́���p n��w���CoۆT�v%(��f�BGјP?(+�V���u���w�̔�v{��4���HL���d	�����@�� wc$5\��#	�47�8�s=��5��:
x7DڅlSE>k����?30���kR�l*]��z�]��q�
��'oh�׃7�����"��:�]P���H�]>�NVв;g���4e�&��^`,�1.���^�&��>k��4e4M�|��*����h�fij�+l�$�E=��Y9l���M���#�S��Y:��.*�ИL�L'�4F�
�tjF���7~/�+N+Y���pK�%-<��F�L�<(��8�^]���3�T��/��5�e��eE��!߃�j\���1�T��!�ґ��E���]W9�d����N�M6l�R"�E�X��E�-��ʛ1��	��ŝ.xsu��l�&J�bF׿�~�O���-$�іe�L,�R��*����p'7 �!�5��%ԛ&�xuH���=�Cz���5vSb'����|&Q
u$�)��g�-C�Z��06�GA��������\��܇�PP���$lS&�O�L�_�2$�>Ԑ�X��Y0�\\%Iƚ��H~�2Ok1�l�HY%dz9�w�/�Wc5��幱�Im��c�j�d�����"P�ޭ�-��#3�*e0����p#ِ��$iy��s#U�m�#w�b��I�;]#�HGB���3� k(^F���,��LY�F���5�4R%�~��N/��x��/EѤ���f��-�՛�
�ߥF��<e:C4�#��u��	>���9�~Uv��5tî�Fm�7'@vB=/5�rvsJ%VVr�s��s�m��s �Z�G���r��5-Ê����2��H6&~�9��UFN6A-�h�:�|�4&®����Oy Q����d����$����)$���a��.m2���>.l��>32L����6xF`��O�~���Λ��F��w�����E�����o��ۆl7��/ �
z���%���uZ$�6�ْ�U��C�+Krp�ӐuִTk���l�t2�A��7^m��yFƳ�l�:bF�MW�!��P����9��wB�C-��S0;����"��
E&V�j�5,;N���q���9�M���麞kZZ��uz:c[���:�KS7֙����8 ?������U����1BM��1��� �8��5!����[y@(�'�g�Z=B��4�p��	6�x�4��"��R2��-N�Ҿ��n�c4һ�N@L�xN�#�t��&�gp������a1�\ڜ�ܲ%r�Ҳ�ܢ�\EM����L1Y��G��8�,�$�҃Y�0��]���˴��}����`��LNԂ��gX`���h��Q���1�KH�yJ��vʦJ��h�$���GInx�NN:�a�[6ZP�n�>����z���h3��R)�\V����>����t�}f�ݎ59��z��7;�[}.ZL'��pqԉܣx���wnՌ�f�`��N/P&XG�3D*���B�al�)�E�ó�).ֿ53�me�{o�ڀ߇��yG��۫+�u�I��W�����!��:��<Co8�+�%�����8�8��}#��ự$����+_u�|�����Σ=��5(��%,�X���Q~G����Y��L�OB�����5�i;̮5 �j\#��*%���|hLz�3G�g�C�I�'�� zDܡQ��a
W�������(���$��D��8��r���hjFrO��((Kd�ؔut~�׃Ϩ��0�&�	w��{��{��.������$�j��I��s�֬���S�\����hpֹp��C�%���v����G�t�.�v۽pe�u�X<�S����UC���F� >+���2�Mu�'��5�[�ΡN&��u�92e�(m��)�l�>ӬТ��Q4M^�g��Wl76����Q���^x<�HD�P��8�)�EY��Vݕ�ѧ^p�Gam��꫍��&��p
7zt�����u_=]�~����g�P Zp�>�YH[*�T_E�p>��V��S�q�H��7A��~�}��Nm{^���yߌ�_CJ��s���H`�qT�];�:��tN%B���zgQ��|�s�#���/�:��ؤ
r��Xf�'<LLE}��"4�Po]^ux��X*θL� �'�-Z��\5�D�� ̸ ,�h� ���Y~$��Cvc�WR!������O�i�e���R^��5�O\y��G�G��_�	Vs~Z�z=��	���^K�q�����'s���Yk=ޅ��_����rs��bu]�rx-�B�2o��h���J�b�H�~���<��u�����oV$��MҵX;�P}>�&����ΐ�+�{2�������c���z��� ����f����#ZڢdB�>AE#�>�UX�M[%~y�sK�xG�B2�I�2W�0Y�R�%w5l����)�����1yݍʺ����ث[^�o���)\.���������i�s��5Q�'<�3n잶�^"k1�d|�_�e�b"�����<U�au}������U+cn��Ø�&�=�B�\��zmh�I�C��*c��h�c���J�'�S����3�����a)<�
���/݅��mМ��4.)v���fA�ކ������}��c7����K�����Ws�ާ�8�#1��d�6A�i�?
ҩʒ@%���~���u�����_� �`^��ک��!<��~q���a��y��X�A棦��T�sp���bq��A!��?���=ԍ7���;~��ڡ�ω~xy�?�gk/�O�s�R�I����$�ƃ�1�m��p���+��b��~�?v���K�5���˪�k♉��-4&MѪV�Q[Dag��ny%'U��Jʵ��$���v����N/���������}qݔ��N��M�����Ճg3r�z�I��a(փr�jdb^T�غa��b���O�}���s��;�O֡��DO��-.U����t����:�sbJ9/���/j���XL��_ʬ���_����+�����/|��h+����,)݀��v�'���VT�8霍�e*�"l�i2F���Q%�w���u��N���,�/�*�i.�?�m��@�7��p�g��NO�9��wR�'H,���Y�k�*Nc���}$z��ޝ��n����w���x�%��5e�H�[x�t:|~~>y�M7i�/���W���W���f�KK���nHO�$�OkqQN4�*��,��T���h{��ލoq"Awʽ�����\K��G-���
����^�����r����@!S2��l�������M7-��k��]ׂ7��[o���Ň��Y^���f�q~凬��%�^@&0��6xf��Fn�k�vM�u�]�v	>B	>��RE�p�cFY�r8��1�eoL�}=��Ķ�zP	T/Yj�y��4G�XsCyT	FTu�R"$��	����p)H̓�^Ӂxa��j�-��~�N!q_���j�T�'�>�@�HU4	�UO=���n����D��7�,w.����M%83Q�
��XQC�a�7�hX.�A17��%�2S.�E�	L۴�զI�I|ɫ�;%Y۲�-�l���Cܩ�M��K�d��妜YI��"�kr�ST�ȠΡ?]c���%s����Ϋߥ�{��~P�������vx�%�f&��Q�H?��:��'����/�<������lO�PG�nBw��aχ���s;R���v��H��Ɇ����hӏ�O��8�j��,4"c)D�j�1ݾ�_������V�����c�;e�ٳ���x���]4����]�;=���~w�s4�������`}]��կ��յ�1W�����������
	���_�4�?���n������4�wsC��m*�!k��:�	LL6���:��o�������j�w�$N�#c�ujq�pz�#���O|�+_�������ǿ�g���O/��k���;����̖;�U��%�F��t�_����,�~l�ps>pC(cs�FH����ȫb�{?�R>S;
����!adȕ�s_�;�h ;��@P�Y��x�2X�x��J4=���k����tV�4��n隙��ɨ�ז��� o9�<^c�H �3]8�1�1xG`��YH�T��d�y��X>������YI��u��*�4� BCs�y�mɨFBHz/��Va��;��V�,���IJ]��1�E��g�v0�,d#������nz��]X��	༾
^���u����Ҙ�uυvl_�������so���7�~�/���_��1��(��e\1�6ſ�e�BS��v��@��S4r���1�~������?�یS�h��s�������CGv� %E�!��Cqu�F<#��T��y��c:}5�|Μ��c����/��2�#Ox�:���n�g?�q���ή~ε�����P7��?��o��t�yVWR�C[g!}K�˸���f9��Z�\ش����R�S�l�7	F27ˌ��J���LŸ�3Wd��+H�N�y<��Kv�9���F���ϯ���6��i����y����&����N�b����,~Ҭ?wzm��-���'?�>��[ٵ��Q��Z�K_������|����Å�C1N���ح�����BojU��a&�\ߎ4�-	<�C�	~�F�t{/a�D_��W�O�����FՈP�s-ߨm0.�k�(����q�ց,z5*2�\>q�&��g��\k��˵���^;6y(��,��q����n;ԑr�8*]yuV�L���<Ƿ�{�ء����G�i�4d��٧�#J
Rn���A��$����"
�9���-��dՄ=��N��Efw!sU�7�&'��[>:?w���3q����N_�Ǟ��ޭ1T�j�ob����P;�������6Y��~���B���:B��	5KE"n	
�5�L����A� zf`��,QB����x�.�7��?�q5�G�����$}f��׾�ŧ������P)e�oq�z��J۴��|��������##x����bg�x��Ǣ���
4�>�8������i8<]��w���_�&>�{�w�N�Y���j�-T�v;LZR�gݐ�}�x��,zb���~���a�,xb(���9���i�Yq76x�3��$�`\4��fڥ��9L�6�>$��V��./�L �5���$���9:�aޔ7�_]i�G��v8���O�+u��>��+������#g�)�p��DR�+f&o���Ӣ܊ ���}!m�}�੩��<��L5�H���X�Q��$d�Z�(ik��7X<��)H�X\����Ignx�G��[��߮5z�>�31y]�ܺ�~���.F�i��*	�)&A�H����K����7=��CO��}F{��Q��3<�f ����0���f���:1;�ؐ2^����I�����Ù	ET[�a����`�����m��
�w)gj���7��Ö]{R��<��(muP�vmW��C�֣ZYxɚ�����^y5ķ���g!R�)�2�m����Lj�l՝z|
3aA�=J,�B�I�f�R�b�벝 �9TL	�-�=�����Q�>�Pg;��*���䬁���٬��w�c����cI�T{m�W�J}RH}��
��H�D�ӧoz`e�A[�c��� �[g�-�� \��~3�pa�Q�BǳY"�.
�lԑ|8��T����h�F�XF3I����%�S�`>�U[p�M.�h����	z5m6'0e�4�"ͅ'NVΠTe��m�.�B.L��B��#�YV,碳kϻ��tj��~u���o�o�����C?++ϕQjT`g|rj��8�&����<U�;�f�6���M���Bx*����6��V�MA��S�2���UdC�Z��[R6}7���'�x�O��^��X}�ƿ����yϤ\�vg�?Vt���w�Z�v!Y�Y�Q�����������i���^ii1�hw��PM��%7�I���U�tɲ�:�R�όTRE\�JH�����"��)q*hsU�;[�:�h����J�m]�����[�`*��Np\Yyb��?�:^�����f��K�[�r�j����ję����"!>�J���Ժ�ۏ"qѱ-�*KY�i/���aU�:,�6v�D@�q�{�@�`�mE��jB��;r�¦@S���(�v;��Ԋ���n���%-�9a4L;<{�~�v��E�Y��H�擐���6a�>�fQv��o� �\;s�Z�0w$�Y�a�ZG������nf���Ku���U�q���D?���l@vMt2�fk�0I�
]�W�5��6�$J��C"bS�����!���ՍTsr~��ptRd�t��'�n�֮=��o�����K����{��O���d����=���$(�/��N��U�y���������%�ӷ���:%��jh	���r�⧙"Ӱ�&y��Mh�<f������q����_}׵�~��tx�Vk������H�����b���Ux_[=s�-O Q�;(i�g(��j���h啶q���B��R������:� ��a��w(k)s��It/p㩗6W� ��t=�tV��7q���+ֺ}or�g�!�Q"�h�l�tb8	u�N��������P\JT���5�5"�J܋�h&�(0�|O��!<a$y�&�`F!�'<�m'"ݧ$�P��tc��)WH���(��:�]p�_G5揫����ך	�|���e������s򑀣|�dw���7�w͏y��u��U�g}H��tQ�Ei\�!&�o���t��u���P�sf���N�����F6xة�W).�t�<K�Hg/ZF���ɪ/�A�e�:(( �"8
��0�f�FS�,��1����Ձ��Ӽv��Ǌ��sn���O m��
�~��Kwf�;ꄩg1
���}���c����=
˪[U��'��������Ifff���w�g���]��"����˶�ٔڏ�d��H�����Ws��������m}��.�c/n�j�'�N��`	[=%�R���\{�����#�N��Y�+���-����� ��A��9-lʹ�՘c(s!��/��re������Np�|0���3VR4� ��i���ͬ|�Zؔ4?���3qp����2�HX��5_Zl�C�#H�L3��:�9���i���<	��7�2���Q����5����H���%�C����I�R���uh�!J�	<��#�+�s����V�}�h��d�0�)�j�&3���i���!�ѭ۬+�����3_�s��ן����]ui)�@t��!bI��BNޑ7� C�]�d����)P
�eB��t8��@\Zy���j�=�: �0��T��+1���67�ࡌ��f,�qλC6xK��O��L�8v�P=o@����"dP�K����RH
�'	a����NX���Ռ����#W�x�u_��մ��ݮ�����eԶ&'<��E�u<7��s-�?~�Q4{wT�D1�y%@�٢�e��J��)�G�/GF���p7w�HG�?p�ؑ���a�^u�>��2���_�ڷwx�;�G��Z�g�k���{*�.Iөxi�� 6TVc�#8�C͝A�:Z�2h��m{BfS�Q �*c��1����J��B'��Y��m����rԙ�pǒ=[�v]�wΚ]`Wc��̉Ss2����\C	��Y��FpŽ���$�&]z�L���>�.xu+M�u!e��(��F��93/_C� D�:嚥l;\]�׉o}�C"�v�3��'�Z�3- [���#���A����s����$�|jy6k���Mȯp�2)�U	T���ȠX�ao��@Y�'}���A��rKfͳ��Z8焗NX�*@"��2U�ϊ�]|G���%x
��)-�gR�J 0��*��M#�R	�J������M4�LQ�LcB	|��=bV���B��t(�v�Z��`S��k����p���O�Y�>������n��{�u�=�~�:PK}z�3�	Ɇ�iJK�R���E�<�x�9���d�6xSc5�l4��!�Q<xc�<
�t�֧?E�t_��P��$3���CB�ǎ�Ɠ53Z[���Wo����s�?]u�翥n�q���W�m��ڭ���X�z�7��n���x!k4�:/ٺ�o���㘆�!���c�[���YJ�����8��=��\#_d�� �^p�6�Pz��f��������W�Us���tF�/BK������G�G�R�&�#_�&�$x�]�b�iu�O�VP�����9�� �R��>�$��>ǿ�s[_���;�]+��Lsv��z�;i;ڙ
U���a�*m5�u4�UH���Ǳ��~���, fWl��H��t8�����8"4�L��4��+�놉1Ӱ�x�Y4E��56���x�k%��i�V?v�����I^G�Ħ"�,w ��92w�r&<�R��g�:{52�l����Տ��!	�����N�������u�u q���A66b}���f��;xm�ǿ���cώ�x��1��Şa%cs�BB�`��MK��������"�UVUVVU�$����|�^�xq|���cF>�ˎ�Ǹ `�1�<xd�Maj?Cжn;r�l�w/��A�_L���C�i$o{LȘ*#�����8Y#nXG`��LpĊǭ}b}TyAFG����e�Rf:/���'p�š\8^A�,�A� �X�69����3yڿ�U��ާa�glz=옝%sqJ���&�9uF�, �@4n����`W^�Wuυ%�^&�y��[��/������|���Ŏ��?��P���ĭ����V���bO�j��;�_㰯���3K?Nʍ���ʤ;w���S��詓Q۝uzq�kǌXZ8�8{��Z�#�Ѳ"���sN����+�usBjM�Mc1:�֊ԫ~+~�5yh�2��l��L{��9��5+�L���G8d�q}Z���p��L�Y��'����76qk�ԫJ�i��Ѵ�%�.��: ,�t��c=>l�8@��f4�i �q��V*t;�[`J��$�� e�N���k��5Ҝo�Ȋ.y�6�Z��򩗽1%_��G�@�Z��:2�M͐�]$)p��x�o/�����_��h�z����Eğ���"��E�r�u��S�n:��t0<w3�yNa��$���-��p�Ӽ�*�@�SQ��Nu:�D�R`66��3�Y,�$B�5T��Û����D�*���э��a�Z��5^�ˉ�\}�\��I�y9�y�'�W`�, ��(��Dy:cTb��	�Yg�� ��)��f�l��°�x�ٙ�G�������z�=�x�W�� ��_o�:��G�c�ħ?}���E�4}��2�g�5z�y�f�gϽ����3U֫��m+�YNT+�ʻ��X��Q?J�^T?k��v�~�l��x�4l,�$���t;c;~ 2ë��gz*�[���ǏBh_��b�i>�4q$�^7)�*Ff-�Oh
�5�E:�i1M�SO�}@��",�ڱ���ʵ�ǠkmP��KQ��ӝ0%u���������\�7�*���FZV��i�Q4al�t���$�"Dݣ��4QӔ��eI�Ԣ�Pz��,�ݣ1Q��HRkJ�җ܊���v�{w���06�u�Ԟ����x��JGRH�C4Mw#0�N�ĪZ��Qj���J��,�z��i'bT#�`1ZG%<�*Pk��j���LG�G@�%�mZ���lL�^�A�����Œ���
�B`LK$Iƥ�)����\E���L�ע��R�T�S��-婝t�$?4D�J0�u����:��E��n�q�kX	�Iy��Ҏv�4<$mf�ê[ü����w����}仏?��o��[���6~ç?mU7����ݠbj*k-,�_����6Oi'�9���*Z�W�铱���]q��K�])�Uտ��S���=U:C����vUHz҂�����|�<���W�T6������e� �Z�p��#��;+n�*���i��%|��������b��p�-��
J��bs�I@N_��� �*7��b�Ͷ�8���ʒ[�~	��\}O*��e�� �C��.(94* �C3��&�y������lַ�8��W[4�*�J�{��6u�j�>:�l��ٳ$vY�Y�k�6� �^���8}2s��ä����0�fw��M:-�9� d=T��Z�x�]�H�-�s�y�-����87?�ַY�����DG��Ӝ�<N�,L#RAMNN�������oH-T�	{/o�`*iL���W��m�+:;��$��͍E�l"��{��� "� 1���E;vNe�Sі2�_��|�e�>˘^����\;o���*���׃u`X�4̴o;�/1��#Y7l�9�(��!q3�!�aS���RV�Չ��.�˽W�c�L����׽�fy�Yw���8Q��M�2����.�?D�>��ԭ�?3�V}��=H�G9�}ό�B�I$��t��3����J����0[���"���:�!5���J�c1�2
���׸:�f+��Gm����-��_�m+s�����X,�FS��F���L�V���G�}�+>y�����o�A3O��	��[������qnݨ�ޟ��g=z�Wf����'GE������������-�(�S��u�)��}��E噑�Q8������+��p��(�g󷭡��PѾlt�l|A�����{ܨi�4���a.%<�t�Z�w�~k\ ��x,z��X��4E�"���S:K��)�zj�*k�%���4=��ݓx�
�>5żvL|'֨��9�A�I� �F�Q�@����]�4F�h�}�s�nГ}�(4x���&oz�����p�C帾�'i�j���k�A<�oԲ��h܎���eS'4j:�;��R���Z�@�����fרh��Iȇ?�[�ڗ~ڹzz��~���v�q��� r�Y)ϫ�����~x�������`����x��~�,�rǿ�M��.3��P��o�X2�
�I�\�骬���Q+56�P�4�/�@ZX�.��p\�r��@�&��y.d�YR𓒈�4Bm/�s?��^6���,Ϭ~��4N4MOƪ�Ӝ�GK,{u;�~_�I�5qC3��O��Ϻ��T�=����w��f�/:�i�9�V����=,9$��}:+}�����6}�$��]vi޾�'�	�c�4���u֟�t,,�j��4�((:�Ғw3�	����'���P'ؔ�T�P� U�&岯:�!�:e�4�:�
�[t‑i��������d�A�iK�}���9k��P&���j�g$�B�����$�K�3���-�hJ���Uxr�]���G�dg����K�(�W��D�HYD��n�'��/�}�-� N�lv���2�٫.7��3~�����5?хw_���_�?�����c�JJU�DU����E���8�̶�{vr��w(�g\�̧�G�,�6��!�i�y��l��+C�mk�o�o�l�Ȫ�:���hs�0��������!��R�uM��2��(�L:Bo
W�	�'R�U9�?�V��G�㢔��SG��x�V�����d��]Q���"�!�*Q��j�l5	X;���hv:�-N�qOG�	��q���NM��D���q�|畯{��W��Ӵ��X�߿߻�}��KU�K��Ɖ������ga��s���Z9�뉈]&g���8�O�%W�7���~���i4t4.���h�6q�u�#V��������Sk���Ys/j_1Z��1���֞d<�ۺ��%�n��2��Y)�zq�h3v��#�� ��DŤ�:n���I"xb��%N5ֿ��]mH]���q�����$@�W��B�<hc�glӷ���\��ܼ.��	���\��x��\T	z�1�」ޓ:ʗ�r�E����2��������K/%���|�V���VՋS7q#&p9��E�?����و����ͯ�7�Y��z/��mv���d*�Q?�S�p�ѻQ�Q��Wi����#U/0=V�C �P%BDPW#YVP�mI����L�Ѱ�ݷ_ݦjCJ����S4SL��%�r�.w�Ա̫J��0�?�� �{�	sjN�R�6�e�\r��79�gt�UP��G��/l�	$T�ecM؉@!T�����:�wXǉ5��K�`�c$k<�H�)��نZ.o0��jn$?ꀅV��GF8R��K;��w2
��3;��7���[�N�W������K���f��{�[.W���K/����8��-q9����IB�DQ+pyg�ƛZ��\�2Ȕ�c�D���9��KN�w�S�#�R�r��>㆗D�r��"��hdŗA=6�h^A�q7zI'�FJ#V�ˬ���3�LZ����	<��O�t������P%I�G9���*5�2e8v��D������2�o� ��x��a��@*�Q��v�`)�j�7l/vٔ�������h��3/j%=��@Q��E�V��E 7��^x��ޙ�RY�IS���N�����v�hV�}���Cq�#��/�S��K�:�W���U f�J��T=�t!��m�8�����F���|R��-eD��Z+�d�i��N�<#ݥ�!�8�O�Љ����7i�̜� '��(�:zt�&p ��>�X]h��ei @R��f���FB�g&(&��H���@�ą>�Ja3a��Ѳ�����&�L`�E@"�n`yN cW��t�w�'�E�����Z�Q�y�g<�zT��}W�y"�F��UO3F�{�.��Of��~;1����r�FV���5�z��֝�R��7��H7}��KF�V["��8jAqZt[0�{=sޛ���]p�qE�.gw=t���^q�5�0J��s����E��sOe,�_q���ԉ4�n�{$�˼ݪ�y����S�+!�^�Ȋ;#r��TNK�6����+7)X�DD���O��
0�ֺg�)jh�Z.�&�HR��]�n�x���&*�PBMh}N��;�`ҡc�zKp9�@��;!)���]���.�t��qN�J_�6�� ��`�"��|cI*�G�1fרB��c�`za�����?yw8�"+V���V���-���e]l3*y�6`.`�HTS��8���9 F�ԟ��p���Z��?%��I���-@�:)�J�Z+
'�m*�c'J%9�u]+�M�S/���ҟJC-fwʷ�a�M]��R�ɮ)�?x�"��UE�4衇T�F$���#d�� i`4ʣB&�7-������y�k{�$+U~�%�ᳳ=�����s�L��sӅ�)�nr�6~��N��<��{T���q�{&�
4#ƊQ�cXX(V��
�&A(*c����x��!���y˴ܮ\���n��;.��<��oy�{O�:��tD����9p��lS�ۉ�_��[����7̠�7��P��V%̪�%ԍ2�Hl"�˺z����d�o�v�nE�/��v�LS��(�j��*fE��Z��nC�vwDv�C�ҕ^���S��@��r~2�'I�5��i�1����S3�=�<M�P~Eu���'4���;;ERu$�.k?�Sܭ{��	ĪEd�t�,^$��������9��|�M+����,�Al�>�@��
�3Ld�dgM}����)ͷ�)8m俕�˳�͸���I�N1�:Z�,� ��r�8�H�+�1�[x��@U�Sʄ�ls��"�* ���O:��;��J�k2�渊�/b�A�4N�O�`tH��ia5�|�&k�\9{�+�|��Mr�}�e~�P����S�C��`<H����.0NJֻ��Jj��m�}��JN���`��z����W.��DǄo#gƝ�$q�y% =� Z���z���^��o\�h�_�{������6���=�M��w��4;mtƯ�4��uT.�S*=���]�O\�I�@ ;ڃ]iU®�<�Dl9��G��Ӣ�5A��a�Ep(��Y���U�{P�C�4�=L���J��*]�����]�9YX���<��X�9�F��(���<�d�t�E���ǏgY�8>��7�+���#e;Q3D
�@���Ӄ�7c2U�I�R"a�H��2�/�鯩��f��V�K�Y�����U+�He�UW���������c�V��=&E(��~�*V?��B@aċ������|�uS�.ll��T[ڡ�N���`�ĸ��t)Bs��x@�Qc�����dL�Llx'�vM=!���hoz��}��O���r��\,D��֠<:��)�I��$�(ZϘ��y�j/�B���'U�=nP�	7ɑј�=D�3��5�T�(�m�ܡ�1Y�cu�F'�ę/������F�����z擷��[v���8~yujO�CT�B���N�9K�����:?+�o51ׁҠ^��2)3"$-�vrdo�f�&�t:�؞w�ד���F:P�nۊz
i�2��A
1�a�T䥽��?C.��=kw�ѓ����5���z� �,Cu���$�%B����{Wrom��6����we�DT�a)�`��27�u�>g�O@���������+w���HV`�<��A��@�hOK��%5�^�9��"0c@e��6�O�O���Q�5�"H����y�;�n:�d�[*��d	�V�Y?x��s���K�D�ԏu��- Ī5N��$�o^Do���]��s�̝�W�9r�s�?���v;��~���.����i�x�w��FA�@�ې��)��B,(E)=e���[�ڐ��窷����0�9�p�EJb�K�\a�d�B]��=�)�=и ����<L���|��pɢ���~п�ػ7��|��)��p��8��c��q�Y����z���a`�� ~�؎��ۑk��(�Zɐ����F�����׆6�3*&���4$-�#t�Fm�!����e��=ԫQ�a���_(=�Ww�_<��7����i �z�":w�'���Cj�8�ڏ���=�(����<2���;r���J���z$n�%�l\��3C%����o|#��-�H�7B�#U@
�9[+E���S�y�bU"e���qO=FX��"g:��鹣���`M�@���HԹp��X	.�:D�!Q�prp��/��9MT>eV�2۠h,�\ń7�5ݔD�@�J���:���&сr����34U�"t�f��~�W�x�����?&�=T�/g/�a��qv�:�+��7�x���~������zf���tʾ-���CB�1���Pb�W#dPC�z"U�;�Ū�v�/���o] ;���y�������쒓����F?�8w��k���)^�TVyF����w�K|�o?~<)��KS�^���zcJ@JW��ے{��	��Dڋ��(e���ϙ�{p��M�G��"�D���+�=�N�3��w^���ԯ��F��o?x��}�`�92�����BO%�8T��Ih:����ԃX��'��'�+Za�7p��X�������0�.C���7é#]4h"�pɳ����bK����P�-<x:ڏ: �~�u=۳������4�L�ʖ��d�Z�Nƀ��ɄpK�"��Wz��UaT�:ˁ�.m�D��K1��ZQH�"E���7�_���9��)Z
9w�@�f��6F��YTeD��#�;RU���$yH���k�Ͼ��o8��`O��K~���G�p��;w���=f��%b<�f�b<pM�>l��O%�TIٷ	~Uh{peD	 Q���\U�1E��T��
�	��V� ����IZ&�%�)-v.���{��CO}׵�G��µ;;�o4�/Ȳ�;gH��rQP{��)�+�(f��@�:�3��
߻h�.��k�'1(v�����W�{��w�]��Ǯ�Ĩ�:x��ʌ9x$���sȌ�3lf���v�o������ h�w���b/�>�𿲛�U:O��_�������v�|�R�_}���l�g���ׂ�hx!N ƨ�'�$$�.1i�]�nvȋ_�Ju�>�\wc��d��>�U��p�I�u�\�V*�8��^ú�^��W���<h�࢓"	�p)^R�t�]w|��x28;�$Ij���c�5���@���I��SLl���f��&9U}����)y���O:��M� �FFU!�
�1�Y���C';�7�j��O{��(ݿ������w��/v�����̫��k�+���'��M�]T�3�����c$����5��CDC�-��p�e�����@'��v;�����/?���$"i��t���]�&i\�F����b�W'��=���zOe_��A��G\S�!���3� 'nv��3�#���ˠrs�̽��9����:U�ۦt@_C:���j2`k/���3N���"��K�Q�CvEbh6HD�4���d�ÖM�m�?�`-�Op��4��|hW�`�ig<�*7����i=�Z���zi��c�V�漐��N˗�a*C�9�y�WK�����;/�p>�7~��i�^J��oJRQ��FG���
̻	�2��a��q���"�w�*=���U��Gԟb�!����f�m��g^�r7�,MG���Ut�K
ˡ�Yݓ'�)}�����B��@��F>�q�>Lȑ�,�,\"<�<>��ы��Z%O�(����H?=�$zѰ!���1��b�,N�Y�2��.9���ɞ��%���Y�Ơ���S�����':�����lp^VKÔ'���'�Z��R�v\�w���t�����r��Ou�����6կ�<�\�x]	���S���������0�iF0��5J�a���#�[�����������(���0\�8"d�^'���@����(L�-T��.�́mcҾ�����{2:NJ�i�+ܹ�Ř�ZVQ0��5�����<Ijӌ�͔.=~����]�G|�]w��]��Cӥ`^����N�q!����r��#u�#-�/~^?"��-�WB���7P�DC�J��`�^${ά�e�ً~�/�x�{.8�1J��=ן��w��+U�R�g�sww?�'?�;���~�����fZ{[[:;���� ;y�T���6gjk'�+�G�*�s���;���8J����k��:� <�yAg��6�A�Ьv��4���~@ϫ�T���i����]ic�'��-`D�{^��̨�uhn\<V�E3f�9�b"�wT?e�UьC�bDW���a�v$)+N�i���Ȃڿ��O|��n\���ܜ��;İ�~�s�'�g�3�ꡃo=�W~>�k��0�5%�����l�L�����,c*X"��~�Y'�_RL���k3`k�����E{рl�|�=��zdf�'���Zs]푘�C�iL�W�RpĲj`�g�AQ^��@�}����,qȎ=w.�T�w?�ҫ�����>�9)��I��ʋj�Nn(oz���Qo�I��cVc���?�_L�Q�;W4 �#Ydr4n{@X���e����c�/U���K19J�޹��������?ybgF���NR��fJv!�)`="��������%r�V�e���>�Є��m��Ɛs��jU�k��J��B�XsW��-D��%xB��q�C�ڢ`lwj�FFt7�:R1�0�$�S�3���G���M����pG�-�nz�d��m��+�	DJ�'=��/���"�������04�~����o]�z�����O���óϯ�|Q����0~�5�܁گ.�/<���,WL�h���!��M�fg,����-���Cg~�U9��^�Θ$�N٧2��J@�>'K��� u��D�ޫU,Z+��.�cQ�=^��_��+�+{X0�d@�+I� $�':�=�"��tv�}�2�}���_�����#�De�c��!�.ٸnV9�!��T����$䃢�b¿s�y��G3y���űI��rX���+V���_~�ʺ���o>u��k~l����~��E~�/[���S��򞬽<����@�C3�� *a3ӮrZ/��m��H�Z���Dq44!O<�Є�~�`�#��$�ht{�:r!1�8��}�A��J5Ȧ�LEL�� ��(C��Z�zme
�|Yu�T`�M��Q��LCx T�h�~�����N5a�y���0*U��c�E����)Y�	�����/a�xJ=�����rN�DR�qE��(eƋ,dc؅�qs��3cq�)�Ӷa$+	}͒e�m��_�@$�����VK}��'?�d*c�YX�8���3�!i����\�R/���rε�8!	F��Ą��!l �$�Kz��gw��'�Y�=t��-���w��W�֗�����T�u��K�ob�
Y�&4�i�uS�m�8��u�X,�����၍n0�*���m����πC�QRΤ��r�r�S':?�&�'����q�R#i�p�(�:�sfN4;�ͬSq��&_�5��G@��XWgrἕ8*$�ߪH~N]c���d�t�E���x��D����۟�b�HhLd+�Z�_L�VB �d��`��x1Cj�I�M�;.%fr������ƢQğ6�oI����z��R�,���Q���{�#T��i"A���9r�SrU�I���-v��^�b������!�l;��Q����iv�)������Z��9e�$5!����In��k4�7��.�?�3�Iiˍ�D�vX��f�I�F��mpWv��A<�����%|�}��V�;#.��'�L�~�{�{֓��NS�����=��E�ɒ��\g''3$��CP�嚶S@ౌ���E��qN��ɪ4��9�5��T#F��{H� T��S$�R��/���Dg|Z�}���T�����8�����(I���h��P�Wu�����X�3"�.���&���Q�#����q�-�F\2���,�h�?���"��'���{�,��3tO23'ya@W���4�5\<��:��rʮ��ԫh6*�y&@֢~B{����1n	1T��8^:�k�(#C��jRjT��1x����%��CR�����������C?�s�,g�V�1��ܕ!%&m��5���룳�o�E(:,�mek���y�q��Jå��"D�i�2 h���9wXA<1�LC	d&_�Gh@G�|�h8��Z 1���8PVU��2G��$�)u$���4�����N@b`t֩<�yT��V'�h��h2��=�/�+���J�WCFV\�ex
j�;C��=�VA��z�Xk$ �m���%SJ�]l#��(�xR'��� �t́�}F��}�P=��F��I�a<25��Z��6�A���@���]�!�U���.B�w��L
�f�Bݼ�J"`���l�n�V�^@<�u[/�*ӕ�OY�gC��h,*������D_ŕ�s`\��=��&Ф<m��"�$iJd�dG����4� ͹	'��&�Di����[f6*��o��0}R�z]I!�\��y�l��<,�� �P��+ύ&�L
"�PcѠ����D�0ƬK8f�O;C*�|��!��h"�B�f���՞YD�V�Maƴ��{?p���F���EH� )��)"Y��Cz�\%���q�,��q��%e�GT+im ��	�n��Q�˂���u5sb�j$Y��:�������&���M����6��5�D���d��2"vbBt����1e@�*�I��쓩�������|S�$"�,4L[��׺E�1��".<�b}G�����MA/�8��r���nB�E�fZ�T�o�\�į��g���-����(v��r�Fwi�|�:��|��GG䪚lP���Z�K����6w�{1'+-(��|��[��iH]h�XJ���
\w���0@i*�A�v�Iõ�HUhօD��\�]����I��v��u���E������j Z����k���-�ҶR(8y�*l�1T3bP?�yUx�ܽ�D�$1u�Õ�݄1��zde1����Cs`-�Ar���ɟ����@�2Lig񫁂d*ԤfX�'>��.��ѿ;���F�
whqL#��^�=�j?�x��Tk�I(7�I�&�$�r��e�C��3Lw\dkۘs���x�M���ψ�~��B�W�g���]Z��	u"(ӪON���OԾ6�:x��U8�099ܡ�ʂ_N�S�2އ}��A.����e���#<jR��c��vV%��`H�̉;�~��<�G���VO\j�~���d�m�?��aܑO����9y����ԃ�� {�F�ˊu�h�����zR�iF[��x��3��#���v���ER�I'�Th������P�<�9���5ƌ�G���2s}�C^h&��Vow<�S��I��#2�ȧ�N<<�\�e�D3�3O�_�SL&�-D�X��&:��G�|�ϲ����P�V�����ի�lXm�=��K��sr��,_1(�ߖ�?�Y�X�R�jhj���oHr�0�n����+���E8���뎷@�
*4S�L�W��j�R�*D����yzz":�qs�YB����~�� %*�ʚT�:|)O��ZUc��Rk:ܵQ1��1�OkiB�5B��:׎k��Kq��h!/Q=V�y����S�1��J�|��y�Do�t�_aĂ��g��Z'��c�Ȋ��H�כ�:�F�����z�-���n��z���K���(n�J&G�)�SuI��yjz�_#.z#��.��Z
��4�"z�a��_��B��A���j���]���ښ�ѩ�D��1�������ۥu���:���H���?���vA����86�*�3-��l�@��E~I!���lV�Z�3�{���R�Se$����%_��M_3(L��¼w��1�ZP
t���9��]��{��η�G2��}R8`�Y&�E��2�/7�E�<OH�?=�hܮ�,Wﴰ ���DO����܆��d�,[jJ#	�3#�� 3��0��h�����J����ApE" �-�2fNn@Ȇ15"5�5�_MlѠgr5�}�o�'-!y���s�B�%ªW��:k�&���]��'L�oh��Y�.i�z��F)%%W�����/�������	�K;��U�щ_�TS,�sV�ˑ��V��>��q���d�t��)ۍBe��I���v~�ɕ�Y�!��81˓�b��u!:�Ǆ#�krdє��ES='u�"ۭUgV�$�t�T���ד���߀K��٭��]�M�C��a�2&a�o�O樚�>/����=���l�/�����,W�L�$9��v�#�;W�] �B��7q,Tq�L�<�m��c�g��wL�E�c���B"l�	k-e$P�:��?I"�a��c�M�i�9��c�� ���Z仏�����Y�<�np��}���Ln�h,\�扔�+J�20�I�X����`:�i�됋.D����:[[���5蟶���܂ie.
_�J[��g�q"�rق�a���&��.Neq�R}���:'s�1�3�!&<�*fr"�ThG)H$4'�V=���~���u�?f�3X�'ﵗ��z]�C.Z$�̓�o���noc���j��M$�V�.�
� K���b�*�2K�
ENC����~�����dr���շ�|���9��1�QQ�v@�-���r��TS2m�2ēi�_b�s̾~7:Q4��M��bŃc����(�+�]3͊{����}d%�/��u>μ�����W�US�e���U�>����P��huP�Uy��<�K��t�L�X���x8��"��Uy��>3Ku��gS��;���Z��<AݺV��Pj�3o�$Wأ��1G2Ǒ���Jc�~��9��Q�Z��b�|��u�����q�ϵ��.��N�Z-�hB�
��N���q�'u�Ϙ�F3YtMv}�^1�6F\ZVf��Jo'0��'�>U�]���sK�7{$CϢ[8�m<��QV�Zǩw�X#t����-��zC*��5����Da�nvF�Pq^���o�eX�>|4�[�:o�*y.����}�@o��GR�=fY�S�,L{Wo4�鞄QJ�8$A��h��3�V���a���:Y&'�0��U[���J����X�ڔn�TO^K���U�a{|���'Q��>Ւ�X�RG9[_n�{�r� �1\�<c�3���+�3�s�ź^K5����r��`g�ʺ{.�:��;#��� � Ú/3�F�rQ��cm![E�73�cM�I���j�#7�@9w@�U�?]��#T� 9q94� 7u�Ί\�}��l�Ml�fo�l}q��c}��	ƌ�<'k�&-�X�'��r.��W���F�<��NN1B=��gn�9G��DbYn(�պ�v��������ߍGXޛ*�Px��9��J��n9�U�X��	�2�&H�D���ۈ{~�Q��߄.�r�YH�Fs�J+�~�oΘC�z����ld}�P>R�^�[o�瑈m�`f1�7{�~��n�D8":��h�|�%̞�������R'$`T{�A?�I�Fd��A��ps��l��7M��#!ۀ��e;�G�D>#i9��U�~�^�hzӾ�CQ\��a�:eb:���Ȋ�6�=�6�W���H�p&R�B�0�(6����0�0����=rZ<[6�f���(6d$�8�j�~1����3��gd��@\V���8*�;:[8I��p+&5�9���N�~��I�����4��ba��9��c���V�+]��ub���h�M���h���|��w�򩌻֫�CB��8F��鉛H��S���T]�s�ly�y������.}퍣0v��Z�rs#�g�="y��V��r�w��1o�ڼţ0c����V2�M�"t���xJ��n�:H(�F���M5�ʋ��z�I�W�`���ڸ�����n!��Lhoun��@K�rlEL��Ѿ5������M�+!&�M�*c�hFK����Q\��6L��_,�P�T�=J��S.pH'ě'[aD�w̐h�I&yg6
�>���Y�'+/�>\*���6;����q��}T��f�c@~�i����s}��Y"�4�B*��#(�}g�>Ee�3�Ǐ�[�TJ �q�YEV]�G�蜙�� ,��a���
� �U�~NH�*َ4Ji�=0U��~e(�ӡ ���Zug0�p�+�b�.R}b�c�H�wH��aVvj�~t��\����SlƑ��7�����N�GI�<��Vd�_2Y��ʤ�K��<-.�1�j.	R�y�z'�
󝪯6$�lg�����٨�Y����D��Si��ԟ�%8\��%*�j�]�)�i+�ʉ3z��Lwn�OHF��P,)�R�ꂖ`LzK}m�8՝'���1���)� u�j-��5X��;�c��k�8��Z�t��{V/`�	2�c��ݗI��I��T�u�/{�Z�(&xe�r@�pX����:x�̹I涓!�N�󷓵8iq�1����ǳ$;���3��;��Z{�(ieҞ_4Q��ЀD���V|`��Gb�*|$�������w;�P��]�K\��T .��%iC*B�0ժ�z�֗���s��M�q����b��I�JR� o��!ˡ�#�.s+s��0wmè=���m�.��@��u�IB�#.����=vg ���4�,N��Ё�=\0[S�0�G�êB��0Q$J��h����YEr6W-?ND�9��O�lS�f���̋�ӧ�i�^���p����))O��Pj�yi�u���d�#S��9U��b���RV�M��i+G�?� י�*[1_I�/�.N|
ҩ��n����N���K^&��·j5Z�z��MV՞��.Iͧ�k���r��f"$��
p�1�u�t�����~;���O������j���럵���;��y��C����Zꆏ� ��)?�(9�]_�<�\K���Mڥ���h�Zo�o����RD�Q\H�	Q1R��w�%�ݾ��+K^QrA�����D�^'���P��Z��]Š�5���a`S��LX?kĵ+������I�8��nɝ[P��D8Q��6�L�,�"^�y ��;b9�j-�9�x�[�]���R圖��
	Qk����*�8�.,(���=j�4��0ٶ@"}�Pe&�����f�M��yEEne�����z���F����k6D�3n"h��!k W�<��uD7�{'o9����~��Qtv��*{2Z5(��$2��f��d:_o�v�G�)R�5�L��(���P),N\ ְ�Ɵ�3���ZG�WWL��뼤�@0k���?���~PU�0g��#�RB�=u��Ż~x�q6�p�Ҝ��ҖI|�Ut��7���D+����W�(M�ܯz/o;�%��F�$}�����̙1pk�e�P��#�句`!c�J�
�mT)��u�k6I�G�H٨?�R��w��}�c1��ɴ"�93�}+b�v�<������e)5MS%V�ﵚ�������^t��޴��ݠ�ϞQ��Yz~���uR�(����"ub^�p���w�ڶ��<n�XW�q]Z�~��62�0��ӛ'�O�:�	��8�����"�@sv�v%����ţ^�������ݲ���y���f{��L&�V*��aó�,��kJŤ���c>T����R(J�q6���E�2��M�㯔r����-�T��:lG��-O�E�S�>��ʸxڣ�]��������?�؄�~����v��>q`��s2I=�<���2����_��+;��+��+;��:鋔�$M/l�ݝ��ۏ,{�n���~1]8�󋴴�'Y/���d�_��'D��v�c��H�QG,Q���l��qţS5��3 fh�����w-����F'�w��!�j(�c�}��u\,�:��r)�y��Lb!c_j���'7>��p�L������={�%�o�ز��y�L�!a7��圉�^Rz��\��`����"r��y=��Fח�|N��%���ƻB�
3j�m�H��1�I6�X^pٗ��z	ɋ���`���\��6'�V�	��c�S�I����p7l��eG�;�ސ�?sK��+�kGc�������1o�XJ1� ��M��a.�I-.$#+�1V�����<�F����(�Ċ߬�����Q�qŃ`q9�.f񷞌o��܂�h7���=��de������r��DǳY�������3���'�����w�䟋+��=V.׳��J� `�zI�Su/p�6	�t�iU�`�*�����3����V�d�y�eY��p��-�Df�!T1#5 =8:����|��Qץ�L�� ������F)I�J�ɖ�e���(ĐR�ρt'��
;lN���{܉i�3��H�<�i������3���ۋ�{i��c�[4w�2Gg臤FM�g���H���T0��{?���wSz�wƮ��{,K#&y`����Ƹ=UH�Z������>����#�4�Q忓�y�e�
+6�LH�l���|�d�X�t�������0�>aCg �:��Z���m����\EN)�+��6w����O$�r�D~�_&q�֭,�5暖T)����vɿf�3%������ܵ�me�\ҍc��!��7DNиƩ���@&���j~���7��Q��:���h#P9˼*����[�~��Y$]q^�Ӈ�) m`P�"1�ɒ�����KI4���W-'_������y�b/yS�S�0���3��с�M~;&�gV�NQJ�T��/�4����eI�Q���"��c�{�ǯ��R�bڪAx���q������1G/�Օ�S�}�b�[��Jvdn�"�a�AtW���}�>�:�\\�D����y���/,����:�&B#D�1
�۹Op� ��[<O��X������ι�sk����<��˧�@K�3����Aν��ng!w�qӌ'�������MW��.4߽��{�+~�J�EB�a�6%`�J�E�,�:�>Z�$�(p�@m8�P/�)�b�����0�p-p/�u� �0��B)XIi���8�}�}w�JF&�t���g�Ev�vpRR�CE�0���}_��-:nܼf��#�'���i��mh�\hK�] h��_��d�n/��O^|勿v����>���ʍ�i��b&�<��Ԡ�P�@#.� i�Ra�sLA��ϨM��R��J��G�-�tc?�hS%㊖%Nth�$t�#���09���`:D��Y�a�w✣��c�P�z�5;4e:J�~|֖,�A�.��	r<�����:�e;�˿~���T"5��{҇0V��bIjKy���߭����~-�:���/���q� �����;b��B���b_����m�ב��E�8b��!5#�*|�Gd�R!*�ɷ��^g1J���6H?�z��'�Q��:)V�5P��s�!�(2F�$�_ɱ\&��Ez�NZ�����xd�����A#�]�7]��O�*��a(~��T����q��2U& %	�:�X���9M�z����S8�R����՟�h�]��z�E�y�|��ds��]�4�r���DL^l�l$�P����fD�Z�!��t��>~�Y�Ņ�W��s}/�s^��� @ܽ����zV0�fffH.<������]ǿF�����,\����Y�=�\��*�%(�Ib© ~�G�C��3���KopQ�`����?��zf2��r����;�h�y����S�Ϋ���<�b���iճ�])�5�Y|���B�v��f��-U��3[�;眙���X���̩�%�Fm=nI덯l�n��0�`����Ku�����RW)�>�8��s�c�˵�8��Z�ͯ��`GP�ʤ�����(��P��(�ɲ���,N|��x*�]m�M��1&t;2&��,�DS=g/X��w
�7��ը4�Kp���r��<P&�ҠX.*��0�ܖ�B�ן��:�������-�����1X�%�l9W	�u����%|���g\7����,����Q�f������y|+<g��,؆Η�^`�9��/3?�#�|�y��,|�� �t2#/Y���[p��`"z�V�����ܐ_�<�:xe�Ef�~��?�Ȧ��:���$���te3�S���]�{�g��P(�Q��A��n� ��A�4X����u+#�,a��#�q��yl��g@l1c\����$:4A�q�f�Z��i�wd�`��灊�{���;|fX7E�e�$�a�{@���vPg��3g��2��i�=o9%u�+2A�T㭠�g��;�:$�69����q�`��.L?p�x��o��k�1��@(?�z?5S����I�Z#I��,Xl���?�w;��T`���m�aנ�v�\��o��F�b"�&|��~�Eo�~R[k�tr߷�G=δ�(�����ч�������8�]������V]�uU���rJ���fv��� ��Z�ŏ�;3sKͳ�:t�+G��X�/iLi����R�o�D(5��1.��D��W(�+��S�<`n&.����l�HC���0ש�	<�%���9`��˃t�2�{��j�ԁ���n�"$Z��8��RX�-����ZG���A )��8��g2(`��db��X�<�V^{<Lވ�%+�А��U��(�P7MCŧۼ�������_Y��M�HD�s}�y
W!�$aa�[�f���K2���¸�|15��F�b)�Ѱ���G�,T
�s7Y��e 4��$����#����H��΃8�4�����U/�9�h,Ph��9�9q�ƽ0����tb-k�2�������=�����f���B��j�D��60�N�lH�7Jki�E$Ƚ���u��*����1nG�|1�_*�g!9���{���Һ�f\���p���S�~x���6ћZ�
*�O���,�0+c�ԩ3�&�«��v�� }ɵ}y/�=ʍ��K?G�� ��.����SQ��]{1�+�5D_n+2��i ��6�r�e��%�n~c+��'�4k�˦����A��Sryy��rkQCe!y�q�֬d!T������%��}�%����&�g-&:�:j�f�69Ɩ'u)��*���}��(='!�m�=�����A��q:��Z�� \�=13"�a~��`�5Vl�&k�[���`�W߼���/<�.���"АgJ�~���/d<0�Lɼ]��j/I�9�M�ABڙaC��2Rm��ME�U.�)qN�-�YG_���F���J@�_��I�Ô�򠸾}��a���<��mk����ϳ�hϛ|0h[�Rk�$&�B��+�c�Z!���7�9�[5	-�X�I�M��ETj��S�$i���ah��ٵ���b��So��Ru��Kٗ_Ƕ���.(��E�����;1v��Vˠ�u���ڿ�������y�A{�t���Q��P�k�����Oő�eD�~��~������w��4��G�~*�C���Xs�P�w	i�2�"���f}�6�5\V��(c�s.n]�;� ot�Zm3��=QS���<L5�5hR�xAq�ן��R=�Ԅ"�5l�������6˰�bwn~ϊ�dv��R�Ѝh]Q�ڒ�@�	?�6��8v��8�L����|�S�l��gl�ͫ�J����!�������7k�.�JB�.���\Y��dNt�L4��uݨ5G����㔵:��S���D�׸(�˅nr?��`�i|������97�Qkܲ�:��3�K'6�5o���3Y�vb�V���l��8]V�S��~�����0��\���v�*b�̩X8�_�c^�l��[��oik��FpN�����rT�>��տï3�����\{��$��ؘr-�����o������QO/��;��('I�e���L�O������֗�W�j�md݄]{2��:g�x6���?*���g[��\{�0�驶=�6��\�Ne����̣���l��GGUXZo�7��fY��Is?"��D��^4���=矿����']�m_����sp�mT��m���J%E�I�$�*便�%�8fk����|X�dM�~��q3h�k	��_������=]N���t��R��#qǂD�����s��P� �����EMC�	�����
jL&��odA�/��{��D��F	��5k% 9]N�g������),�@s�C 现@��>��x����nW����L�l�Ȋ��nשV�u'�����S �D���X���r��.��WA&�;vK� A�<x0����{h)��o�r�2!7I9���@�)�*�<U<���yE%�ڊN���t9]~�%�V��y�ُ�\*\V��zU����Gw2��f\~]"�гa"�Xt������u�]7��n�i�[�bF���t9]N��h0E�x�ή]����?�������v�9�(7Ѐ���r�#�3��]���i��_v����_;7�p�x���}�? /xQ� ����tyN�gۉ��.�W�-Ä�,�Gfgg��x�{��}����.�H�{6����1�h��5P'���_���<��?M)�&��
��%���r��.��
w��lV��$I�AP���P�5@ܫ�N�R�8��j=�~=.^��m���G�L�⺓��P������>xٻ���c����O}�S�={�|s�پ+ᵰc�32�Ȣw)x�c�Q|)��6�$�CX"�*���*���:eq�b�`�/Ѝj�Ƴ�v��R��5��x�������#k��ߵ�<�B�	�O������q@SW�X�H�q܌�T��t���ao�ﭼ���al/�yZ*�Ѣj���H� ;| ;E���:E�	��xG�\��{��^8�4�}������|�OB'�FQ|�Ȳ>7�ƻ�!ib0L�/6��*�5�zqP�Ͼ��%�8!6"�v3�}hэ*՛����`c����q#����|���덀}i!�gq�]o#�N��}�Rp�������v���8�E�?I⾙��.��V�!q�yR���)C⎙i8w� wdB���7��뮻��p��t��9���� ��gO$e_���lX	p�D�B�H��<��k^����������Ї>�۷�k����G�-�+�T���t������Sz�c坴����ěX�c_X����^�����F����z���n
	އ?��F�W$��7	�����a�1֌=�#^��7��Nt0����e뙀�x.H���Il��h�oE�kT��T*znXw:<�� ���g���f�{�%��ŧ7�AYk�#�J�u麾�d�`�e�91�~X*u3��"����6\fYi.}����u�� ��Hlf͍�.�6]�4粀x���'����o��믿��������Ç�����Ý�2{���E�zmU�v,'��|���Z�X�66�f��F�r��� �A�w;==�4���hl����e�~jj���m]׎;h���}5�|�vj�&�+��sjsx�������%�z�_�P�G$��N9�J����n�F}k�M߀��)PL:����yek�a�xX�Z�B�=5�������׾k�9܈�?���^���V\c�^k=�:�n8�׺�XN��6�S��oI�ڨ��L�n`�R���A����):Ề�����L"�X&�I/�zF��6k6�����;��{W�ǷB.�qu�}l��O
.x� �$�E�(�>w��8eo������w���Ǯ��j��ѵ�^{�/x��?��?}�����B$��.�L�&/b5���&��'r�|�����V^0��3Ū�x!!3��;�]�{H���:��w��m+��	%��*O�i�c�;��;8+��ĥk��G�[�mx�qKl��g��(��%@E_�1�o��@�ժ�vqS�~�x Z�ӯ��K�VJVf�˳���W%i��0�{T#c`d����dy��7#�3�_�6�Ĥ��o[�4�09��QC(P:;��uy}ۛ�t�~H�Ի�I��`ԏlk�*]/o��z=�1C+��^���U��=��O�����q��K
A���'�u��7�BԽ��"��e�&��	�٨X=�^�%q����/>��?�?�o��ozӛbt���4��c�]�$�����OUWW���43 f����K��?��b mXA��!����^;�4�#�0�:�v��CY�wm2��l�+�2)ٴesVZR�#һ�\`�`�3�ӟ��|�{_f�򽬮�|��
�]Y��2����=��o�X_�|��n�ʉg�=������+Wزڲ�;��+K����?���
[��~b���ߵ����/~����쏂�{f�U49(�cs�1�v�]���ğ*�,(Y  ��^��ܧ>���~�����~����ɑ�H4�XcKa�P�U������S��?O��q�r<��U�y�f^��P���KOׄe����(��翑��O�ğ��������˗/㋚Nc�5vRM\�tI<��#ɯ�گ�8��$Ap�0��1�B_2��%�9��<�}��gkP𫫫*�:���`"Z��Ye��;�x�1�O�9ئ1�O~�w~�y���p�������?��}��� ���=޼�n�n� Km��}�wy���Ǝ�N�Ō�F�ʯ��ʵkۧ���/��{��{6>��y� C�4���l0���q�'>�P��)��������
0�&�{���q9���x�p�����[��ex\SJ��}��Ȱ���2�6-)�Y)���y����V��s;+�)���1~�&S��rn��0�;�QM5Ƨ����0Ƕ��g��粄��yѻ{�|�t�ó��V���Ső�?�G��-�/�P�11�nwM^�~|�֚��0���\�L�+�?��v){���N��'�|r&���7/;H��+2������j��w���I���Ղ�w1����S9�)  �wȘy�w���o�fn�<��u^G��eQ̻=w��m���3��͹sX�s��m�\�����v?a�޸��v�����KW�b �tU��@ ���x1���.��~����ذ/^|^�{ �[�6���-��M,���s:a1h�#��G�ۧ����WVʠ��Nڻ�P�v�w�-�������N>,{�����ϟ`�c�$ݹ�c(�'�����#��1����[p�o�c�0Ǜ'6fΜ9��:8��c�&xZN�ܾ�Y͹?�!>�����ϳۮ����nz}�������v����ޟyu6�p�0|"%w�@�z>�>��fY2������I��n�������|�3v�۲�7Z+�?0�<���z{�����Fǥ�1y��a�� v�v�=��x��y�N���]����v��6�W��C�%`�эY-���(��(qr�]w������n�~�ӟ��[��[�06���ի����r�O�����H�O�I���&�;�n���6=�;m�z��_ߝ�;��}��;m��ENHp���{>�x:{�y�-E
Q���{�e/^�[]]��s����O}�S��!^c?�я^��������si�>t�ԩ.x�)����>��nĻ B_��{|����k�̺n��_7O]�pL0y�`B�M��L�[�@3��p,���?Ը=s�h�x�iF����?��̾|��Y��O^ӻ�����ޖ�ox�R;���S�<�pd)"��?^�}��/����/��/���/�⡏u(Al�3ǵ���?R|o���̲�n��=�rP��i���{�[{��IF�C)�-�s&0�V�u	 ����Ё�#i�� Sf�b\�����ȭ�/J����q"x^��Z��a�r����FpA�398:���q,�����/R�T^$�r&�$ڠ���7S
/�@��AI5)-ɵ���u_�B��]��IT�.Ǐӡ�,öx�(�KVVYv�?�wHW�������m�Jqq��s?�3�pߴB�����E�0�I,����q"������s�����=Q�ñG,����kc^c��Gx��螖�GZ�h�����x��q|o'���}V˽���۔���X��)/c.\ �cR����{����eߵk���,�H����8�}��ۨ����Xeekcw�ʥ!~�DJX_Ծv�����_��@',�e��~/4�s�U~�]M"B�H�{�s�A� t����=�Q���R��>j^���}�>�N��-Hd�F�yt�xЬdX�h��m����%O8֭tpR��U ���&%w���0����O� pǉ1Y鱷��39�߀��َ� 0ւc�z��_������J3h2�s�=ʌ�g�e���h��l��b|z��"��l��^�����,���p��C������6�<\�xc�;�_�������˿���_����d�W�^=��~��>�8O����b�<�ϸF
|Q�w���,p��ˊ�� �$����2�%�`��*��E0��!P�0��z�ILhM���£Վ�`�G���fK�(c�<�L�!Q��~�h��Kc@�|@XC@/��E;�o%�������+(@�8'��N��u$r�Gm��2�h �)qr�5���0E�m;�K9�S¤���h�=� *�f������Za{Ĕp�J�����ɀ�-\XMJ����� VG=3dD�=�rV���Iø	���br������X=.�5N���ۄ���Mx�1��ϭhғ��g�e��[5
�MFJ@:�w�N������R�l�2�AJ%�( ��w�ԩS���	V��	���s�����C�ffm��/��� @���ׯ��~5w��n�������eٮ꽾�{���d	�y^=R��hx[[q���=&S��q�x�����e��"��K�ӝsr&1R����9�+�qE�?U�T.�P��F�ǅ ��b����'����ϸ�z����!�"�����]�L���SO��s&a|�G�R����5��:<�����IT�� �Xm���pŢ(����}���F;w�n�d|�
nDD�=NJ0y�}V^B+�\9pO|3��E�,'������d�����;������]-���z�\�� ,s�\��:��{�to
�r���'�]�z7�$�L6n)�w!A`���r�� �> �+�y��������.6M:��x4���~� �|��_ޅ�a�׻ ��f�����c΢w��S�a�;���a��w�n�hg���~�9`��'�.�n��<��\��_����C�y���Ƀ�S��Ws0�3.�A(��Z,��#
��ܧkk��/I)�s�WP `�t��=���Sq��RIъDǱ���G�g�A݁\��gE�&e1���Lc��Ȧ�i���0d��bhY���"��^�F8��\ܵ����M"�)rr�i"���y��9Z�{��vZ��or%Ϝ^�;O�,��k�h8�|����P�`�9�1LpH�ޑm8Y��@$py�&E�%3p�a8y���߸y�W�+p~m��A'�<m��t;n�&���s��"�9�j�d��p�̞q$-��b���qG�<����ʸ	BªG�F�����6��c�(+�$����Mn"XY�����e�oR���l5�[��-7��?<v����Y]]}p���a�7�;����ٟ}��qd;����;�������>_��_������)��{���9jeU0m�17�h���� �Q��I�|;Y�NH�O�&ar�Q��N��׸����>�K�v�]�~ྏƉz��J x;0!�g(`^���׿�ҿܾ������I��(р���̙���s��璟��iD+ ���ko|�ׯ�x���GW�l�ٕ�`�׺�����<���q��\�p.�E N�w_��֕W߸��¶�}m��$3C��"V�>���=�6>�鬜�/�OH�~0�x�[_�z��w�\��=0iz7�Ol��[++�^���VZ�48�q᪣�s��7�n�}�?۽��؈k��u﹍G/^<���Xl��� ��0���b���u�O�|���`��^�E���@e�k���>���/~$��ݭ4��$d�=�o_y���|�]��m�l-�=�B�k�����d��w��8γ>k�6���zk��+�}�����x���������Az�=g>t�}g��G�T+�iFD�h+������o����n�<Z�����7o�<�}��Y����4���vwwEm�9,�]�!���Taw���t'��8���3�9��!�s��K�-k}}[���o����օv^z�=���\�:;2���aNB�&| ^�|����ÿ���ܹs����"<*����x�_��k�GI��o��a���v�_}��������om}������{��+=|�#�l?Ny����dC������G��}�<��W�����w���ߕ+��������G?��յ�@���%6��2����~�ŷ.?���b�]X@���:{���Ӻ{C�?�������i�HH8����㯼���޽����?���o~�K����_�>�����<����W�m!bjG����9�������{�٣�~���sK��Λo����[����?�m����V&�ܼ��֗���7�����փ���v��M��y�ů��<|���m����@�[+��������_�������ȟ�䭻�ڴ4Tx���������>���ܷ���oL{���P�����~�+�����?�ۆqb{>8!�W��Oc��~�#��hue�J`��Ip�̗������׾����я���n����.]ߗ��'I�����Ǿ�K�Zm��jJ
����ܸ~��W����9{��ޭ<�_��7����~㡽���鍍?zࡇ�����O��O�>K���k׮�gri����Ⱦ��/Pg��￟�.]�h�3�<�e�Ǝ��*v��Ǝ�~������o1�D��\=}�?�#7p���;Ϟz��Ir��˭I`M?�7��6׺�k���k7>󙟚J���/�D�{������� o26R�$Nٰ��R����Ц$����L���_���C�=�����7uaoC�����:c�_zS���'�ݩ���g�=���w�����X�Vn4� �#�*�~��G�w����z�S{��}�s���#�'�gm�ӎڰ�p���n�Hl��ɟ�k�'���_�k�G8=������� [�x�+������፿��r{r�����h������^[��4�O�g��tW�����������OMi�|�s��_�w�_9��P&2'�+ˈ�"�6�	�y�S���/��_M�{S������&Ġ�į`+��r}m��v>��W���3�O�����ށ��-�N�����}����t�t{{�`z�CL��u?�-���,���m1l���4M�N�3
H�s�t0-��Y���@J�	k����w���~���3�٩c��?�X�v��~�(��EǤdG��sg�v�]�$>{����=g��4B�G:�����\nn�]8�(c=����}��b���0Q�i��Y+^��7V�V��*q����~\|�+��t��OI3���4��/�;&=�y����~��S?�7����O���W��nmoE0�10�y�ju�����c�����aj�Ng]��ͻ9�:p9�}ֆj���n���؅�T���	��q�,7q��tD���8�W��y�}�Uv{衇��t��������V��|6�c+��S��C��_�p�ʋ/��j�Q
����2X�'��4���Yg�#66�Md>��X\��2���4 (�3��:	�ƒ���㝅��L;��E0��>G:��2~��ߨ �=�
o��-i���5e.%5��\�Ջ7+ ��]eI*�p>qc��+�Y�?�+�N�����$��^I�B�k6����$R�5V�ۧ�$M[pi5��rQpdG��(�d����j%	�8����@lu�M,#�������#��ʿjI�s�^��Ɉ�ã��䔨L��oZv:�D�P91͍��s
���S�K��C���I�%Ȇ����k�P��9k ����-��&�9r��D4�18� ('*��R& �?��Y�c{�a���$鏕�9��J�G�^\������(���)�6N����vt��y��0
���b"b6 L��p���iv���\P:w m���Ա5Q�X�Z�o}5֑H3f��hmy��)$	����j���|��a+�/��ĕX�E �m�6�����xK�#!4ǢTa��k/���4�U*أ����k1\��6'](C�a������F�EQnw"`>�Ƽ��1���?���i+u�=�١����/{�J���@ }��Z�=�ֲYpVGA�c�������''Ef����e��U���`B1��*섃шH�R7�ֆ6��P�[�U���%�y��5T�䊢`��Hs�����["�[$eJ*s� �*A���(�a}��$��z<F�r
FZec��� �;�o��P��U�b=�!I�u\��cX�n��EU3k�T��m�(e�Q�����h<�%��O��\�� ��c��i��0�!H�<�B8�I���}l�E�q�+��-�"b�XZWT�Ӫk���u+��%ƚ-��J�u+;yKsҲ!��p]����(4i�Z�xl��r)��4n�UY�	&-n������ڿ��p��c�-'-9- �_��X�j�c���ص��i����A	����+v�"Y�b�26g�����J+�΍�q�F�K`��`����X���^�8���mo�X��)��иprNL+pл�i|Kg�g��0��ib ��}ӧ���nF��Z����x��K��+��Ʉw��Xw��JM�Mb��"l���̑�d�h
y����W�T�r]��U3x�x}X=�DۨZ
���{���,��iR2�dsx2H9������pU����z+d�bP�w0ض����y�;;&����dF7��`�;\Հ��X�'ؐE��A�;ǲ�	����S]@�"�k L0B�9
����V��y��XjaLF�p�К�I�#�>�F���y����1�hq� �*�����1aI2P�N�+'���?�Vj�E�fȢ��=�A6M C���,'־}n��D9\V���p*�qR�:���}EdH��/TVEF�0��5X*|��]��
.�;!1L�ʜ��_�&oil_h�7Q!�Ʃr�O�0���,��}XG�2�����?�$)���(�}��p��}Y�
��^��y��O!���8o ��ʯ96FA+��p�#������ᒏT�N(eAMn} /o�ܴHD�	&�<qQii����x�K��e��;]4z�� #�=�+�9N#�1�a�r�!R����ÉOZ�ZgE��s��Ƀ߮�v��j���	����4d�ː������}�ؿ"��Fo?.�7e(J�ۣ�,Ƀ���NXcKa��`���D�W:�	͋��)�\���� �I��b0,!� ����e�4�^x�Fl8T���c/�
��(�� E�F�<2�y�8쏡T	�*3�h�F-@dJ��"y� �1��ϕt�6�`�$�`�,%,-���{�������{��U_	I��I�5�Q�E�[,h9ji&��I6#Q6iQ!!�8��vy�����u��b��yS��%Zk���k\!O	�:�	#�1�"J��j��ϩ��(�^�ʞ9�f�K`��pCm�sxLҵDb8xu�OjM.�T:k#b�M3�HUHE�_�GQ�8IH3�jN��p�di+Aa�Y�p��WJ�2"tZ!�Wml)�K�X<j��r��4����vΟ�;��`|f�1#��n�"0�1&�e�M��K�2q6K�����E�,n��n����|��=�"�\*�+(�$o�UƉTQ�Ɩ��?�F�- Ѵhk�WM�ɋC&5+t���7�=����d�\y`�
��Fړ۠$�18�B�|z�Vp��;��z�!�g�@FV�b�R��HQԚ�� �\��vQǾqK(����oظq��(��j2�/'�qx��ޗ��?��1#��O�&�K6�"��������g���f���'Ym�(uL��CO�� ������%	v�����PD">���D�we[b�øJ#�θ{�
*n�(1��Z_�@�Qhk��Yx���[��%wt���/���������� �I��D4�t�q�	�7	l�y��^�hH���c�ZIO��_�&-��f-�4�]����R�������q��O2�vQ)�pނ&7�xr&�A.r?���7&��/N���\��d� �	7�5��uNpk�����`|@��	�ցU��,��G�OdJ��v6+ȃޤp=��Ű��sZ���1�8�0C��Ҫ�����Z'�U$#g׌���̜R��R�eq�N���:������=2��?����͵�(81�?��Xc'��?�F�?�8��Z)�x|�$e�S�`dL�]��M�����;�ܠ��T�,��(Q:��9��cyg7���c�8�2�k0�ON�8k�
k�ݦ��&�~O�k�7wz��G��7_��l"��o��p�P��"�OoI9����(�,�D]Ч�نx��GݡG�����ʰ^f]c�Y(�0����Ź\�W�R�!��	ܢR&S�s�x���sv� Hx��9ֱf�����o{Y!\���on���nlD�����s�Yk ���-��2u��I1�iS!~�Բ�`��Q[7L�aRSFIz���K��ދ�;>IY�4�(��//�/;EO\�G-^�U�D:�pU�eo�r@8n��dU<&P].����k!�Jc󷶪B�!�cw/��f��)x7�V}tw/#*�pyq��[5K��q�w��B6*���^.�������E2��qMO[k ~�K�KЏÅ����Tg<�9�R�ӮX�oJ�I��y�A�A$|����yeo��BhLERf�P��ST�d���'J)�f��s�w66x2�%�p�n��7vr���n�;,�]hYnx�YM ����M�ڪV��{F�%=���E��q��cA��E�M�t��f�G߯:Y�w �]�ޞe�qZf��fB!�NM���Q��o�^ށ�uokc'��?�f�(0Ec}�s>��͘��-�!��c/T���F�y(�����$kllRHV�ɥQ��5n���x��{�H�9)T�L�e�}#w�E�9c�uN�vymc��Xd�WDotx�����R�1&i��t�
��{K*����ϳ�N�5 ��u� �����*(k\=�
c����}����E=�F����}4�8��Q1���$�T���'�-x����ac��O���؈J�~��1�wY����M��E[���*�*�\�ʄ���ܙ})^�&!7�.�ݾ���JptK7~I��nDi	2þ��j	��X>���K���U�*���X%f�y�@uZ5�d�7Y��c�(�@��~>'�al���
júh���%$�?���)�2�M!gGR�����/M;�(�D5��4<�e��O���n%Q��C/�������";
fb�I_�p�)1]�򅆅r�$f����q���r��`_��4����?7�S /f�f��)��%��O�I��G�f�vG��p���6��eG���������jǧ/p
���^���&b�{��I
g7
�����S�~�}<<4IҢ�L����M��`�+)�]�	��t�u��e���1ʣ�$�z����O�I��J�VoFʼd�.B�b�=tL��,▓w�w�]~{�7�!���æy���gt+�)Z���Y�$7\�/ F�Z�!QiP��Z lM�ǳv���[�#8�"�v�iG��i�w��0�o����� #�Fwx9��H=�f�Q��M��ډA��� ���?��W;��g%��X��^�j�4�^�������uZ4��g7����Z4;�Y��M�sO���&�*sJ/|�@\���?��@m��8�ts
��,Q�q�9xI�~���T�I��6V0a��$�6nΏ!BB̞�8�^0��+|�>ˎg�Ɩ��?�&����� g�xr�@�[V�X�t��G��G���w��c{̲��/�>�<jф�^�9��^�Q����?w�z��Vfm���4�&~�UZ&��9�]��������"�lǆ��i�� W�TA��*�5�fy�ƍ�I�� �	7ɂE�T�N�=x�}�bG�*�`B�
ۺ|�2�t*�N1�	U2�x�>|;V�\ؚ]�5O�m���=)�
�Вhdu�-�I0V���X���*M�x��a�X���a���|���ע븸�o���R���Y�'�J0~<Z���>" 2���[ t1���cR��+��y$W�,(���9�U�h�'6m=^>��fGp�1V-�.%�����a�f���}�fYU�<x���ǹH&m����/��/H�߱�����O�	)���UZ�\�9��
�����wW�gi:���le7@�P^��͘%V,�&Y�i��[pƌT2�v��M�k�BVL�Ċ/N{A
i�BW{{�X���a>kDh���_*����#$�nF)ga��v��qa��ڎ��{f�)���p��)�͡s"G,��$��l80�ذ$IX>���u��h8�i�r��?���-_�gui�'�u��ƃ_"k ~i��~Z��8���c���WW�<�F'i�f�����g�EіTkb��z
[ŭ�� ���ߐl��0�
�����Bc��ڲe|���7 �$� �	7��S�AT��΀|Ѱ�p�jB-K
���2v,���l���S��� /��_�g+&��n���me"&]�>#�;�c>�U�(E�Z�����)
 Dy�sl�4�T�I�Y&��p�F.���˓�Ȏ
/x��GxJh�$'�]Eք����o�g��R��0��Ӣ�.[<�=���6�-�(DÙ��d���*�e�*�'�<��^po�U��� 㠚��qb��[�Vi�,^��N����(y��ޛ� ��q�X�^�Z0���Wخ �Y=�{�F�X0���}%̪����U���X�[4	���ϓ�~Z��l�+n�@)}1x{:�v�)<S�a�Ež;F,�c���N
w��<x:�1��{oY�Kb�oۗ�<�k��
����Q��E#+��a��w��aj�vǃV�b+=2�f���p���L�~�a�����������X�'ܤx{��2	U:qM��P�|�����í(�|R�ѩ�^��VC����G�H��p�T��+i���x��D4jKc�7v��>��G�8�ad�D�%�q�Q�"�yz��em��(� ���z�w��<��H*g*?�B��������]�ػ��_b��/<e-��WY4���/D�$�e��z;16RM�2�9���|����
Xx��C��\X�+��R�a�NWG6�1�@X4��و�b&'�95 �l� ��2�-?�����a[W�|?WMڲ'ka[˗dE�꜐��j��W����z�)s����ǽL-�4lu�+P��M��e��O�Q�#+XUU�6tI���@!Q.��\���&d�S��ǻ8uy)��Ul��E�-"�FC9/a��LQ줋 ���a�p͑1�{債>�T���\�Ȉ�6w"����t����n��Ԏ�oȍ�IKm~6�Y��A`'~4fǔ�)<�rC��-����S�)f�-�5 ��B&�/
�Ȩ��ӻ��9�9Mj����g�$k;^Ӓo9jQ�/�Xs1I��c����崊Ŷ��JV���"� _�N��`��:Q�4��ll���%���:�ᇥ�Q�fɽ��Ib�;��te�S.�M����c�x!�&Y�k��^���V��ES7xQ/(4ԘOq[���l��/���Y�KbU�?�2]�n�_��c.<��e=y!����4�8�a����Љ��h�c���9��{a�8��I��׆�Kj�(t�G�tXÆj���
�W]�8&�1���s�axI�����?�&�����p��}��e1Dc��)�I��c��#�;~�Q�p�S�����F�*7C�y�y�
�ЩH^����$��$�EVp9�\���G�(ÐYq_^Y]�l/��Zm=Ac'��?�f'<�(��_n��G���Q�Q&�!2�dvc���4G.�R�&�[ܘ]T��!�fx�z]�w^�V��*��(f�;���X���{��x���j5�*l�Fl~uj�}�g�T���;�� ��)�b]|s]0�FR�<�	J�&��W��:B�ҟ,��+qzM��-���K�"]�*��P�ɪ��x�ȼDG�XN�x_ʦ�M!��X��j�{	5ۃ�&::�ԯ1,��b��uDC�&6m��vV�h���7c����,*i_�s���J���*Y��I����k�����:M;|��&��� �I��㉽MrBC4�(���j���ݨ d)L�NUFc"�v�n�H��~KZ�nBV:��[�e�;��2=�`r�,�/�����Q2E�h�جۣ&is�t1S�NL�f����*Ģq\{��G��Ф����֣bV|m�77vr��%0CMT�w����#�g *�&��4���Ӌ��0�E��r�r �T
�O� �
A���(p���0�<޽%�^kW����`���sb��{�a6vN��a�Tl���B�Y�z�\嬱�����,�`�Ԛ�=d��uV�X,c���s��}�B�N^�A�`�Lfg
~J����lA���ã��<xn���LT���
����~��J.�1��E�7\=vA\�{'	�1�4g;je�{{Y��n���W˸ ���샧tr�â�#6�����hd��]x?���˞���E �&���%u���˞��ͤ��!�Ҿ�E�]���㩅���G��38�9F�"o�|�Śwz	�	�2���Q5�����s��dMx�J�O}^�>��K�jձ1�i�)�k�'�t�F�-����MZ�-\���N�"k����6$�0��cє|9��(t4���Y�b���7��h���_b�k�vX~�"C&����y��'T��&,O;[�
�췔��y8h�t�S`TϢ��k�E���?�K�V�	���s���g�^Ǵ��8�;sK��l���M�Yv3y��()����X��y�1��+��!�0S٥K_\B�`��w�r��A$n���&��8�`˾��YFfYUg9�XI#T�Yc���q����m�����c�`���j2z��y������o��+��l=R��>��X?SJ@�rΟ]AGs_�c�`�+�E��n�,Ii��� �&Lg�G�đ�&�k�Hkgj,���@;U��qݏȃ�^hl��\"���E��&<^Q��:��v�̛ocW���)k ���H�  �Z:j���D���J�K�0ɊTI�5S�M7<��Y��	�R7��܁�0��#��#&(�s7������h�د����d�z��xF�'Y�IV>Z`������ܙp&�v�8�Q0}V^)���PLQh��J���6atG���s06Sl����?F�7v���e�"�&t}�]�T�I��d9�S�ג~��._~���3���<��Ǣ��Bv%� TUe����u����
��2o˾�Ի��16��
����S����I�YY�Zl�ӕ��d����y�.D#�ͲX�K`�-V�t���Q%+�ڊ(�<�˾Xy��ֆH�ݚ1���Ym�a��i��RA�:=����3����B/n�YmWc�V0�������v��m�'D���X���7y��|9Xn̨�Sc�c�7�0bL�W4x���1�@�de�y<xX`ĭN�Es�sJwV{G�[L��v�����A��j���]��A^b�����m�h�gÐ������ӔI3�h>˶أ8�#��4�޵�X�;c�9i�ПXw3�t�� ����>�*��H�?�
Q���Tc���<�r��Q�[�����������4�8M�Z5I?�t���$k_JޤJ�Ƒ_k ����H�bC" ���_�a��̑�Wݯo�8"ˤh���X�	�S�W�Y4����s�L_�>���w��cֵ�H R����m�p�δoI��7c���� |c>"�>׷�1�P)~�˩Z���Ld�ԝ��5�Q�&��U��p��>�`�0 b*Ի�X4�@�w>D,{���G�{���=��D�?;�de"o~i��%5W���W,��9&D]�>g$���4l���E3w<�EM���ix�"�^�:8�Y�J(i�E�'G�P�6�8J���fE�&ML�z��*`�o��q�|-�h�m�Z6�^����f+U+Ր�(:v	��%R`�&�7��Z4���Ȏ`C��2�G9�T��J򝂥 ���5�x��*ש��D#\����B4��bo{��22pKhN��@�3���!�$�b�UCu����4� |c>�Ƌe�-��#�:�撇EC6�����ǏS��[@/���Up��tjx��M;^[�V������f^9!� ��wMl�Z[��:<klI��%0���n�5�h���˹ oQ��4ʘ�E#�6g5<x8P�{�X4̶�4vR�r0i��|���@�ۄ`Sp�f5�"�d=��{���7Sj��01��|�m���+�8C�l���rX�'�Jdǉ;�r�\b$EkQ�G���-U��b�K�Q�$-f#�1V����a��h+���M�,d���&_�>��Lu��)w�Z}ӖʓM�uy��%5ˎ�3��'�H�)c�������Q΋��3��.̂�qc��z�w"D��ˬ���&Z��Zz���7�4� ���r∋�	~�d%6u��ܣ�/� >���~W�������͑h!�<6��H	��$�I�����jR�Nѷ�(���Ȗ	�&�<� �	���%��qJ�(U���˛��
��M�c��h.XF�S3/�c�;��GqI��$�}@6���B������-� }0��s�p_&k ~	�P�N'�::���+$�V	,���V幺ti+t^���"Ģ,���K�V���!A��/m�b��<��!���-w)Z�ڒ�Ω�K�V�s�m���4�X�K`��U�0F3��7�aj��H��J4#\�E���Ң��р�,�iWp��m^$g��lE]�\�L��%ʃ�ȹ��ab���@ei0|��\rT�;->�±R1�#ܛ��Q��N��z�V��9ϒ�/�n��s�	A���4]�����5<���O��� Yķ�yG?%
����5�$�c��&I�Y���?x�F�������b;��0��<� 7��,OD]\��Y�*W��V�Rw�E3=B(U�T�ƤlT�<��TV�ƈ�?�}�!�B�Y4�9�Mv��yD��&B�\� �	7��
T;���Lĭ2�ʳ\'��&�P�8}�L-�l��D���E���:4�e����my��+6f�B������d0�S��i�BL��-'��'緻�9v5�eI�4=Y���_��>����Z-�b�f�;�?a���ь�c�p��(�uv�1/ˬ����hX`�t1��g�xN(� :�q�6��Րƚg�͇9˕*�9���X��`���<�)S'�52��3v1j!�ڇ�c�X�R�a��m����:5n�Ft{�縦�6k�8�����"!�Y��\��B[������p2ċ7���U�<r1�8I80
�Pa���Ao�X���-�%�y����*c�Q�Yn��/T�-<��������3��*��p9��?4"j��">Ը#�#���&���Q��3E�[�X44x�WLD��ǆ��,q�4jܛ$�X�Kj��|q�`��Y����w�]���|@�x�^�p��V �<��@�4ِ{p8����u
�.��aS'�����z�d�2���[�<��Q�u?l�E������D^��H��{����d5y��h%�����[��U�όX-�d�C��+|wvkgGֳh�x�Ģa7�$x�F1�N����I�#�4����Mi��^�����d�q�dݧ0��}j���ϳ�N�5 ���3�{�Q��B�H.xe���z,iwDG-���6 8�s����o)�h�������+���pE���' �p<��ON6���E��;�d<�dь���Um���X�9��d}���s�=�;�� |c��m␳j�+<88���p����hd�^[�ʽ1x�x\'U��	����p0�xV�̤����#
#�)[M�
q~�vIuZ4��C��8}1xw?l�8��z�g`r}�G�'ݐ���_I�����J8�h��I;5�8M 8�ξq�㸭���&��R��	��ifJ��6���'CP�5���BgG�j�m�=oߙFYՊ���E�����fW�"n ~i����� �L����'J���|[D��yΞ~���>f�,���o�Gm��Y&�Nϻ6�ѢѰq`��&��Є&F�t��腿7uR΃�O���|A��>Fm
<{��R.lٛ�����[�Р���2a*�X"�͹���x�5�1iᤴ����ΦA|�Q4�[ѐ\0,8|�n���;��_�mN �:5�Z4�p�����X�K`~v���H��[E���Qk�f�ܲ0��_*6�K�j�p��1��qҍ���'�$��K�q>-d�p&2����?���R���3�8��cBڑ���[�S�ԤMԄh���o�l�ѳ!`��::!�ˢt#��1�i�9L,̌;�E]R���O��$�_����O�ގ�P�_A䲒�ԃ�ĉ_��`n�
���_��&��b�R0I��a����v},��&ɜv�g,���âYD�'5�<EI01&ﵪ�W�$qc_^��h�q;$�Y:�&�h��`""�˙���ߣ�3�a{�6�,���d���uw��`�\7��%��O��V��RLg)c�g
�F�"r©�GP�=tH���g�wC���I�YIϏE��/%6��ش�e��a��`s5�& �����Ӳ/33�	��c�_�U�Ou�r@��K����$�<�G?���8���t��җ����p��}s�7�H�,�5 ��m�$�Q|Wlr��3 3��w��n	����M�N�blq��eh������WZ����x��Q=xC�TC�XT4�q��?�l��n�����n��16 M�tar�}	V� M2Ҩ��{~��g�׮�����B'��~<��{B4�d�s�ʕ��vL�b\���'�=��c�G�0����&�m.�>�'z������ػ��o춬,���!9x�m�F�s+Y�g����E����ڢ�=~�C��,�ݍ	X���c�+8����b��oG��q�b�}461�e��O��q�e
���(�"_G'�V��!l�()mk�Ǡa&Y�qv��!v���V���rc��M�k
��l �z��d˅���4�f��M�Y�{�qG�wa��I�.�5 ��B&d�^j��hG����a	�:���?�9���9�s��޺\<��d�5e���{�ǜ3~��;ךa:����΋���<`y�������
���q�T�<� |c�m��&����ڧ�p䗧��̱HGK����L�Y�Q�P�~�4ݞ�������<�8V�CU���;F��K�1Ԣa��_�I�s��rX�Kj���zd!�2:��M��B��e��� L�'��i��38�`8��r�dt
�B�w<�l����,�eUc���אŅ�b���~'<xԾɔ��X2c�e<x�:7�x�o��[J���M~y��%0a=���/.U���1�5=�\b�S8 y^a[YS %ŋ�������Ֆ}��\'�T1-���#�\2R���עI|<x�c�3rq�
��C�ؔ2ݶ�}s��=fRDR���-�F���-5t_���'���$
����X�K`�Mh��MG�����D�b2�,�V ���"UPk��&_�?D3���15
��$�͡3ah��D�L�����Z4�*��w>��ػ��?�V��BY���o��\KX�,�N��%9Z$G�:]��{_5y�4�a����6*��<GW}���V�[ V^{�ă���-��~A�@*��ڷ@��B�h��a�F�
4�߁(Rc�^k �1��b�ĢqB
���,N#j��s�.o����#෗E��Sze�e<�G�ٱ��GMaUz!�Vר���_`����17QD���5���X��-n\�2DSJ�F�Z�� %�.-�Gd�Dq�N�jkmhc����=<x!��Y�{�z���w��հ���OT5����}+]�ؗ��o�k�e�`7���'�ob)�hB�������]�)�~Lt���xX�V{~���mp���?�̘ф�;*�âh�G�(<:V�˟�/}3Eɇ����ola�Y�^���D	!yw��>�hZ����:	���yTQbs`�� '���p�>욤}?h��\��z񸚐�*���9�q�kՎ���5��%���-#�5,�3��#%�/_vz��
���)��/2¶|IV
���)��ƅ��e0�xY4�K:O�ؔ��\�mą:~��Rb
Y4��:�#[�_,��.�ă�U�R�`�l(U0ۭ˱���e��������XfĦ��\�3�q>`L�X���{	 s�O�Sh�h��t���iKd�j!/_O<z����my�ƶ)F-,��<F�5'|�=eY����ȥ�޽ F"�1�c�Xu���)����4��墌�!�J�
<��g�#(����
W򻂏I�O�����X�K`�ݹ%9&X29�3W1�ؓ�ۙ���:����ۊw2�P�s�-���{�Yp���-QӅ��9<���&=xwel�s|r�=�
����2Ex�xg8��t��+���Z�$L5�����[��D~LvfO�ҥ�
�!��<(J�ʛ{�w�n>"��ɳ*�ڢ]��93�Dv��m�Q���D�2O'����~�ʑ�6��&~$G.�"ǂ���i۷<� ����aq�1/e��+�	��>W�+�G�)��U�h\�F�0@i�n3O�P\H���?<s������q��]iM��!^F<%�M����a�8��sT�����w蘜@Q��5�� �	7Y~�}_iL
����Y�I!k��eJ/��*Y�"�������-�����;����aê�;�U �?'��ԍ�
|qgS�7R�Vw/��	kB4G��d#.c�8����)���Ч��l�/�Ej��!U��+�{�rmu,��c���+L�&�%�U���?5K��4��H��TDU�b��&�!&��Xx�v��+�Ҫ<�h�~�c���� ���|�A�������f�J$� ��J�[~-�Z�σ�p{�Ig��e�c���E��b�>-L�Zl���eV�<x)��֓ZƎ��ܯ�]I� �z�ׄZfgGw��e���-C��s�O"��F����|<�����Uo�f�MP�������Z��mB���T<��v9��c�@�{$cBte���<x{��y�������M��ii���nR�����>����+����Ie��b����+8�Pe�'>zWAtַ".:R̞�SN��_��TJ�|��}e��Em������e^t��0L�F< )���)��Xw������r�{�8��3������'��/�#� �#��
�F��;�>��=b�o��Mq�Ɠ_k ���L��7��Q��8aA����$q�~la���h�FE���}�*���	6̌Q����4Ib�p+	I�xY4�f�:]CJ��a�:�$��S��	S6��d� ���|�,�-�6� ���)ɚ�����\g�e�o�Y��I���3�s��X4�������Mwޱ�G��cF��/%q܃=Y�.�P���� =�x;���U���c�ώ��x���`a�;{�%�{���%��Dj��D0͑������gElh� �:�re�S�h�'DS&E��Q{I.��	�&$�����(�+U��ĺ��������=bcX��*�-�%O��U�o��*#�ES�Ӡ�vaSk<�����Z��x]��6�����I�C����]�<��y���'k��Zp1
2���-���dѐF��/�X46T��4�5����)��k.�HcO�m��m8E���p�)%���ƍ'~	��Ƽ��5�z�QG��� D�'����Ƀ���~��Yvc�R(���N���5�ˠǊӃ���#h��>��f�����
�m��g�q��:�҃/�SM˾��O�U�|���<|���F����Q�����]��xi�`��ictl�i[r\��7�ÐP�ok9��;=��L$��'=��<�/�5 �-��.Eک�Ҩ��Q ��?賨ݲ���ixV� d����al��$V��t&�-����V9�ܦ><�h�'��~�����z�hʽ��rR9w�0!����+m�Ɩ��?�,���|������{�hȤI�*�
���F��Y�VU���os����6�h:Fq��H��Bf�q1M=[���㐎fEW�Wr��)�x,��� _iCqv�H����=Y97U�pM�r�;�����Cd�k�&"q�0�)�S��B/�B�Ɩ��ol!�j͖P%pRC�K��V�e��LOz��߆���D�>HƯ�L��#��D�J]n^�3�)iI�\�l\m�'�
�Ca�`渜t�1���N�T��^����T��x�-�(/P5>=~Aɦ�u٬�%1Si�4#i5c�nOR$�f�!�2��h�7:<�7��l�Ӣ��n�(>_2@��6!7�r�m�_c����<r�9s��>θ%:�߃�F*��V�79[y͍ɷ�*��������>3�J�Ɩ��_#L���)mk�{�T΅!v�~>-�������g��b�nCVg��qeՠu�Ç��Za�1xǢa�΢7]���H�wɢy��Ż7lÃ_>k ~)��{�3.S�ҩJ��>���j�%z�q�(��N��~R'A�,�BVK(_q��e���a�����s1��g�`n"nIo�j�:�$��hj ~٬������6b��:0��p	������lu?˂�4����6�1h^�mG	T��\Afc��/Z��b��G��3�a붳���$�ͲY�'�j3��� ?�4)� ��>��){�J��B4[�s�~>�1�����ɋ��{������x����j�L����»`�@�o�m4jD���y�����7m0�؉����!~���E��t-�Q]y�Ϣ��g!�iw#ɵ�fW�hdMX���*�-T��{���BH��2Ë[���ȃo/�g�\�2����/�5 ��J#�[N�A���PJ;�Eإ�P�u�.����i�r��Xý�ϗ�o+��b\_+���y�rZj��w�D0��s�ny�	�f0p:�{b�rK���*�ds�x�UŤ(��H���q��m���ӫg�Юw���C��;�G�֦�uI��n��#ĝ���}����+=���rb 7�Ï�!��Ł��>����M��~�A�c�\5��]�1x��p�% �$%�g���FX6Jx�WW�J8>�ECO�J֥��O��w+����M�X�A���[]�`t�3f6�@ޤ�Zi����
>J;<g[��?8�-���Q6��
y��طw��4@x���I����E#�,���i�ܰ�[�
�M��"��&��RX�'�п-c���+l{}f���w��afzRJ�du�fFZ�,,���:eR�t�Q�;����^iۜMP3��cyk6�*�n�:�"�LF�|T/(&��&Y�͎d5y��e\�^:�3��1� ��Y�K`�[2��*����swla�B%�m��O"p.ưLx�?�[p�=���׏(��Ϣa���(_��ҕ���mj�'��g/ݓ8��P�S�;�aH���1!ؙ3gF�X�'ܤ����̟p�o��b��_K�B�ݓ��J��I�1i6����[uAހv��k�Q�Of'�����|�����G�>��4K}��~=x���������#�<6�(�á�)$����c��/�5 �4��\��~���-X��<
7�E ��(�ɋG1�P�Ng���:0jw:���;Q�N�NM�}�<$�Ω�Vtz[��1&Yki�,��hx��c��T��{;�tU�3�*����n`Q�?"VW���G���g?����T���RY�K`�fΧ]����!�!�v܅0!1ձ~(g��qI�<l�d#��q�
��Ö}<�Ɍk,�a.C �{�N���0b¤�9�!G_�b_M+�p�_�e���O��g�J�H��`��
S�mkS��
oK	͸��*�J������F
��R��T<gF���sI�bݽ�n�K�0^����I��iգ�L4�v�4X3��z������E�,� �	7�����\�S[���� & �1̂��B��4���69ü�6�%-��]���Mne����J<[��& ����9P��R�[n/SDD)W�6o��p�u �ȦW�s�1\�fu�7�"ð���k�~I`i��
��&���؎��'-p� '�/����5��?M�FX��9]����ۆ�s��w���o,�u�%��.��]7��������
��e��b6([��"���;�b���ݟD��~Y�y�O�q�H�9Tv8����q=TT�D���:Ya.��'���r���#�Qä�HD���T�����V�ԚN����O|^u?�h�Y4�A�T���vx���%/O���EY�D|G���< ?g��(W�̭2���X�<�;B�_��$&m]� �����W��:���Ը8!>O��v�h��P���ul}�#Q���r��8N,2���bc�a��p����_l�N�h�����ϴ��`cʮC�q�����>�Aq1*�Č�������+��@�	��
�`d�I�����>C _A%��S�m-x.�X�3'����[��sO+5�?bǲ��� 9�k����$�㗬�/?G����%������޼�)l��+"8��p��ip_��8�F�,��q�w�Լ�b4�y�赛"L��d$��Z4����m"� ��A�$� �	�4���l�^��CY6�����<y��-��!��u�+���J�o�6S(Q����V�b��$��0X"�e�F8��/v���e� Ԏ�2:�		��j��~�JS -��\�>�r��7MQ���=U�-��u��� ��`����R�&�9K���ʇu/5'�6i�y�#�8�gK�fl5\�<x3��@qs�3��)<{�A{tNXt�+�� �Ա�9{wZ�'ܶw��ҶZ�ٟ����E}л�Mn X�^��Vk�����<��B�,a�:C!�$I0�`̞�`���4r��(8F��/\9׫�K|R����n�z��@>�l�\۵]u⍆��ʴ�c���:Q���
�r�Z��b8�VlE8��D��4�
@��6L4j��d�i�p*)�?6�}�c��sk���C%L
ث�"���j��,׷�� Ql,�$���.��f�ULE,뗂p�o���U6P�C��2W�^m��%��O��ij���2�ޞ���/������u��3Fڡ�Ќ�Bx���sR���f(rf&ǖC �1�`��A���_x����K����s���j�{}�
pv��+����%�:��&�2����*�Z-�:��0���r1t7$p�1�� ����W�iL��t$1c��i�+�8�C����� �,�H�&J��?1Ӑg���Q�@Y�� WEZX��a6��r�<3	2��e���SRƫ����q���A��'���5��X�'�vvvl��[��� ��~�(~SS��k�t�LN�2Y�2���1�߳C9ȳ46-�t��X_��@���۹<�7�5�p�����f������3����]%t����������`Kg��� ? �5R!]RP��&�Z��~���	ꡅ��N����-���*���۾�ӧ��n|	$1Ʉ$���d2#�H0<$� ��i�'�2�(�F�B	((`��0��2���`�1�;vb��۷���sٗ�V5���u���9��3���ڽ�����gkժU����̌?�_4�!�ycw�`��U9�NI,49&$��^���5i���E�����rZg�/���v.�W�z��.�Y��T�!VB*�)�"4H�m&$/^���Ҭ���S�[�n�o������O�)�x��y�����<Mj{�j�j۴��>t�V�J.�{���_�bt�˜h2��5K�i�X�L�i3F�n�t�k�J����CŅ־�}��S">�67��Ez��B�����s=Y�v�,���vJ��ȿUI�y.�&0S$ֈ5�-8zo}�SeԦD�<�n?z���$Idۮ�6Ѭ���	��5Ֆk�,^�B��^���:u�Wۼ�Ҹ8�I���X�FNs���^Ow�p�-��e#�ȮI�@XT�~W^��H��]'j��&���ٳ��	>`�?����btss��tk�n�I�,R��l�4>�	�e����k7�'�
��Ћ���dst��)b%��EJB���5i���|��O�:�c{{]Uu�y�l�dDԤZ�4-p\O�h{��v3|u�M�uߑ�l{e&s�k�tE�I.���|e�غ���rr׉�̇C��b���s6O��)F����/m���F9>u�L�x��3Y�c��>�D��X�k��z4ڐ7'[�c�j�M�Y/���'=5�*b��$�֕����]��sV���Q�M=f�Hĸn�T�B2���n?��Yڣ��4t�9�˳���]U
�=2�I��l.��"�����ɩS���33����dT���������~��iV�N^|��cJm�8}��UI2�j�Mg������[��r5���ܙ��ԧ�T���!�9��3OG�EO��+G���
�����'[�+�^����w6O�����X,����ʗ��'۪�o��ۚ�4�
�d��R��֥��˗������������͑#\<��߬ݷu�omO_=v��@��63ץ�ku��W�%����ħ~��JH�h���?�㢝^'�V�~d�K�)[�IB�6P*y�������7N���|JV�T6�%�_��Ym
R�/���zÜMŔ&�T^��+�$���M��cLܘ��_��~?�LUŮ�ujm�6Չ,++�|{�y�;�^m/\��I�7��b�(
�S{���O��a��������DW�h,�_����¥����?����4�++[�k_����P��5�S�H��x"Z<��ͭ�	�{>�_�X����?>O���CN���K'~��~��#�<2�ζ"�A$��@������n�?�=�)���[5=;ޞ�����?��ϕ'׆�p59����l�X���'D�U5����؞��������8�n�D��X�8��:��w���'�"�ۄgZ˕JT��ܤ��ͫ[���g.�SH�N�k���w��ʻ����ͦA`5�p�ܚ�ſ�ru�#�_y~�9�Y���}U.�v�����{�a�%y�`1��5�V���ի7'��[	��m��6�qlm���={�,e�#�<aB��9��#��:���^[���my{�*:�ioE�~O�����4�ɓ���#���+Wo��Ѥ~�hD��E�B3O���Jq׋�_�g�+�)	0��J�T����V����S����'�s�֩�����W������'�<O	"KE���_�DO���7�{o��omO���V����M�̉����7$��i�b;-+�A�����v5ښ4���ѱͭ�w�,�Oc��7_�"n\��|��_��_y����6"ч�H�����_>=��B���B+۳��zP��o�8�~��{���c�AoR�\׉r�S�Dz�7`��MT�2�j�Ɔ�s��L�e�h8"�#�^Wl�J��{˖�x�"��=��Ʉ����R}Y�x%�}w%�l0H�]���oV>蔈R������l�� m ��7����~V
&S��Jmqi����H��N0�ԈoN-D�(� ����D�O�B�'�ɒ�����Kح�������Q'��|c�,Ѯ�m�j�{��M��a�;!��Y+�K���n@�"qV�S��d�u�/���xɼ("��@�c�Sh{��'�P�i4z��uJ � <,��+L�s�r�j���3R"�H!D�L�����k �ޓ'O^�������7��駟~���"�G|/"|`�)?Y��~�ڽ��~�i�i;���,î��x�	��{�q���%�q"w�X ˮ,���J",�vt���go+����%G�p1�Um����Q����5�m��s)��i��" ����a�0�X���7��jSv�ô� �@J�;t��?<����L�4&,�>寚`+k.��6�@[�N�m�4T�7E�6`�4KZD8c��/u^.L��&���y�` w��L�iiz�RU���2��-γ���f�ia�Q���p��m�3�+$��H���|���.P��5��6+�#�e](�T�Q&U����!�������3g^`���C$���yksu:��K���L�:�Abu-MP1fB�N4טx&�"�Z#�e���K X�$y�kDt�C���ly�i�F�%�Ъ�ZY�CD�L����wK~�!fMc����C�(ȷڻ\k�`{*3�q.D"hɈ��Hf����4qGgH� ��/�E#M��yLba�P*�Vl�qMDw+f;v���NT^�zm\&�}Iڻ!�[�ji�?�J�����f�҂��]�g	�&\π��q�V��;؜���:�ݔ�I����׎;C���,�b�� 	>0�!�[�xY��<��Y2�;3�3.p�'H �֖I�n]8 aM�o��-bn���&"��+��͆<��\MF�	U��ZC�B�*�"[��2J���8T��lmh�y�C���YΒ�/��:�q�m$3s���o���Uض�<���-_��v�'��趤Z�����ˤ�1���҈�4������9P&��pJ��1�"-ߝm!��JuH<φ4[W��5�0=�q"h���L�D�S�qK��UU�]�7n܈^5"|`W㶬�!n�֨kء
�D��1+8Į��B�1��S^EbXV_�s-�5�(�I���%�mC���ڻ`VggD()�@��ā�3Ң]�a	31�Υr�lX!`k����������
�ś�����־�kM��������y7�J3��k�Ԛ���I�Շ���3�L[7�K����&�Hc�
�om�F�z62?%qo�Lƾ�j)�s3
��^�&�Q/ئ��YH}����s�Znꕕ�������^E$���Uݖ��s7tlF����:��:��_z;�U=ϣgVî�Կ��=�Wּ>m��Ě��*׎ֻ����u���i+i;��~�z}��������IU~���� ��7J���O�;�k����U���&m����Y��v�
}���\j5��],�g�َ�бy�F���������R����A�G�fx���="J����;��A8����n��0�䮛K�A	�7YY\���7�H�a"N�#�b�G��p	>0ؓ��6b)H���^BE$�0�������7 "�D �/q p`�W�e�M2@D���#��F�ި���H���~��ˈ��E�s�α��	>0��68�mЉ�X���B�J)��ׯGM����u�o���Mz�"|x�?ֈ�@��"�D$��`��>b)��Kbg}"|x��Q��88"�*"|`P&(z��G,|�E."�����<bYp㇍N,"HD��q(���,"HD�.T��X�7Ѷm\�	���C\d�XD�v?�Pa"|`�&�����G��H��!ƃ�8`�CĂM2LD�����@YMM4a"|`�q��"E$��M4� ��1.`D�q�SĲ�&R
$"�g����#�F����h����D��F,(�����C�8`���
�E$�0�3K���-��Cq ���#"���h�,���E$��m�o��E$�0���"*#|`��
"�x�v؈&"�G,�h�	�����G�戥@/�[�/�"|x�,�+�8�7�<(��>␈��F$����oD�^���M5��E,�� `D��DqHD?��	>0$I�ÿ�Eֈ���m�A#|`�m��F0�D���x&k��@�{	����w�F,���8"�,�څֈ�� �=z]�H��6xk�����>G$���X��"�BZ�B���">���X�X��ݰ� 	>0`�/����g��4��(��{6��;>�v�?/�v�g��mA�{���ui������r�}�{�X��t�w���E���,����n[�_�g��w�h��ōq#|` ��UR��~��a�$��A�g&l!�"}���u|�;���Ed��	���WW�2d���_s�[$@�i��|�ؽ��	i�B��tn,�g��]����=wͥ���W\���Cw��#�,�v�DUU.�RD��?w�}��|��~^��v�u�Y¢v �"�^?�+ӵ���%�.�v��k���������� ݙ�+����EY���&�p	>0 T�� ��9���&v�����ZD�y���<(����`�ԝ�� _�|���}�up����t��,u>��-+�P�כ��4H�0��_YYџ1ή��.��qZ�q-��ө����g�fK~>'����(�=W^h�]�Gd�|���v��={���ُ}2���ׯ�۷o�" ��o����ĉluuU�d��o����]ڬ�ٿ�r��>v��q������F���˳� ����>1�9sfFή>��ʕ+����eЗ�'O���@��������u�]w�>a\�c�r�|��_�p���y���w��[[[������}fhөS�عs�f�������͛3����dnA#"8D������s�����~���رc�H^{�5��㏳g�yf_m���A�(�C��&��K/��{�1M��������q����1��|@�, ����^��ĝYb���L�gV�����W��	�k��b�x�;���������o���k_�{��g���0���w�x@�cz����/|�mll,4����������(�������?�nݺ���	[7>��p�g?��=�y������|������i�=�hE$���(�ӂ��B˄��q��a췈
"�f�4w�}�l���s�-m�v )���-�	���Iז��A���>A�F��~�i}�O��i�)"/�:-z?�:�F@��ْ3�`����"�O�ȇrP�3e]�zuG�n�~ ��0����S��z]E>PD�]?xG���k��t��;�ue�e��Z�tvx���e�EF�q�A�L�v��uķ3�u8Rs$�T����N���{������#�En������W�^/~���7c�1�=�������&PD� O�����*��*�T�'�E.�NKt��w_S��G���E���^.^(��.1v}��"�>CӅ�u,ʷ���_��t��e��uc���g�� �i�垏~(�����ܸ:���{&H���W:3�a��H���k��58���%���/`�D�Q_8t��Z��Ev���x����Ϣ�D�]�?^�h�n@� PG�~��u��g:��^]�~�MZ�ӷ�����p�px�u��3��$�۷��d��	ܑ�������3M���N,Y�#/����e۴h�P�Ce���r%vWF�=���������8�J�b���	>0,�E���}B[NC�m�Ε� �q���};�����٭+8��i����/Z3���]���m����S�]�ݟit�:ݲ\:?��	�G��~�K:��+c/3B�Ⱥ���/*ן�U���e��i�NX��,��u�)�/�0B����ٙ|�����}��]y��^�����#|`��w�`�;m��ؗ���ҵ�d�u�s�pd�� 2���P�|��cQrY��&���j�6tw�v�2��c<0Yd^Y�޽���ǵS�>��{��"�B$�01��EU�m��	����N{t^3�,�{!��l\�]-����X��8�t�Q��;��xxA��D���y�76������Ej�������	tgNc|�8D~9v�a��~��"|`�?����������l��~�&��e�<��.M|v�rWS�K�tBă���ru��aO�Ʌ+peFP8�~�E�1^n�v���v�:������n�tQ?�������շW9]���`l�B��B#)�'��H����������꫚ �������讁h���'�d/���l!$�݈�P7v����o����d9���ȏ6��/��� ��v�".�a<XP� �}!�ߵk��Ȋ���׿��qAϰ�!��n\��Ǖ���SO�Pnf���ᢽn|P/�}��U<s�{����'[�d��`	>0t������Z!�l� ���,ҺQ����� �-������pD�� ��9�Mh�~̖E��i�O<���f�:p�,K�t�.]���q�������Dz(��8��������c���/�c��?;Y�=�tPg��2\�P�=L4q�S��8����j�- v}�A4 ��L�]���)��!݀`nwk��~��f�f�~�%p�����n_����5i�n9�2���!}�����g�q�x9��(D�ꁮ�ú�F|� |`�ƃw?z��X�����]s��`?���'�E�J�u�EξYĕ�%����տ�@Z]7EG��~��J��Q�����~=��&����P�2����d����H�ab��K~�����ny{aWkt׀.�uObګ�E��B��㰮����]�X��[��0~��l�w�]D��U	i4ф�H�����kjXd����ȯ{��$_�\�ȹ(f��ձ�M��.�D��^�����}�Op-�������y2��������TVE��0"�x��߻���t}�g?�"x����}B������o��ۏE��5����D{;���][]���͆�=���o���F�@	>0���{-�u5n]_��/w/�w�Y�^��~:_tw��eZ48���K��!�)ŏm�6^�UF���`/o_(�c��]B��7v,�N�l,PD���V���bY�!/��׽��܋�z/�w�����%�ED��澌�l��B�(�E.�{��M��3:�/��w|����b��	>0pW$n\�X�`�5�@��60(� �T#�L4��d���C$�������8v�&"@D��M2�h"�i�q�0"�k��~��"�hF$�� ��ud_D�>�,j��"|h0������m��]����m��v�ڳ!���S�ԾV!_�X��N
��H�v��}ʑ�ەu{���jϢrv�]���������~u�����u-�G�a���+�\u��,�"��H���g��I4�h�n��~� r�	Z��'��ɥ�ƙݼD�Z��2�)ĖE:N/�\��u����������)1/���%�u]�$�L�Xv3����jFLh�df��K���kf$�21u�v(��V�6L�,'��W�{ǔݜ��]�  eIDAT���[Ru�_���f��2-p�u�zC|�w��i_uSOjG�D.��7}��''����='�3Q�Ċ��'P����3kYM��e�&�i[�u4��H���i%EbB�*C�>�M����f�h���5I�&�!$����2_#m)E�ә�&���|W��y.!���U���ۤ7�p˯j^��͈�y�fAU�S�iEB'aM[�2��"�u}�o�8�պN%��6�Znڜ�����7�	 �\A�����*O0$���[25����n;�-1��t��`�g��8W��H5�%D�Y4��H����IJu������b���|����1��0���i}=�G%�S��Z�k��kۦc6������AH���C����М�m��h�A
ڿ���iX�D�-�;[��a��\�O�A�t��_�CJ}�N�q+��� j��p�u�z��e��s�(�����&uy�͍bN�9]ߌ��)�X�f<6 ��z)>�0�&�0	><*�Э-q~�s�&o����H��5�m�7�qb�P�WY������z�<7s"T�am@0��M���l��JA�k6g��>����m�+�Zs��͊�d��[[P���t#���l23^͚c�����u֚yR��YϔX��cq�Ml�n���c��H�5�O�v�8���e>8Q����m<����H������۲�9��!��[��=�� ��R���ϥ5D��W�����sk*!�ɵf.�&��S6�	�}fqz�i���3�N�������n'3C��!(����8�u���ފ1�4KV�t�(�|n���X�|��%�����n�c��[ImK�6d���sj��+���Ӓ�p-(Z�Ϭg���Or�Bϼ�zk'te������Kr��l��*���`sf5Kz�8h��ق�g��d�[��Z�����I�Yc�`J�J*D8eF����Ѽ��f�-xOY���$�SP+{�Q�pܕ��2ۖ�ڗ�g������1V�,)�ֈkm�a3���^>n�A�Zmzd�HQ3p�G-jڀ�6ổo3����1+�Mg��_��e��M5�3	n��j�̳���:j�7̴P�Q[&�S+�"��Ԕn۵U��'!t4ɸ�&"�!e �!Qș� �0�1D
)�C�?�)��նbo1Cb�cR�9�4�c���,�����Fm��}&zD�����MfM���@>�(��$#-Sh�&C�Ը��elגmX�Ar��չ�r)=W�YH�~Ia�vЧ�2�Y�%Hԁ���#��IN�i�0�h��A�TfE��Y��# ���	Aq�^'����ř�,���+�v���0�� ����Y����U�v��%4EJ��݈J3sC�ڔR�!����1+"(�}�m�k/�ޅuk�XHS=zM�G��B�Q�J�H������D�cCh��l<1&ALӓ&������n����P�I��Q"Ի���lۂ�Ը�Aod"��Ґ'vɰbVH��c��L�'�%"k�܅��S� BlK�,%ү���{y���!�5���i�N��]1��Q�	mN����������ֶ��d~8�!Ԝ���D�n�of��ꨨ��)��F��T�3����ՐҜ��OS�W�,���/��}�%��2�2�,������֧���	;�'��9�(��fUc$�;uaP�Mj�XZ���09F]8M߆�����U��`�5��J3\�-=30s6Y�D$���y+�`�;���*Y�ț5�U��]B�'�w�������+�@c�v掙�	���;S���]�m"_�&Ə�7j�z=%D�T3�l&D����3c'Śڑ�#�:Y���N�O6 �N��,��XՔ�u	5�v���D��2�)�k(Zs5�$�L�j�N��%CV�6!��Ͳq^���Bt&�#4'{D��O�-���[��� [Y]a#*oJrTn?m��ڣE�`Xi����,�fSj� a���$�G䜦=���H[ޤ�0�6vA��Zz.pG?Jm�k�cͤaeY��I�
Fݲ^�1Y���2�1�"J[�f&!��W1Ӣ1�@ٚTl��va�%	����l8`�T�F��x�$��&LD����E{���&�1�_�	�#zݷΈX�&9M��B�&DʔY��Ԛ,�k�	��7TLr��=s7��)b�!��
���#��Ŵe"/(]C�ݾ��'<Y��l�j�͊A���-�cV������C-w�gl�$,*�5��K�������4ߌtiٲ�����F�)�˩n�F��>�A�w_e,m[�!K���r�Y�v��o����xTxZ�
��Yգ��k!�Mmn�A�Qܖ�QR� A%e�=��h��q�ܓF�ڟ(N2M�Q�����+�Nglω4�q8d�8� R�Dl��y2�fG�ڕ�K���	�{���?�k`&�m�1�����{��P@ՙ�3jcA�������'���|�lKD�����v�z�8� ��C�P��5i\Bw�ٔzj��kں�����㸽��l)��+�n�M´�cf:��jM3�k�<%��(=F��3�x��7vl����yM?�j��&�9��9Z2�e�K��'^�uz�y�D�P_�;��F��H�!5��vGT�
�]��gi�:X�nb?x�ir����D#��ۙʬKcb��hW�jz�����4x�d3s���
�b��h����I���q~P{i��,�)�n�l`�h\��ڦ�Wf)�9#�#4���9tN��;V�ſ��)�|0˅\�V��^0n��E����Ռ�166S��w��;ԩ�l�F/-ЬIB��~�z��Ŗ�fC(��fMH�ç�(C�H����-�}nti�ݞ��&Kh��\�6s�yf4~�Ӯj�JrD�gߕ���<�u\�UӴ��4�7Te���j�����9%J�fm��qb&�X@��t�B�FӐ�mf;HM�=�ѥ��y�b����7��f��v�����,�W��n/��m���as�K��Ԍ�6�HS_�v�I����6,���s�9��?bnc�h��z��,e��]�<X�Q�y*�M4a"|pH5��R�pzll�˹�L:�;�K墕X����vo�Gi)�%`n��z�<m@Zܘ`���'�\]�n�Pp{�ٙ�i��^h�������W��S[w�A�|nRB�$�|��* �Lr����vh��2���yxC�3�v�Q�_ʍ��3��A[3�uc��Bgƻf��+h��{��7>���C�0G�z���##Ȕ��'$(S� �Z���\5�DJ��,�,"�s���ۃ2T��*�2t�
�bbꎐ"�WD��!$?�TkMz���7��ǣ�3'cY�j�V��~��&��m�f�$��
)����jR6�#�&b�_�vg,��G,�vq!��V�e�����������)<]�e�f.D���HI��ƣ��k�����iA���4ɷ�9Wr6��(�~�n�Q�\�r�B�L��8�]G�da�X�Qh��4����i�Uh~JO����LI��C\� cLKU�q�ٙ�)�p'�zתf0��Ie=��;���"|hH���������fـ�ʆ�Z]�)��e%1餗�r:���ηڸI��J�3�Y�huX�<�Y?��O�8�.|�+���DL�1��t�K���HS��
�S��[f��f�dQ�����+I��ҳZ+6?�:T��?�'K�~����0!��H M���bŋ�Ҥ��u�y���6�{4&���2jKcB�Q%5�1�LXY���ŀZ��&,oM��E�
Ҏ�<Ӓ.�� m�l��O#m_t���>W���4��,8���ya;�z�L{ؤ������F�M|!,\K��Z��-[އ�ɍ{�6���L�[�l2ݦ���C R�T�@l`H�hr�5�ת"��H��#J�\�G,��JaA�f�ͲfoїZ���R�\k��H.E�F���^5�O�_dl:�AFک0:<����)CդZ;ϕq{�N��9v�h���T�L%*%M<I�&u�����٭�b��#"q�E�z���|���L���b+GzZ���3 �Z�l����S�Z�C�����?�+�q�T�03�$L�9�H�-``iI$�&����$xbf��oP�WI�*��+�I�6�:b��TDܷ[ID��s�;E}�g#'̈́Z���c[� �B���g��4^ �����++����ɨ�F6z�#�Ba����[���4�'IO�o��,M�|��F��Ѝ�m�=�F�zSUS7���jJ("���T�,ˮ���U���++�ZU�j{ďYe���b��d��m��/�^���\*�+[�Z�%�/Jk���V��r��W� ���O3�CFIyI�DZ/�<H��s'I��p��&혴�4m�O�
i��ք=��J �d�`3)+>	OV��R]3ٴIB��:ѱY IR�6�|E"�^�$�j �2M��;&��{V��4�HDGnq���3��72>MR��J���[#6XY%�� q>.k!z���Ƽ�Ī��^%44�I�H�#z���T��V�SVS��OD��&�)��+2�֭5��p/�m/I���W�J���"�	V*�⩂],��*�:�>r�S�:��p�Ңh��V�_�f2�j���
u{4�g�㘙HH=J�pH3����'��T�ʪH��IW�oUU�q��q�"�C$��@Z��b��D_O�V+�E�χ�C>�LX��q"N����h$��E��"#"��CG��bY�<KSQ��vc_���t�֎eS٨�Q�Q��#�?"����Fu!�<ႄC#R�rlH:���!S9Y�`2�������)�S9��ԁ�l�$�3ci�y��$#�N�<�XtMYEmD�)	��A)��k�|Mm��,���9b)%FD���>��aX������}�_Uc��D�D�$��Z�ȩ��_e-9i��ԩ�|�E��Pr�#w\1���j�D�ȔO����l��n���`��U�^Fϧ�� ��&B�eL�������b��O*5����������Ӫl�� �(]��b �r|��ֆ�M��x'�o�, mii��G�*AS4�e����$�^x��k"��_��_�z�ڵ������{��������D�xǽ/�t2���kkkk���q�?��'���G���}?��#G�K_��ذ�&TV��
ޫ���l����_ۘ.���"d_ۓ?��?m˘�>��G�{��8����?��o{�G�H�!����GIX��.7���N�������>�g���:�I��W��Ǟ�f\fk�5�.g�9٘��?��̵c;��.����sϱ�._��#g�q�	��U$YӰ|�_��g�4[0�b/?w�=G����?Ώ��Y�F���_g�_xa�q�~�c��YU��{��c�X�"�C$�����C�f�?p޼=q��w��'>�Y6v]�3�w	���g{��엿|`���3����H����~oe2��?����坔����󗏭W��C=t�N4>B)i�C������ߞp�߶�ʢY�*�Pj�|G�eݾ}{哟���C���,~�~kH�Z���?��O|b�� Ԯ�������{n[�v��c%����C��Z{��(~��~���_����{���/�_�"}�GN>����S�M��������-��<�K��K?%�|��}�?0��wh@�����US>��zWy�o����}b��?�ó�|��'���_��������?K9���p�����ɟ�ɿ�q�ֱ���O�o�z���7�>������GD�����y�Q��*���ī���{��>�H�o�������[wBV`F��*K�5!��;(���}�;�d�`�����w�)�Z�a����es�؅;�n�~�wVW}�Q���v�ś�nݸ�����_�jz'3j�<����/|鎶�~�_������K�~���w���g��o��o�mA�O�c9D��=    IEND�B`�PK
     o_�[Q��0�U  �U  /   images/a88da2ca-7e0d-495e-a5bf-cdc1eeca5e78.png�PNG

   IHDR   d   �   �M�m   	pHYs  �  ��+  U�IDATx��}�eE��{�ݯ�LObf`��$ad.�	Y]XWQ\1�((k��]WWpwq]�]&�5�E�I��Ȑa�c�t��U�שp���h�k����u�Su�9�j/>���k�v���xZ�N~���� �:xQJ]e(tuH ��0ٌ`�e�o�* xJ����^(W
 8�HH��"�h�B#��(-�O
�R}��Υ��_�x�/PW0����Z�6j��3��D� ���zܜp�H ��2��h&c ������Q�ejL1�Z!��� ��t�>gh�rY�Ѽ/~�D�� ��R*����{Ċ�+��� ~~�Mp����_��𶷞}��𠹽{w���������Р0�4pp��Ȍg��p�PdA���6�g��]4��!�I�;d������ 2���k�lڣd��i����j	������������{�����a�Z��o���ǏC�@���������oh�(��d��Sh�h�lG�����;�����o��}"�'�'`�-�Y�f͛�����_�^���ܓ���'��`x��BF��d�`��4S{*��.��9��/g����ߝI���T��c�e���󩧞z�Z1×~��n��g�dooߟ!�tK��X�c�U�һ(�!�(�h�8I�.IM�-�ӴAs=�$!��tJ1�e�H|f����C;�����'���|F�{,��L|���!�y��c�]oT�<��ɩUk׮=��h^����֭[��o;�Vɽ��y�s��y��ŋ�{��ժ#�A�SOb�`�N(�J�qb_���w�"�:�/eNc��/u�f��� f�� %y ΄��=�K��$9���Svh�=J(0�Nu��@����wl�r��ŋr)�Q�7� ^Vp��R�2�����3��n��!��t~^�W>���I�Vԁ��۷'�w�ɤ�ǵZ�Ҟ�������+d,�p�A`�]b����cǎ*���><�9�4���!�6#¤��8�{)K�ST�Z���dOOLL��C�{������緶o�~t":�+���I�U~�P�9���Wp��뵝s8�I M��v��;<�&�~	��%�H�#�$��1e[��v�8���<D���WRoo�Z!�z{N��H�"��sS���'I��Sk)k�?1\ĭ�'��
���J�c��5��S���%�Iw�E0�T�˜�,bD�3-/#��1/�is����b�ۣ�Uˉ$<_� �!\"bu�>�鬗����f��G=�Ԍۧ>c����WN���9
����#V��R���דkx�Oպ��*H�Z|�S����.�Ӫ 	-�e��D/��H�[��UO��N�*ޞi���2u��F4 ��Tߊ�s�s߷�r�8e��{(c�FH��5=�P�����'���z�
�����rd�]��^Yt�W����R��	�4z*4+��P�!$#G�,QHU'� �g*c��}ߚ;t���+[�9���R�]��9��*�#	MM������9F�Y�֪�����mk�&Ec.��؝o]4��#�ꩡF@��IVآ� C��nDB�	`�:z�����8Ozjʴ2K*��=����@��'D�,��t����q�}���/���-K�D2�Z�4+!�t�j\G��W����kj�#��;������|��j�I��H)*��0�>�K&��45���^�s>|�׆6?�A`d��o����/R��P��Yˎ�p=�����c�V�k7}�E�~��K� ��8���79�a2:>OM	!|!I���9%����ܼ�п%}~�?�s�ҏ��mG�\���S�+DiPFv�Yڔ�t�7�Z��4֌�q�N��38(c���	ɽ��������{�B�꟎���0%z�!!�����߲�L�3�8�T��p'�O<��j�0uC���<�]ҁ �����;�E�ViJ�+=�/�Z�d��GhP+��q4��������я���+�pTA!�8�Q0񯧧���dk�w�<k�s�	�@:ŤC�����쓤\�%*̚���O$�Mn�]	��V�bɧ��+��>Q�R$M?^@L��!)@�O�N\��Y
��|����~�O�C�����K;V�7�埛e��f���5��V�|�-�á���HQy5� ���a���N��d]�kh�
�kI%D�!IEmW]���^�פ��ܿ�W���2j�Q���~�85�@�(�[�z;L�?�<D�	����
�Z�
YD��n�z�m�ȌEX��f%6j7&+�9�@��}���W�Q�SQ�$AV5���ñ��3ڧ�xw���.���|,�Ο�j|�#�rY.ʥ�vM��"��B��^h��d������?	�I^�J=���$I��B�/_]��q|���f���y <A���b1��hY;}q�%��D ��ET@/�:����W?���\r�d$�pM*� W�q3%\�MTB�z ����a��]͸�y^����Q-_I��D�;i�)�#I��/%���pu�D`��n�#�N�%�c�F�|���7� ����()]�MjO���<x�e�\�㯭�RD� I��c�Qb8f��j��Y!�%c|KN�6:Lpd^%�p���-=>���\q�{�pҮ]'#��~)��F"�F��J��yγ�'^61U�� �����kg���`��� ϝh�S87d��MO��Z����&g;�����d�HtA�~�
��A���jx�y���f�AH>f���[�Ly�&�ZVJ&s�e5�Q5T4����b,f�79m����"��cpz��K��$��P�DK�ӂ�.\uo�
������3г3 -�i�x�=m�!�]L6�|x�D��=\�XUk�$�V�Lt+�SH�&�3�X�<h�/�q�s�KgK���|*>��-��u�eN�r�9��y�ppʝ�sH�4��5k���+�%�Q�L�L�n5����>�@�v���y�D�5�/$�bzo����R���*�S�s^A<������s�G��3)�qe1�����#���uu L�7W,����}_���ht�����޷AI��јvmn��1�U����դ����`�lRdLZ|�c�5�v)i�N#$6��p-I�#"H�=C]��E����A�	���r!����
�7 ��.+�i-���<��B���(�ӒS�!��H���&�ȼ���O���{K�љ�K��J���&<�E���߽픓[>>��"�v�����~��aӑ�eH�x����-�J�%��j��@<�,�Κ�r����B���
��Q�G�#�����Vr�:*�<�y���R������	����0/���2v&<������mDj���%5y�Wb��ⷔ� �'Ε,�l�3^�!��5��G���W��Kʁ=�<o��׳��w��1��,טA��P!D�,�9ʤY��D��gpߝ B�Ժ��L�21�1F�<�d1�E^�;,��e'/����w.����C���c!��T�H!�i�6)R���R�@R#�(�������5�"/TZ��b���u�u=���Ln��A�[��~CV��Wv����Z�Dz�r���+)�����v�#B�V����j����H5E"j�Weqj=���s��=�)�?R$.$Q��y2�d׀!��f�d� ]?9�;�#>6"�x��2U��Z�<'/���0j��Р͐��[Ԏ���������Iy
x�����c���Zp�b���$#X��]�)J����Gz��4r�3X-*�[^'*l'�a�r(s0��.<V(�5Az�sڊ�zj�K��P��v8s�1w�����h����[����I\�F"��P�q9�\cW@�G��Z�aK�3�Kӑ!+E1���zV�t�F����D�������vRB%�@�~�W���U���J��Bc�Bþ��|.��H�1/G���ዹ��z�gM���R���(�!���C�9f���6��'D�--$(�X��Z�����]�~w�#%Q@��X|������^'qr�*ђ_G�$H�$�;*�a�p&���o® a�T�-1�� ;;6by�̬:�_Y{��T�8�
���V=���bD�>�ݯ�����ሁ��+H�Uhf
���:�-e��<��AU��J�L�Y�8�w2�ƟBZ:>V������ݔ'�/#F��6�M�&&��F�cj!�����g1+iIp~ə�XR�!~�D�יD+v3��^����M;s�I7��(G![!m:q�9��@	9e4
3�wO�������Q1!)�ܔ0t:#���E�j�1o�O6P&2�#br�������4H�pf��KE�Q$%�l�9���0�b?i����y�eO�IfPv�YR�Oajr���b����1����`?k�AMt�!,��w�ϐ���q�GލRh�Ɔw�E�h�P���//�8�x$=����l��_�O��\�iXEAL��9� Kg1L�t��_t��p"~���XR����'b)O��s�=z����#�؍g���X�|�qT�Q�SG�_\�RQt�� �@3+�7��_�}�ލ}�����[���+�.(�V�~������T�	��;��� �?��<��������R"A�/�:��d��T�%y����]O!ĭ1H�h@P3p䫛�_�y�ّ }�:N��[)��#}�M�gCV9�}��>r�O飣���ȋ��,�ڦd�Uup��՝��/�n�:�1�D&/4�c�����>�"!�����}�ek��%ړ�QA�! A8:a���	���T�~uUC����}h5�Д[TD�����Ȋ��#��W$/q<d(�R��-�N�J�<�5$	y�H)rv4��#vqd�������:/�%j]�i�qZKgN�nR!���u$` A��Y��}$�,Qb�`�yY�zR����tҞ�zY{���gM��i#JlYZ�˨�YC,��9�	HU���QBJ]��R0�T�����&��� i���q	)j�Oq�>�9�M�N(I��ޕ;MM�"}v�9�h�&��b�J��׭m �Q�tH�2��S*u�GXA��L�$�p!$�(�3�U۱����{�1�E� acb����G.	��
��/�B�O�
HbiɁI�O�G�3x��ƍɕ j�J� B��e�݊B6�#��� �K�C�X���\�&�g���SY-���2o2V�.6A)XI��Iɴu!+�0zE(I��.�+�~�ժ�x)ZBi��K���Y�ۿ��~��}B���"OK���
�:)���B4���o<�3�8��V8�z��������r�+�YG��;��y��c�>Z�r�o��j�:v�:�9�%�v䛿WT��X3��lY�ax:���f�%�3������nmM��������-Z��ܬ�y��"q w��X��X݌Q�F���wOL~���&���k�)R�¡�9RH4s�4�
�����=Uy�1v��mr.�?��~I�30�Α�=GS��u֋�T��6|��M''�����X|�Ww���5m�/~���]RR����Lt�{�,w��!;tK��t�>���/���x�̓�Zt��7��I���Vtx�P%ǒrg�Gh�p���x�ݣ�{�X,����<�,SW�6.�ł��@��R��g�*q���$$�mE�D}�R��0�W�0=ݷ݉2�ܷX�#+`Tk�8�~7�,� S���i�����AY�����qp�^+v�1.O��F�����G�'P;R�\>Le��e��N�p�rHÀ������-9�E�t�7v�\�p'�i�"�^�qR:J�]yi�sn3�c��\��Z��'x�y��bZ���dF��l'����#ʠ+ d�^�Ra?�٦�k�n���	o�xJ�����_F�E��e�L)��`,!��$��(��ʄ�����2�h��Sc�b�5'��є1˔�v-i�-M\�&�Lԕ��U��@��`���lDI**���JR*UX�|L�:ӈ�C%��7���S�l������#���OD��:ΊX�]��Gq&�m�U�B0BD��,�(]�ig[�ǈ���e�A�d��f2�&''1��_��ځR�Z��$N��N����8b����?�
pu{86�a�V<�
8Fn1f:4�Ix�	��>8VVS��i�������V7pz���N�1�6E�"�����敚��@N��н����۴+a� �>!����sU��g�{0>y�t����w��{i�v�l��-�(��,%�u�\�d�A1"�a,�1��5�!��
����c�T��a�zd~��4b�c?��%�=2:��z��
�ظ"CF��Y��$y�i����
^�iy�ą�&��ϸ(�L�>�$�	 m+Y�#R�l22�W^�A!Ꙥ=|R�V��z�T4���>rya��U�1<+�a�����t~H�����s�H� ��}C�X���w��z����'�K��?YVf~%vc# ���f��1 M��
L�N�3ZT@f��}�dɫ'~�ej���s8;rr��OANF�wa8y�T7�v#+�~4�*A�������C��r�H��Lmf�3�0�Dd٨��8��;沇p`�Y��!e���&_����O��"�G��ekf�g�g�^��������^i�R��{�F9{MM�����,�2�9�2H.�Jp�*���c�N��}q^8���k��{"��3�y��T�Vo�Xެ#<Tz~�#~��?LYs_��?���!��Ӂ��|�<Dm~�d�.�4z2Q��y����	���%�"��#!��^X�.��q����(�1�22NxF��f+D���s�}Z��k��7�G���ly4�t�J*A��}�u�.&�U�c�V��cC���L�_�ߵb�{�09}>'��r�,�B��)F~���~V�9���Ko��2ڀZ�U�52j�;��d8Vxw/�W�p�M*�Ǔkߵ�v�Ow���+����m�j���/�2L.SZ��}hjXuv�MU�pVǌC����2�uA��Q�����{�ފW�(e�����}�_�Q�J���UON���7,f���]V��(n�K�C��fы�Ǉ���s��3����W@��בFT�U:���kA���\�~S�dȢ$�׊�#>�@��M����"�]=��|��}g�!��i:g�@�j�I�AO�E��� ��#�Q,�,iG�����!�Ɖ���گ��޸v\��h
����pd,,�K����e�r�v�#6�� e���%��E�D���j�I�#��-7m�A��O��p:��/�cLK�N�ӡ�_eH�={<*������#�);-i%��%;��a�:Oճ�_����c�s����H�|�3���d !(�?�yT�w��qS
�թ�9/��x˝�E��������NJ�z.���0���WH)��?���΋=����?X|�b��w�� �4!��307L=�a�d��4�rc�����C���0��K�6������ˣ5u�"��允
��\��!��3�7�4w�Ԅ�1��Qha" Q+�J,�[y�p�s���$�����,dTX�BvZ8&\�`#1��*���sz�~�����P�k�e^�>W��F�Iҁ��3����؏��I/�c��@D3�NNqu� ���	�I�N�?�����ޖ�׌�5��҈�+AM�$d:�:G2m�~���.������Ԥ?���\$+&A��zS61<�#sQ.�q���	Y�֩iM�S�����M�6�-��j�y��ҷ��&�i�ѹ�:���1]q׶�ѹ��B�)�4�mF�"�%���I�� cQkoH���	�i��>y�&P�&�H�0@�dIy�)	|�!!$�F*�NN������")�<��SJ**8�O)�0li�I����̐�Ț�:֢&���U��a���-lt���"n�R� &us�k�������t��z���F>�o�XN1#\h��=�x�^:ި�y,2.;p��<����y2.�s6�a����n���K�7R$< �i����J� �V�L��NF�(�0Je���'׏���Î�������5��	͆ޙ�(��%&M=�e��ap�����x��\�$^����'�ݯ[�.,]a�����"����KA,�����x���,l���m������ώ ��]�I�fF8Z�F��
=��fW���	�R3a:&k$�!��љ�:��'���ӔL�{�O�JN�4�LW���c�-��9dy�oP�i���
Q�#M����o����^e<&!�I'.Ca}��'�pt����}Ǎ��+e�x�>.�u�~�C��t{o�������{aj'�<a�U]vbȝ�UO�m|�k|���@T�P�]���{��� C4�2.z3�t4�Ĵ^�V��q6>Q`��tJ��{QD-����ܪSw���p����h�L�Fx@���������&��on��kl嘹C�l���['.SZ�v��f�!���c�)
S]�F����t����_���?
�a}�i�u����Y�e��������?�ڛY�8�����EFV4�-�O�ʎ�@>������	;��[PY��(���ڥEq���"���߅$WO��B�|u7�˰*Qx؎*�!2�i�dhAkPC���s��lL�Wq�0��Sc@���U~��B�%��P��3I�L���5������'Fw�����uˀ�U=6�ڽ-�diVj1ȸ]��B�.%�U��:d��m!R�:4��_p�)�]rʅq��M���܆&�2�sX_�2ֈdq#�xӿtU��}�$���W}nū>���J�0���|+ۀ�4=��s�{���=���(޴W���oX����T�Y�	K�]�ƕ�2ӌ�F�u1s��}Z���������B�5�����Y���É(G",B+��lƓt(�Q8Lh��_�9|�P,O�Ĥ�gU�B4�JT+�D&��7p݂�]2R/�����iB�;,��BR�D�5T�{��_���/]zm8�:�w�s�s[��^�r}I��E����hr��+4
��}��Z{���Į��d��G���?+��J*�����W�b`ڋ�H���$8����z��x�s9��s�!#�1�u�As*j:�D�7=K3���Jq�[y��>�a��X�(�C�d���j�8u0��INs�̟Q� D���1�n 3�&�{1Op�UVv��>><5�����jF|�MD�C��D	_�啾Cn�ؽ�:��x�h,��r��:q�cnz��#N��BΑ�Q��61�X�C�0Ъ3_J��T�E�7������j�e�$3W��0�d�ZOfR�86A�f�D{1�VQՀ��'!��b��rRTP+��ޥ�hI,�0z(��Ek?�,bt�����A+��ԲҰC*43l�3�+q5~b��і��� �v�uI��=�U$�EmtFX�FPV�QJ+���@� im�ŸML���K�(P�s�N+�j�'��LM�M�;1%9:�j3����z-�ɨ�k��B�M)�i)%�U�4@�Փ&5+��y+@�UE1���i@(u�Yc��|rL�T�mL����0j�Q�ʌ����	�ʼ��+#t���HcxD��8i24�}��Om:�4�	��B���)��~hBmIY�� �d2�,���N�M�C�m������M)�r;��xsOQ~*�·�$I���ޮ���Tذ�R�%։O   ��ŵ�
ѕ�]�f�_R�����/���b���V�O���xKA��xb/���qk,
�8xmD?N�v3P���i����@@\(N��.��dAF#C'���HM�H��I�i�Z��q�d�, [�.����4:� �������[ԋ��0���M[�M�32	�A��K�cq���j7��Tl\wh_�j�5����G��c��<ݻ��Y���<�o=�o�EC���.�ڹ$�n�D��c K>����5�)��퓪������D4o��j��~���*!m��Y{lS��7���"��M�n[%���-�W�yZy�YX����g�##U�\g.����$�TËa�����9}��N����*�ݓd�)�`��k�%:C�7h�!$��@$�����swu���C�r����&�X�ث;AOGȧ0l[�%
Q_�Wٝ�޼�v%]���YII��47�K+&.�=7yOk�jz.X�2Ŕ�P9yh!���V�3�D����:�NW�0u�J��f��������\�J�'����1E�`Ж#�v
�v�a�f
 �A;�o&%aO3�b��h��&^�(��@�<��e�T�M��z'x]/����֡7Ӑ���e���mo"Cq	�l��z��P2S�A+U���\��h|#�L�Y��ѾJ2���/�٭Q߂H���h���e�w6�]��K~K��dZ���y�gR��<��-ab
N��}~~�uD�kl}ּ�'��l*�Νؖg�Xئ,p]�Џd_e�o�Z�9x[[�Ҷ�ڢNP�����I8�N�Nl�)j��Sl���fp�!%9�w��\��̣����@�.0�d�Z8�ё��L~��^xKc�Sgr�w�$�]�����շ�a�E�1�x�s'>>^�W��:F�#���r$����Νa��X���x�v@f���mg�?m:�i&�C��*���Z�X=�@D����rc�/F�g���d��u9)N��Z�m�j2,W�5`����qϽå���/�YxnWq�g�� ��l6$�u��G�"Y,�J/ =� �]mҏ�n��7�/�N6��u�����+Z�i_!��E��w���`������،S�IG���J&�&�t�;��2�ξ7���d ��F�pbD��v���qN{��q	�Y�S�H�W)B{-?i)|�mʥs��/(���9T���c�z�jY��:'�73_L;	5��~#�4ii����pN��Z�����:�#�%��.4�)]�02���a/xuk�q!���B�~�����)͚N�5U�RX��/I�fm[wdE�X�~s9jR3g�7P��T)��{cv��]��Z�K�1��("�&�Ńȴќ����� �mU?��fT�zhG�UA���iMRj*���pB��Q�	�ޭˋ�V��J��?Y+��6
�WBQ��H�m�$�H�!�n`�d��ʽ���{��/��ojj����K��^JE<=.+8O7$K]���5�AT�xB�eR@%T�&�R��'CM.�F��(��N�Ihh��$�������+��Y
905��kQ0���I�����Lmk�����#�S��iK�T��m 1��%I���c��.���Z�o09q���xl\<ܔ�rz��L���<JKY���;��0�K7�u1a�6��Z8'Lն:务]�/���,	Vt/�0'It;"��7���I��,��$�E����S�	j�v&Ձ��\O����ܵ�FɵԙI��񭨯M�(�*}�S��S���m����DY�ɟX�fҢ�yӉ.��.z͕nA�j��(�OR�[ ��'����ø�S81׌(4稉�7:R�-�tB�7�|�W�g��� ��Ք"R����&��T*e�[� ��2�l07�\?�KǉI>�ŊyВ%����_]���hhӶ�v4�>��$i|	�3Q��Y=45�@��Ў=�p�(ǆ�wJ�]�����fB:�;R�Dv�������S��Q���?OG]�q��#�)z��fh��Y�����"���Iw6m�ޯ��R���*���	� �����H��Yҗ�#���)�ʮ�qu����\,��Zhj�5��eVoN]�~�5.)+�ml�b.P�����,c7qY,��*�	''^���N��e���"F���~�
�LW��O���ܲ�f/����I�/��{n���V�y��z�'��ٓ�=�̏^앺��c�����'�Z�,��Tt�1m��Utb��q���W��߯�Z��oB����t��Y w*���M����=���wnz�������ջjǞ?���a�uk�F*1'�S��`�A��& '�"�����-���p�k�F��o���� ���8�3Z����|���}���ho�K�8��toF��R�8��"]V,g͑m�����sS!ъvmS9�x���f4q{��2�d^��w�����S�J����c��iy^��/��Rkt��@��|u��B'm����%�[9�{����YfS0��s��!��R�$�ri�9{��k������������D�>s�S�9�C#n_( �O��*3uI�=��'e�O��0;@I��,���E:�>c#N �Zsjƴ۴b��4	?����Om�5���-����&,4u]�P$�?و��|f�uϓV����F�2c�֫�N�$�<�'��A�Q%:��H��TJ��3? �X���]%��rDK	JD�l>Z.4���B+�Eƛ��9Y�2n9+=���w�+#�N,�G-o���bXR_L��1�L6���A8�R�jԂo��;�G'Պ4%�I�鲹�����V�a�ੈ�֊Jk�����%�A�U��&��n��;6C�e3s'����
��rF&N�Hc��C^�뫻���ŋ����4/�b���~��nM�؎��~Y�z��k�ߺ��Y-(�t�9_�r�1g�B)'FN���?��>D�Cjy���q�e'V���kՋ4_0�r٧z+�X�{�PpO�u)�:@�l�u�X`�*7���=��4���+�O��{%�N���"o�tִ5($��Nn�����������k��o����ٙ�Ki�4g
vE#���?�V;C�z6GiE�.ǌ�,n��$�m�ɍ�� �.��W��D�G+��8qo�;���#�F�%-��C�L��h�
$�7p�a_޻��ת�n��\,U��>ODNH�ט]2c���+&�`Yo8���K>���[^�h��9�Gt׾׋z(/��P�ۋ0�D�`�D�9'9s���o��퇯|߭��}"��
oD����޼L�үp�0�	B��h�#3�@QӋ}��}0��#a̒dJ%�Ƅ���pj2��*���hb��#8�lj6�Y۷�$.TkEs�ϸ.��V�c���E!�]���H��"Km�,W�G�mE6"���tM^�D�V����
�z�{:�T�"���G�ޱ(
=c���=m���N�N}=��C_���N�nk��?Q�^ϒ���5q����.�K��J�iz�E�:\Gk#���F��s�Vz�����5�GGZ�q+#ۯ��	�g���$���Fi<0��B砨�w�	�|2m��vB�����H$a�b�T�;��4UB���m*�����j�A?��DD�_�l�8%G�c�WV�ξ�t�ƥ)$  ��1�*qrޢ�������B����#է�Q�C;����`i-���RL/j�nZ~#��4��f8��������M3uM����#�Bq���Q�tj0�����o5�-|o+�*�[���n���t�c��s�5H���𡹅�wF����C���P��BqQ�m��tɄɘ.t�_ߜ;���Ւ�aX/�.*�{�k�N(F�ew�ۤ�z�����F�$�hf��~˕��5ǜ��6�X�� �t�������,�h�B/3��M �m="��xb7|Ќ�S�L.M���eBc���w������8|�ڮ�;OQH2RD��H��L#��mշ�A|�D���j\���G�L�gj�pj,�9IP"d�p��I�a�*����x?0��jN��B���Ś�S���_NE�O�V�Y�gH"����j�Pܺ�H��R�ã�l\K���. �`{bxv�κ�6�8�d����i�G@+�YTH\0类�;/�<��4�KK���9��W�E���é��if9K+OI�y�x$F�5���09Zzg�xP�r5���N���9S�3#��e;���b�wO��Q
�9�����T�9�B�0k�o�'&^4��*���ܸ�'$�/0�J`��2#����b�zt��>��R<���:5��XקM���(ɭ��ҁ4T��o�m��`ޒ�4���5��n��Ҹ�V��(���y�S�95��Vg�=a�Uݻ��|j�WKD4C�*��r���&+���F<�����{&�R(�P�u��]�{DW��8�x����{B����Z��W���7x�{�&w�t�S�F_}05?C�#��՛kj�/�מG�:a#�8�}���O�#� �����8�P���z�Ю��'���I៝p��WUW�����|Ӿ���S;\���j�׋H[�i���^��;z�+��������o����)3�س�%�e��zfW��;׬��N��58��,a=m6��l�"��.��X)¦�_�� hG6S�B/w�\:�ɔ~��hE7iw���v�?�HY�<���M���}���@��_p�3^~������#�{�>x�_ޱ`�@e�P�.��֬���fQ�Ü���$�&���.��)�0���xq�5wL��6paplD�A�Ә�V+�����y�5|R?l�y���o�F��z�o\���-�q"*�<h��s��=�E�K�Tl��W)(�K@\,�C�m땱x"y�=��5���d�ʬ"��V�D����#�n����o\�%{��'�P�߾ş���4� �^.Ň��T�B���xaK\Z���i��K���q��-�8I=��2��,R?�4�C�֨(�O�-����AL��SZz m�=Wj%�^򔠩XEA����c�+���{��w�Qݟ�>� ��}b��6\d��F>#H�t�>]��e�K[=T� 6Q���y����&�H�\�;���x߁�қ n&!%ӥq��Z�M���Z0/Z�;��UC�57�����*Ѕ]�$!�9��@θ�#�ԐY4\�}�?�գ9^�H��R˯D��~V���|Փ��K�L�������Y����,���ڧ�:�a�>�C@��=]F�Es���m�%T�œ�f/���E���"�IwJ5����(\�ҋ �v�]-Y�:as��ǡ��Q�'J��!��fqI]z�օ04���>�ʚPCCf1h��X�$�Q؃�1fn�u��Ycj����|��p�8h+^��}3�9�,+o����M�h��Җ�U�ز�;\pM���f��������H�c�bXU$S��#��7��G�d��j��AM�]�����LW�5$�9��⤴��P�I��q;-�]NZ+�&�� -�Po+�a�2TJ��̣�(���ϖ���#���H��?�\�,Q�Kf�C4Bp�f��on)�/�+= ����Wn�[[�)��o&4S�}�b�#�Im���5��י�i�Zd¤�Y%2O�����@$�%�&���>8��\}��T�rmGIh����Oھ/���,���t�OK�[D�҂6��@<�܌RRf�<���!dW�k���fS�t��i��J�	Kݡ�UQ�,R�sȓ������t<�����)���X�Z�01���6$4d�Ҕ�� ��i�OD�
c����Kr��f9N(�W�4�:���y\�t)d,<��!���d�&$�ܽ�ͺ�V�.�C�v7��8��;K��N�.E���mn��Z��;�~�T�p��������2���n�T�"!��ں���7I-��]w~����~����!�e1�e"�S�Ǆ�Z�/����)��ӂ��޵wǺ�<�Vο����v���c!�L=l7��4��4����b׃7�޹��H�����<w��+*���Z?��J�17������l,9*����ޥ�,��ٶꪙ[�A�鍂'�r#��/ش�P�tߍP�frFd��K� Ҭ��	�p�I=�K�^�����%7y̛2T�la�J������y� �g��l��
�\����̹|d�����iis@R�;'�e�{Ka���щ�%�a�^�N�-u~�K��.�[pZІ4ٴ�"d�#�c,x�Fs�����8�ⶐ{�f�iwG9BA�. ,�/"82�<~�e.�y!�v-
�� �3���;��2��63��91SS�ƙ�j�P�+���w�j���V��i�)�Ԇ���d�.�whOkO�e<�F���ƐѴ�nO�VG���j��o�w�|B�qS����z�ޜX��D)��j��AA��h6_�����Z]�ik��*��G��Gy}[;%2L]����JTE,T���{�AK޹{���ͫ�~��ybܲ}ؠ��������o��^V�z��e�2Ng�'d�@s���~Ot;)b��;Ś��l�G����u��!�s9�_�{������8h�.E�ML�dN����)ɽ��,� 0w��J�G�"c�n�A���u%�� S�	L5h�n|��6�X���u���*�=�7V��k9��[B��^a,ڪ�6V�%���㹤m~��7����"��U'[��?�\�:���/�;5"���{�|��׋B���Qo�HPb4��`xx�+FF��c�Wa0�8�j�O���Gd�~ں�ObN��%�7�3�@;%g`��8����DQ�9J�^��Vt�T*�訣��1::
�wx+W,�={�0���d����TE?ج�e�벧�;�, �3��ں���0:{]������d�i3p��-�D���4yʑ���C9��믿��s�=~��_�7<2�.���fu�Bu�?+�8��ֈ+V�{Uq���Q�f�hm?LpG7�͖5fK].�,���`�^.t�!S�W��`����I�C{�[2� ����(�$���8L�^�l�-��r�E�y�k8Zk��{�n(Kp�q��֭[�\�x����s�B
n�+2rsҿ{ȓt� �'=�W��|Ԋ�{N}�a珎57|���_;��yǜ�zś6n����n{���^�쿜М5�߱�K[��:�����ڇ>?0P���α��u?���o>�䃟��_}�c{~x�]���3�{����e���M����\�ƿ�?{Ȓ���?鰷�n�u�-�=�h���F���<Ֆ1��H`q�(�)2v�򕯼��G�Bdw�q����h�<�P��a�!�`dddC��؀�i��g�s_���֍���������J�{�����G���F���b�|�׾q��u/xN$�/�ع��������a���W������ǎ��q��vͭ\y�.~�Q�լ4��ܷ��η��*[���g��s '�~�_�@���+���u�\��D�m�����y��8:�w��7exd�����k�<��C�c�8��c���/��4B���?Ж�я~֬Y�ۆdΜ9Z��8 �����vo+R�n�[��1ZD�{�9&'������W����Dpص}��/DSSD�����b}j�T���#��w֡0ը����U���8�)�+w�#��(�\2.��:��?��2�k��)�h� ��wТ%��K>�����b�RW]u�FƧ?�i�3.��Bx�ᇓkr�E�X�����U���Bt�s#�{L�ϰ0�'^hDh�I�:E���)Vk�a�y�h��LYc��FB���X{�p�I�Z�����=X?�:q�ޜR��%�p�m�mp�%�����I'���x�0����������)�T�r,ɨ=C$�y�۪����4F�M��%�Tg�u�X@/P��i	6R�6Z��\�'i]A~@��C��E7�V�5�8��P��#��(',H�SM�TfL�vG�T[�X��Q 9]�:�ٞ�{fWK"�Řy���݅ju����`���!�nxD|8S��t��lH]f�+BK�Iv�L�t��I,;��@�BkR����G�r�ǚ�R���`�ڬ!��B�'n�'k	؄�����C�,h]D:�Ecf�l��i�|��q�2v��#��M��S]s��}4VB�|��q��l�YC���:�D0��3���a�j�X2�b]K�y�,BtV�7�e.4�fbS�Y�!#L�S�?jE���\��f!hX4>�\i3gѵ��]-a��H��(����i���9��R�RPi�yI���5��ȕ�3m��4��#Y��b/ָ�1�9���$�g�N�$-A+d޼#�]��ˤg0�Y���ٕDbH�f�[:�bo�B:�ǖ��u�̲�e�P�
�uΦC�dw"��ĥ�d_�gz�:�q(Oc�5�HS@�����HS��l��#fD1cT���y���ܹBkqO6K@�6=S1Ͷ��3�L]!8���c���%0`~gv�5��䀔�"��s��>���!����>{
^�?X�UM=����.C�N�cu�2��d����/6��_C� �����Kh(q��a��<�GO���O�E�$om���/���6M�?���<�Z�;*�b9	�߿C�ɶYe�N�N6@�Z��a��btD��2���i�`+�d�"�i�-T��ɦ�M���F���2�@��!��0[m��:t���h�璳�@iiW�[gVV���l�����5J���h���y:��El9��T�q��Um iʴ�L�Jdv�v1!�@&Z-_��Ԑ��2�2֬"��Ͱ�\���6�N�bm�P�?�|ZK3ݽ"��%��#�,�,�����"X���X�6�`c�5�w��Do>�Ѩ�� ?�gv��yRd+��>��U��\G�+1s:���fQ1t5B!c��v�s'�/N��B胭�ۦ�gTrH�"d�y�=�G�	@���)e���d�Mh�V�H��2~zҾ}�9j fz���L�h�\%$����j�+ee�5��6��r%'s�$Sfٔ�qgf?���Jo��t���0[fܖv����$��io��B���e�8�Ikꌚ�>I�;��z�L	B���3��R��:�0�/SCy	�Xի��L��DQ��6�I<�m�#`f�)K�ȥ�@���%�0+�鍃u�3qm@�7����G`Ȃٶe���B7��x;������B�����Y��%cq�q�ˤ�S�]9:1{�۬!Ĕ" �!rK�Ȍ��3b,���>�T(��y�W�6�����r'*���$c����=�� ����"�Ӿ͆�h6��:�E�&���kt<SWH��gJH
�+�v!����eu��2���;�(��<����f̘CA�����lER�S�T~��6�*c��"���q�l�>���j�?�V���~YIK����FX7�H���G��f�d���LJ�۔9�������@`*3'�И+"�鋛�{lx�WI�B�Z.e��vߔg��.E��d�Nj��R�Ξ��vg�6R���	�r�� ��C���7"iR�(d��q��*�gd\������H9+�����lm �Y�+� �ƤTo�lL�fepa�i] D�O����La<.m�BYo��+d��'��V�Uk�2d-�.��2��Hx4�1eR���%���ȴhNZ�9�S���A��h�\uf���
�Z�R�1�qH��]8�j��1w���2���������5<���Ӓs��l��7.JS��5+D�t:[7�� �3��H{�{�|��NJ�h3ɵ<�{EE�&�`�z��y��)^�����fOS�@k,%��l9"\	c���W�i[�)��E�P�ᦘE@eL�,
��uc9&uDU+}�èm���b�%B�h:���H��aK*��QO����y�0��a��P0U�f����Z��̢_=<'?wyK�<�G���V-�T��CN�T����W{^�{�!ԛ�����Zp��qb�kN<�d�;P	�����*�秬z߻�s!fn1�OT'�Q�Q��̿6o��z���YAHOO7���(t���B9���nX����|b��_��o,��%r��#��]�}����H�@����q���>��E<R8��ǭ|�V�;�y+ja�׽�g���J��%`��ms���/-�������u�W�^������*�u����ɯ�>�E�����F�j���۷kN�5'լ dx�(���������0z�?~��f�cs�R�g�|蟾����e�?����{�E�4t�"%����v�H3���}�1��+�`�K_>zч��/�H~��;��/�e~#�?a��[����)���o��[Y���;��F�_˔q��ö����w1w6ڬ �6`��N?���:�~�D��񩈬���j[�tWU�y��G���W��澡��Zy�k4������$e�G��L@��H}(4�z�}�4��jm��������YAW�!x$&x�%�L�;����<��䒳�_�rYhi����ڬ9��5ƌ���g��
B�EX�����"WϬ�T
�<�Ǥ5v��@�?����2[��BH[B�I��Tk�k�B��r�Ob��6�KdV���{�+RfuP������lO�?:��D� �	��>��'sl�ڬ2u4O<�Yς�+W�5�\�+5p^�����n�M_���3�<��^شi�>�t�R8�S�}Xfۉ'��ݯ?����o�^�*صk�]�V���W��p�M7��А>�j�*8��#��k���J@�f�dI�駟�]w�F6�a�HpA��җ���ߟ d�ܹ�X���?\#�!��H{��G�`�3�8��!�/�c����L�m�$��ں:]ө�N�dIS�z�IY�"a7n�믿>G*~���0��?�)l߾=9�w�^��ꫡ�H�"����w�N~#�o��f,�C�ӏ~���1�[�+��qw觱�^�;F*�oذA�e�wܑ\�}F|w��������yL��u7�pC������>w����HI{f�������dHғmO��#щfIS� �eKr|��3P��8�(���޽֖�#"�ZE\�o�]4M�y����$��ϧA���lN�����N�ά S5��7�ٴ5��0"�d"h0)fk��H����rćXF@,�d�	]x���u�&b��c���ȌsH�O���G0Ԝ����
V�.E.�J�H�P��a5x�����e`i�a����
�Ϧ

�;���Ԛ[&�$�A���#T?��1,��V�*���Co�T_1��1�S���Ȩ>�#��(��T�U ���҅����:�.�(*���ݫVѸ�Ru�GPR��L��|Z�9"�
ju<� 9W]�cx���}����X������=u��B����y��σ�h�q��aJ�Y�-&?KG�
�c��4t�d
���t6��$����
	�@�t�yL��z�����	�ޙ��y�:�MW���꿩�Q�qOwܳ]BWPP�E��z"L��c�&��z3��>�C�YAH9(B/��uw}f�,	���˾2�#j�nW��@�c٣ �C���`B�[��Ľ�g>)+�6�WS���P��zB��/�a�+��ȥDnQ�*�##�wI�&���O�d\]Q*�{��Yپg�-X�v̷v�ZU_��SQ���6�ݯ9�ս=�^3>�f줚��j����]K~��ڨ����!'�Կ�λ��틼X�}�E/�t�z�Ԩ��|�|�wѩ����r���EjլQ_���u��v���G�8�z�=~��Z�7#���� 3�0Na��h    IEND�B`�PK
     o_�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     o_�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     o_�[Z���0b  0b                   cirkitFile.jsonPK 
     o_�[                        ]b  jsons/PK 
     o_�[rfƣ�  �               �b  jsons/user_defined.jsonPK 
     o_�[                        �{  images/PK 
     o_�[P��/ǽ  ǽ  /             �{  images/0b351edc-7875-4477-b820-546ce15be531.pngPK 
     o_�[$7h�!  �!  /             �9 images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.pngPK 
     o_�[���� � /             �[ images/bf314729-9196-4b76-b154-4ab11fec66f9.pngPK 
     o_�[Q��0�U  �U  /             t images/a88da2ca-7e0d-495e-a5bf-cdc1eeca5e78.pngPK 
     o_�[�c��f  �f  /             j� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     o_�[��EM  M  /             �1 images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK    
 
   2E   