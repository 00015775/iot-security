PK
     �]�[���4�|  �|     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_0":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_1":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_2":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_3":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4":["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0"],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_5":["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0"],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_6":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_7":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_8":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_9":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_10":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_11":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_12":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_13":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_14":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_15":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_16":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_17":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_18":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_19":["pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_1"],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_20":["pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_2"],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_21":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_22":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_23":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_24":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_25":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_26":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_27":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_28":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_29":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_30":[],"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_31":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0":["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_0"],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0":["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_5","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_3"],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_1":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_1":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_2":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_2":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_3":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_3":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_4":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_4":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_5":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_5":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_6":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_6":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_7":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_7":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_8":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_8":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_9":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_9":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_10":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_10":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_11":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_11":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_12":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_12":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_13":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_13":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_14":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_14":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_15":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_15":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_16":[],"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_16":[],"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_0":["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0"],"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_1":["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_19"],"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_2":["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_20"],"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_3":["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0"]},"pin_to_color":{"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_0":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_1":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_2":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_3":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4":"#ff2600","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_5":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_6":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_7":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_8":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_9":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_10":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_11":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_12":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_13":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_14":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_15":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_16":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_17":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_18":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_19":"#FFE502","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_20":"#96d35f","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_21":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_22":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_23":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_24":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_25":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_26":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_27":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_28":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_29":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_30":"#000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_31":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0":"#ff2600","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_1":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_1":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_2":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_2":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_3":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_3":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_4":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_4":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_5":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_5":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_6":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_6":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_7":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_7":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_8":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_8":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_9":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_9":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_10":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_10":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_11":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_11":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_12":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_12":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_13":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_13":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_14":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_14":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_15":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_15":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_16":"#000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_16":"#000000","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_0":"#ff2600","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_1":"#FFE502","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_2":"#96d35f","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_3":"#000000"},"pin_to_state":{"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_0":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_1":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_2":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_3":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_5":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_6":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_7":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_8":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_9":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_10":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_11":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_12":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_13":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_14":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_15":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_16":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_17":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_18":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_19":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_20":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_21":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_22":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_23":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_24":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_25":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_26":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_27":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_28":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_29":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_30":"neutral","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_31":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_1":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_1":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_2":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_2":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_3":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_3":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_4":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_4":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_5":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_5":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_6":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_6":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_7":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_7":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_8":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_8":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_9":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_9":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_10":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_10":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_11":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_11":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_12":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_12":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_13":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_13":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_14":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_14":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_15":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_15":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_16":"neutral","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_16":"neutral","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_0":"neutral","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_1":"neutral","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_2":"neutral","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_3":"neutral"},"next_color_idx":5,"wires_placed_in_order":[["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0"],["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0"],["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_5","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0"],["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_0"],["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_3"],["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_19","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_1"],["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_20","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_2"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0"]]],[[["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4"]],[]],[[],[["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0"]]],[[],[["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_5","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0"]]],[[],[["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_0"]]],[[],[["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_3"]]],[[],[["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_19","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_1"]]],[[],[["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_20","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_2"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_0":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_1":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_2":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_3":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4":"0000000000000000","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_5":"0000000000000001","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_6":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_7":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_8":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_9":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_10":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_11":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_12":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_13":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_14":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_15":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_16":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_17":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_18":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_19":"0000000000000002","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_20":"0000000000000003","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_21":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_22":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_23":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_24":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_25":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_26":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_27":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_28":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_29":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_30":"_","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_31":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0":"0000000000000000","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0":"0000000000000001","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_1":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_1":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_2":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_2":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_3":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_3":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_4":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_4":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_5":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_5":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_6":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_6":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_7":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_7":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_8":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_8":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_9":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_9":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_10":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_10":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_11":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_11":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_12":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_12":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_13":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_13":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_14":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_14":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_15":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_15":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_16":"_","pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_16":"_","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_0":"0000000000000000","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_1":"0000000000000002","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_2":"0000000000000003","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_3":"0000000000000001"},"component_id_to_pins":{"431bb9eb-13a9-40b9-8288-d29dc7f633ad":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"036be6ab-6325-4263-b477-7689cac6bdd4":["0","1","2","3"],"c934ab84-79ef-4ab8-ab64-87e30b03885e":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_0"],"0000000000000001":["pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0","pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_5","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_3"],"0000000000000002":["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_19","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_1"],"0000000000000003":["pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_20","pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_2"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3"},"all_breadboard_info_list":["cf663b0e-137e-4ebc-a058-da9e925d582d_63_2_True_1210_130_up","3a19d390-e0fa-47cb-bd71-db8874730c0b_17_2_False_685_280_up"],"breadboard_info_list":["3a19d390-e0fa-47cb-bd71-db8874730c0b_17_2_False_685_280_up"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[1101.25,402.5],"typeId":"23db5403-7550-740c-a02b-8b3755757442","componentVersion":1,"instanceId":"431bb9eb-13a9-40b9-8288-d29dc7f633ad","orientation":"up","circleData":[[1082.5,545],[1097.5,545],[1112.5,545],[1127.5,545],[1142.5,545],[1157.5,545],[1172.5,545],[1187.5,545],[1217.5,545],[1232.5,545],[1247.5,545],[1262.5,545],[1277.5,545],[1292.5,545],[1028.5,260],[1043.5,260],[1058.5,260],[1073.5,260],[1088.5,260],[1103.5,260],[1118.5,260],[1133.5,260],[1148.5,260],[1163.5,260],[1187.5,260],[1202.5,260],[1217.5,260],[1232.5,260],[1247.5,260],[1262.5,260],[1277.5,260],[1292.5,260]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"2e7dec78-3909-4d6d-8f08-f82815e4675c\",\"explorerHtmlId\":\"5efb6b6d-ba3d-4243-8693-2bcc1b9e11e4\",\"nameHtmlId\":\"2a28646b-98bb-4888-9d3d-b3a4f1a25b0b\",\"nameInputHtmlId\":\"198e7804-3b5b-4fdc-a31a-6d1e740a11e2\",\"explorerChildHtmlId\":\"83d3f653-fd8e-4084-a5e1-72e2e22275dc\",\"explorerCarrotOpenHtmlId\":\"994764b3-1ddd-4a4b-8ea5-6f8655af55d5\",\"explorerCarrotClosedHtmlId\":\"a43685e6-4256-4c0a-948a-ac933c1680ba\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"c4f183d1-59ed-4dbe-8638-2ac1df25c968\",\"explorerHtmlId\":\"1b6b7a0b-456d-410f-b5e2-3e7cfe69dbdf\",\"nameHtmlId\":\"e42ffa7b-bd7e-483a-b724-968982d87e4f\",\"nameInputHtmlId\":\"db881c74-4793-411d-8c74-c50b477c3849\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"9839704e-077d-4657-b881-3770539d2d55\",\"explorerHtmlId\":\"1402ba2a-c209-4f04-9116-6a0b05a14171\",\"nameHtmlId\":\"42d6a1be-fbbf-46ab-9937-e08e42291efd\",\"nameInputHtmlId\":\"186899a8-ffe4-484f-8d72-4e729bfed361\",\"code\":\"\"},0,","codeLabelPosition":[1101.25,245],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"SEN-15569","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"SparkFun","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[717.0136135,88.496435],"typeId":"f7a95729-a811-496b-83f5-7789de376adf","componentVersion":2,"instanceId":"036be6ab-6325-4263-b477-7689cac6bdd4","orientation":"up","circleData":[[692.5,155],[707.4992245000001,155],[722.4999985000001,154.99530950000002],[737.4984445,154.99374950000004]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Ultrasonic Sensor (HC-SR04):\n  - VCC → 5V\n  - GND → GND\n  - TRIG → Pin 12\n  - ECHO → Pin 11","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[980.8046875,87.19999999999999],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"c934ab84-79ef-4ab8-ab64-87e30b03885e","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"8.79601","left":"573.85321","width":"758.64679","height":"561.20399","x":"573.85321","y":"8.79601"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0\",\"endPinId\":\"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0_0\",\"rawEndPinId\":\"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"647.5000000000_290.0000000000\\\",\\\"647.5000000000_282.5000000000\\\",\\\"587.5000000000_282.5000000000\\\",\\\"587.5000000000_575.0000000000\\\",\\\"1142.5000000000_575.0000000000\\\",\\\"1142.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0\",\"endPinId\":\"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_3a19d390-e0fa-47cb-bd71-db8874730c0b_0_0_1\",\"rawEndPinId\":\"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.5000000000_290.0000000000\\\",\\\"662.5000000000_252.5000000000\\\",\\\"692.5000000000_252.5000000000\\\",\\\"692.5000000000_155.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0\",\"endPinId\":\"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_5\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0_4\",\"rawEndPinId\":\"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_290.0000000000\\\",\\\"812.5000000000_222.5000000000\\\",\\\"1345.0000000000_222.5000000000\\\",\\\"1345.0000000000_575.0000000000\\\",\\\"1157.5000000000_575.0000000000\\\",\\\"1157.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0\",\"endPinId\":\"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_3\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_3a19d390-e0fa-47cb-bd71-db8874730c0b_1_0_3\",\"rawEndPinId\":\"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_290.0000000000\\\",\\\"797.5000000000_252.5000000000\\\",\\\"737.5000000000_252.5000000000\\\",\\\"737.5000000000_200.0000000000\\\",\\\"737.4984445000_200.0000000000\\\",\\\"737.4984445000_154.9937495000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_1\",\"endPinId\":\"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_19\",\"rawStartPinId\":\"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_1\",\"rawEndPinId\":\"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_19\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"707.4992245000_155.0000000000\\\",\\\"707.4992245000_200.0000000000\\\",\\\"1103.5000000000_200.0000000000\\\",\\\"1103.5000000000_260.0000000000\\\"]}\"}","{\"color\":\"#96d35f\",\"startPinId\":\"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_2\",\"endPinId\":\"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_20\",\"rawStartPinId\":\"pin-type-component_036be6ab-6325-4263-b477-7689cac6bdd4_2\",\"rawEndPinId\":\"pin-type-component_431bb9eb-13a9-40b9-8288-d29dc7f633ad_20\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"722.4999985000_154.9953095000\\\",\\\"722.4999985000_185.0000000000\\\",\\\"1118.5000000000_185.0000000000\\\",\\\"1118.5000000000_260.0000000000\\\"]}\"}"],"projectDescription":""}PK
     �]�[               jsons/PK
     �]�[	���Z  Z     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino UNO","category":["Microcontroller"],"userDefined":false,"id":"23db5403-7550-740c-a02b-8b3755757442","subtypeDescription":"","subtypePic":"0b351edc-7875-4477-b820-546ce15be531.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"HC-SR04 Ultrasonic Sensor","category":["User Defined"],"userDefined":true,"id":"f7a95729-a811-496b-83f5-7789de376adf","subtypeDescription":"","subtypePic":"5a738b76-89aa-4728-b8e5-f09c859dbb14.png","pinInfo":{"numDisplayCols":"17.75472","numDisplayRows":"9.29339","pins":[{"uniquePinIdString":"0","positionMil":"724.31191,21.31240","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"824.30674,21.31240","isAnchorPin":false,"label":"TRIG"},{"uniquePinIdString":"2","positionMil":"924.31190,21.34367","isAnchorPin":false,"label":"ECHO"},{"uniquePinIdString":"3","positionMil":"1024.30154,21.35407","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"SEN-15569","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"SparkFun","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"ba153158-cccd-4fb1-9320-38bebad1b7f9.png","componentVersion":2,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     �]�[               images/PK
     �]�[P��/ǽ  ǽ  /   images/0b351edc-7875-4477-b820-546ce15be531.png�PNG

   IHDR  u  v   ��:   sBIT|d�    IDATx���}tSwz/��$۲0���Mblc0fB��3���@��0�b�!d�qN�bν'�tAgڣ�rf��i��Ճ���M�8�Ms�z��� N�`L�~��-�/��ClE�e[/{k���Y+kY��O��g?���S��ҡ�D�P�C���{HDDDDD�;����_��{�R�=�p����V)v9""""��Ή�:�t(I�R�)xZ�Q��5�cR�GBנP�@��x�1�cR��+o6I���t�|�&�I ����W��ǙM~��<>/(�^h�J""""
O����=�p���`T��F��:ix./M�8�IV�0<<,�0������ ~�}�M�Kb�J�/^:���Q��)��ӣ ]��+���!�L-[�,(q��~cP�Qx��+u>HT�*�GT�K�N�F#�0�����BN�T���@{��c�NQ9*���!�S�=�p�n�DDDDD��abg�{�aR祄W��="""""�G('v�~I�v|b��
[�M�6ן)�B�;JX�&"""�^�N�dRDO�f੅�`�b���y��A�����DF=T*~��"�bb�������_��g}� �L|v;>��f�@�|y`��6��~�PN�JU�Pث�B�GIDDD^B1��^Jx�PI�g9������~�1��y��\oo/���@�Z����80w��Y���G'Q�f
���c��	��0����'�C
���䎈��h�P�:�aLv��0�Ə��8��/�ҡ:m�Ҡ ^��٨���w��cqyX˸�˸�Ըb����q7��
B�b�J��X���Z���qu\e����MRʕP��{`<�}���R�a��A�<�,]�q��G��s"�������m>=?*v�~I��v\���H�����_�W�J�@�g�DDDDA
]1���1!����(F~�r;"""���N���);`W�*���	F~�r���`�#"""

�r�f��0e�tk�f����봯��f �S&&�ݮC�RA�R1.�2.�W,6����O�P ֋�y�q7��I��f��b�`xx `�Za��  � ��������"��<x��:�����e�?�S `||f�FGGKllRSS��!�2.�2��q�b��1:j���H��R*��?���\�e\�<n8`RG����`�Zq���ޅ��?�6�������9Z-���/��#�uB�)�o�<`�P�B�|ǟ_W*�P��D h��q�?>�v�Wg�˸�˸���B��J�9s�tA*\����xu1ʸ�˸��L���������z��c;Vcn������ݻ���|���>�����ݻHNLD�R	����	L���X`������͎/&&�y��]�����BZf&������(�k�Z���?}(��"<����8f}��6��1���F�oV�[���pa�P(`���q�q%�+�@.H]/D�q7�qCYd���fý{���ڊ�`�Ղ�y�H���%&c�}p���� ��#QJE,���0������F���`Q����b����ܩ����)lF��� 7&����q�q7Xq������˸��	���&A[k+�:��א9/��x���`��8J qJ%�J$ƨ`�����������'�=�RRR�z���.�Z��ƕ6c�MPR8.�ZZZ�~�ʕ�D�0c\�e\ƕ�J����;ר�fɒ<Q.D�q72ӟ�|U��Ʉ/._��cu��j��Q����qc
̍�A�J��]��f5z�菡/-EFF�#�"v4�=W#�x�I�ꛦ@�`
�����&�)�e\�e\�X,V�_���~�q7��"��d��_��G���I0wv`��W�1
t11xT���}�O���B{{��1"�ݎ�oa0�K4������:��d�o��a�ڄ�9��&��$�� �T���x�_���＃��nIbE"��� �&�D����(�0��r###�M}=p���`W�A(M�*H���D�u4��?��ݻ��$""""�DLꢘ�f���1|�7��SWWP�����k���gQ6��t��W��!Q4aR��Z[��#;I�� 't�X�ɱ1�{���ٳA������(0��R###�ZW�m"�;�2�r:j��qq���Z���m� !�r�a2�MY"��������(����B�sc����e��F��vxW~�kV눈���|��.
Y,�7��|�C==r�c�����~�vÜV(V��ЫE&uQ���Z�#���N��,N�D�݆�S��J�
�J���@DDD�b�@4��ݥؖ�,�Y��5O�C��`���54`�ܹ�Z���
�����s����{H�'��9?>T��A'Ʊ��ӽ~nll�!�q�qe������u			�˸�BqC�� �L����z����_H�X,�tu ���m0�X��!t~�%��^QJn
@7��C�^�N� @�MY!�q��Ұx�b�~gxxV��7H�q�qŌ+�����;V���Ì˸�+s�P��Q���/��T���/�P<�Q*�Q����,�PB��.N"%��@������D�/!!j��q�q7hqŒ��������{j�:�J�2.�7T1��2��혫���phn���cm]��~'�PB�B�����=��WU(��K/��^�1.�2.����Q����˸�x�P��Qftp�PȾ��LT
��^ht�Uj��h����^:��P(���u�J����.�			���^Mkf\�e\��5�X
E��!)�f*)�2.�70��2C�3�'�J���.���(xZεu��!�*]LLFGG���+�x�v;�2.�2�$qŢT*#���q�\1��211*����ƬT
�G��P���P��/^n
fܹ�*W /r�͆��Q��ĸ�˸���v�,�g\�e���5uDaJ�b&�F�t()X1���P�Jc�����E�ؘ�(�*Y��B��J���nΏ�ؔ�6G!""""q1�#
sBb7�Ǉ$��oʙ����(ېh��j4rcF���,��B�@A�Mِ��������])�x�P�æ(~�����w2�����:�<�������a1.�2.�J�A�<|�rیω���q7��"^9{)��C%1P�	��K��?��Ǽn����+z�իG��~��|y��	Q�-���	Ld/Ď��I����%9n����Ʉ�f~��@���ʡ
�BiP EQD3���,�+uQF����/>Gl|<F����G�v;�͐{aK���1P�Ѿ��'v،C�Û/x���ĩT�
����Qx`Re2�z|u�#h�ڐL���vL���Z�B=�O+�|Z�w쯼��ݎ(lm6�\����

{�(Q(P L�%"""����.�:�ڝ^<��>�R?O��&��		S�#Y����;�?P�v;,6;�=���P�i�Oʩݑ�8N��Z�>��  �ͷq����#"""�hƤ.����M��ۛ^=�؎՘+�ǳ`u�?�-�B�Z7f�#5�		r�h���4��� �Ä �m\���.�2��,��`�Z�����Iu46m�5�������CDD���A�{�i�3����*�P܌���۠��?�{(DS�4jԾ��-��.@��2��I5�v�PV���t�ㅙ�0���/+�'""���J]R'$ ��߃��fHU�6�s�h�j��B4E�~1����� ��q ���#;E���AY�竺=ې�Q��ݏQw���gBbW�gJ�����$�()�%i�����ꛤQ���#�����U4��`	�����I]�Z�y3>�������H�6F�6<U�W�y����6��Q�� P�w�3�[�� �a�ԕ�03�oECKǔ�7u����h����X��3Wd%��$�U��P���V�0[��kB��IΧ$�Ez$͉��B3�zM0�;Ө��ك�O���G�؁�Y}�rпk9�:6?�f4�t�� �9% Z:`�o�}��1���P����(�#'U��7�a8�i�n(5T� �T������R�π�]����Iա��է/OIn�vJ���Caf:*��(�L��A��I]�R'$������e$��b�����2a��j�!q�rV�$�؍ӈ��t�Q�|��4�q��}�^??ntK��J[`�1��[U;a�o��TI�03M�=��.�"�@W�F� �]��8V,q\��t�$/��b�����9�Iա�j�󮼐 U�_���-h�Daf:��lsܬ��.I�FyAJ�fKrq�� ��B3J�`ܽ	m�&�w�|��+�B�!$��bT�_����]��$�%yYh�ډE;O�d���1�p�ؚ<��_��B�]Q���B���)�����s~�m�&g���HҨQ��.˿CR�(ңzG)�zMh���o���AR%�rbR����p��e��Q��`�b�� ,6�J��/�"�����'��^�Ռ��x�I|��Ը��� ��+nt�>���:���˜�i��P�w����[��:��iҜx���L�<�ԫ��:	��s�*]����b�P߈���h�쁡����0�����fA����8Ū�+U�IS���ls\ؾ��(q�V���0l~ʭr"er'�o%�G0`�¸{�:{�>��ӗ/m~J��M8\+w�k~�><-J�$�U�W�����g����U��r$�6!�5�7:���F��)��5l~����`��*�^�S��*�����2�Z���|�#�%��(�����?�	]����ڂ�ؙ'&`��P��͎�+����^%vb��&�3�s����Gб�ȹ��5����h=�t�^��4���gO�	�J��=DI^�ǋ�����VSg���\����k�����f���:{P��%JL)�XP��Ǩh�pT�&�-h��ASg���sRu��v�y��1����vK��-I�vN��:��B3�o�qU�v�#BE�����b)��r;?��\q|��r{�����Ϸ���oEݞm0��$i����9��k
ڍ:�����^�O��o-��(�NH��?z	��7�@F��:����Yl6Xl6<��z}PbF#�+�l��TqgJ�H��wocw�_���6�fck*��=f��4���#p�J'֜T�E}��V���rR�n���z��
����sKĎ+�f/4;�r����V �zMn�[CKrR�S�����dm[E��9�q��b^��A��M0���V-��b��n������3��{1�}0[Q��ǎX{�IV}5�7b`Ă��U(������0[��TeMҨk7E�Ć&u�y�����������I_��yX���{�R��g���J��%vR����I��	�_b�K?F~َ��|���:bO���iHr�<����6���]mA��RwoBCK�V��X��<����C��R��e�����ݛд�nu�;J��ԕ�WjBr��Q�di�#����B3��ls�w���>V�_�;'ޙX�y�?0b�m�p�w0[a�Ќ�T�֯���j�5���0��PV�ܣS*7�a(+F�ي�3W��h)/�s~O�|�B\C� n�;oX	�_��I����Q	��N&�$�I�:*ۓ�/���(_����Hä� 8���j���~�0��+I�q��	&�
<��V�$$ub%���+�kb���5���Q/A�`�xu�t�l5ቶiH�;J���O�i��tęr���	�/��W����3WP^���-�><-�U��T �)�U�v$)��-q0�7��܀�*��.W-�u|�;���*li"�6�7����/4;�f��%VBYx��VT}x�ys	�d7w��\AҜx�t�����K�r�|��g�8���,�ñ�I���ZQ��<�B(܌��j'>����r \$�z�$�3��wl�j̍~�mƥ�%l-7��h���=Q�����0n�#&�Q���	�����{�3u%�=v�44#��[̔�(�FG���#K��ێ�1K��v/X���&i�h{mϔ��+�d��<%u{�9�	�֯Dݵ[nI�q�&$͉w�o�".�m���ׄ�w?F���:���H�`�-�3���>(���C��{��J�4'^�q�$'U7�1�	[P��3j��A����_�
	^�>/�r/l{!��TF,S���3.0��Y�~%��e=�� |�#4u��|6���,�+u�F���5�{��܌k�|Z�s���N�d�f�æV���ǲ?�C�Nn�>���1Y�&<�J��S\MW�4�����d`�"ZBmӐ�F0u{�9���0��n�6g�W9)Z�,�FI^�dӢB�1n����dO8Z:B�
�{������ӽ.�_�lǏ��P����*ؘԑGz=2~�:���q���	�qq�%%�n�atx��a�'<_H��혰�a�c:[|<����d�ȅ�{�T�gm�-���<�8����g�8�)��t��>ga�]�$_DDN����/����S��e�����`�b��4�S������9|s�"�{�C��F������v�Y,Ǹ��ݎ���1O��%6bޢEr�I�R����bb�������_��g}�߿/P+��C51Ԙ�΃�l���-�Y���ʊ�����$R�]7[�Nh�`Jw8��G�4$O�w0M6\�1���(Zp�exj�#���{cc�]|����LR������ہ�۝�u7O�뜺hQH�7�]˳�����s������ΰL�����q�g��{}&��[�M�x	ӳ�O��ݙ�����~��;�q=6�u]�S^���M������R�]7ݴ�$�ڹg��Y�S��q�X��|%U����g��d��w#�N�F~Fηv-f��'��z)��ԑ�ع2��$�Ŝ9j|��9ѹ�g��3l6qo8���0G��Wmw<�������fO��!n�(/ȃa�S���"6��tp�:�.@s�}��|+�!/?#�+� ���j/ݐ<f��'��z)���E����P�Th���x��=��B9?]U����F��U��u�~q��2�&���q��Ձ��w]!6/_��Wc߱��� q]ﾇ���b�'p���o�-y�q��E<��2<�jYT�'�ߋ�[ס��)��kr3 &�U�}]�3�P�w;��q3>��ɋ8x�d㐋R����j��s�O����R�".���_$�E%yYh���l�!eB8����$��q���|k'v�s��B�B��lE͹&�w� ���ηv:�h8O\���Z�G�6����gp���{�9g�'o:aL���:"�($T�=ڂ��J���|�ś�w�I|k���E�yM�7?#mJU�sּQ+I���ϭZ6��-���Lꈈ�����FU�WN��^�y�h�ϸ�$u{� ���,Gv�Źp�s�^
��q-�I4}/jvn��XVr�dSm���2}�պH��ʤ��H&����=�$�;0b	�F�MXrRuAm�ϸ���������}?**�b�êJ���-�[�,jΓh�^�۸��y���Bo�-z����A��8�uݴ�9��m�7��7T0�#�r�� !�}Ͼ�ix0<����q A��i2{�Ed\Wf�Ǥj��DW��+�����\�578��uT#��L���;�F��V-CG�P�.z��<����i��dRMì9ׄ-�\�.��A�h�V� &uDQ����T*��
T*�����װXş��so��I��TJ�`�"\��+H1�]����T	N �����T�����ͷe	y���,xU�h;O���z�v9���0+?8���2��ȩ��F�I]��Y>���Gg��y�wa�\uF]������סP��P�����4�Q��~�l�	���i��$g>z�� ��>���mbv�j�������Nː+n�JҨQ��9�:�TA�F��Mn�ih�@��Ge!�3��q��ͬ���nv�:�:(��z�D��n��d��|\����4�H�v)`RDm�Ch���;��G֜�ٟH>��l�|g@�a����<����<���;���6H Q    IDAT,$͉��}2I����-�v�LҨQ�g�c��ӗ�~f�oD[� rR�Ά*rOդ�s�l6/_��Ϡ��e5�=$����{hl������k{���W�'�v�8y���?�_ock��鏮-��w���Ps�	�cZ��#�:""��`ܽɹI���R��}Թ��� ��O!'U'�vEz����	����J�f�di6�:����N���e�;�1��j>B�>����?(y�h;O�����|4�~t���h����D��:""S��0[QQ�w$y~����(ң��G��K�f��f��0n���t���)z��F�EU$�on�4�h;O���F���PŤ��H���>}�Y6��۳%yY�>sE�΅I���n�lE��+n���"I�F�F͆)�N�bתe0����|#���������o��cDD<L�\\\�^4	�%8���&$Jm.SO�d�03]�ꜧ1L69��9&t��N�:[|?���X�F�,����jl""
&u!*F��J5}�>�(�ʐH�
EP^/Q��>}Y��j*���>�$/K�M�#���N$��ߢ��-ؼ|1��fmz����i��1Q�aR���P��������oJg6��9o|�	��A$�6��@ݵ[�*]��������T�_��<T�����&׺�a��ŲĖ�)ɇI]����\�+}��K]}���F��0�o�Z�aE��^�O_���%yY0^hv&�9)ZG�ˇ���y3�=���  K��L��A�(�tDD�I]���i�_���AsHT���j�JT�_9�c��FѧdV�����AT�a(+v�Y[�	��Fne �5���JN��An� ��\���D�]�����:"� 0[=�U�����-��ڂ�T�s���^��Id��f%��?�ڿ���IQDbRGD$���#^=/'U��i;ö����k�4F��i�(�]�����O��HCVr"���s]E�.���řIQ*/�C��%�f%\���3�  �]�"�u/l�MD��03Ezf�;g�q�zM����K��E��<wo���-0�7�M�2�ބ��[R}��w�֯DE�9��o�s�ٱF��n���S��L&��i{m��}�\5u�x]� 
G����d.'U��^���p�]�Q��w�àe{�9���^���Y{�#��uO@�Q56E'9���"=�w�:f��N9~I^e�(/ȋ��I&u��̕)�f�ø{��lC�ύS�����^�=�۳9)ZN|���P��U;QR}d�4.o�9��۟�^ۃ�^SD~�&�Z���qpL�du.���V�;�	n}�6���֮�%u}����)YbQ��+��(�;�a�a+���,��ن��+#�bǤ.J4u����T�(u|��8�K�P����O�]l
���v::�M��}�$/�Q�+�C�F�'͉w��Ä.��^���K7�.6E9��$�������M�=H�p�Pä.��8Od��<M�l��Aҟ����#�"I5��ls�l9}u�n9+ܳMY&""
Ur%Wf+�Vf��xS4I�v4 ���L�HN� ���p��Q�++FN�M�=0^hs�DQ������>IDDaN���x�U�W"'E����M�f^����K�ύ4L�DyA*����������﹖��VT��1eŨ(� �w����-�>}��<��M��.f딵tD�"��FE��y��Q
CY1�Qؓ+�2�7b`����Փ��-0��4"�8`R��֯D���S��D��QJSg��>�$�U����Q;�U�Q���)���g��0^hFaf:J�]e�VʊQw���QX�3��>s�g� 'U��usĂ�Ξo�"i���1��@��/sRu0�ބ$�zʖ�0[�1�><�ܾ�zG);V�������H�Ҡ�H���+��ك�w?���DD6�M����t�������$��?���+80��p���?,Gݞm+iު۳����LV���l��w?"ѳ�O��ݙυ{��ۯ�7w7Hꮶ��j��
^^����t&uDDv�K�b]3&i�0��03U��x̊"��Y$΂aR烵smXk��ܤ���VǨ#�N[�ɱ��mU�n�;۰{��!̝fBRRt��Q᫶;~�����f�˸20[�w:���7��]1f�U��B�_V�m�%$|Ez4�t����y��I��~�j��Z�q�Q�R���������!��KN��U�(EN����MҨ���P��Q��N����*F���>���	���䬘U���hܷ��ݛ`��r$q�W:�Y�E"&u^���~�slԺD�q����Ά&��#���%�F���Z���	8���T��圮�%��2s�����7w{�S(����|#w�L��4�;�W�zM(�(Z:D�j��yA�T�(��Qw�I���''P�~<ܲ�[�N	d��: """
?rW�\��������C��l&uDDDDDDޒ�b�:�L�V�(u&���� �oq���*fR��Q���h��A�ύ0^hƀي�w?v.Aj�ډ�"�dc�+uDQ���Hиw|�^���C�0.�$�3a C}�ǥ?���)��;J1`�F�>u��E��{C�J9���:(X�	s������&G�l�lE��Gg�� L��ԭ�X�#�R�{�`��ݮ��9K-D�o;��H���df+�O_�r�iܽ	%K��4+/�CE�%yY��ꮶ����.Ԯ�_�~�[�jO\�XW�(����(�c��U;a�oDCK�v:��=����F4u��j�JT���������nݼ���
�I����ԡ;'U���?���᪢H��<Y����b&��+��BҜx��MҨ��Q�/�0�#�R�rL�;U���h���PyA��BN�n�}d�d�P��h��m��9m#����^���i��䡩�Ǒ$�T�0�����6>O���7��{
�M�=HҨQ򰃢�di6�V��e�%u���h�5����L��MN��W,���q�¾�Ez��&��\���i�#T�f��૜T��>��(���sw��E��K��/����dUw�����H�r%(�LwV�\-�B���U���0-�P��hn�R��P��&A4��9�:�䡡�f���"�����)�7&'����4կ� o��#�g����-��܎���&7s�sv=��1�����%i��
�l���&W�;J���s��p͞��>���
�4�H�ހ�:""""��]mA�槜2O*��h�왶�2y/Z	chh�pTU&W�Z��2�q�a���,�v&�B�Vw�e��?�ꐓ�CÉOݎ��ҁ�<f�;�ϭ>s�y��wor����Kv��{�C (�<�j[�p�\�[ ϯz��O��b��Z'���t�i�m�&��ن�=�7$�OnL�"Шz4#�݇e"&V���sS��>�jb,�q������3c��$/u�nI:�
&L��vE�Y��Φ�H��؅����4n��U�
3��p��m�eCKJ�]�Uw��m
f��%�W�������2%U�|1��q8x�"���]O.��Gq��.��e�}��g�CG�Z��x>Ea�\[ߠ�1�.�L���+&uD��e�x��$���ĳ�p;� ��w^�,���EX���Ci�j\""�ʹ�+�C�^O����zf�_�ufBu��f;�֯DyA^@S���{la_�~%�֯t{��j�]�Ȧ�geM�
UɆ�gϵ7YCK��rVq��®���Qs�	 P{�j/����L�]W���;�]���'��|�Y�Z�b�W	��B�䛁W���	���(b}���˪N���A��;/��  ���������5.���K|��t�,y��r6Ez���9s�ʖ7rRuHҨ=&��L��Օ�e�-E����}����n��L7ƺ�-0l~
���0[��2��j��
�d�[;q�uj���}'�㍀`��}m��<�s��E2&uDL�krB����`$vL�HJ9)Zgh�!L1�JI^rRu�H�Mi,�4'~��,ꮶ�03I��4N�6�9���칾�%���.���S �����E8���:��ΔXI��1�#")��9�|�0M�x�ٱmA�S!gC[�	�~����f��$5m������kKա���?{��s����j�w�pt��$����*iN���n�ȑ�y����1a��H�����r !!a,!!!V��^zD?2fW���#���?|D�1�;����7��N�fK褊�Mb%EbǄ���TQ�G���0^h������C}#��7�:3�9m1'U��Ι��~_LO׈E��:��K@M;����w���vT��������E�>e�	d���������P(Rl6[�7�x�b���h4���[
 q
;  �_(�a�4h4J ��Ð���x��i�YG:Ψz�\V����N���n闟�������ݛ���g�J��B�W	S��+h�t44��9���2eSs_�����U.��l��p�d��:]zJRZ:`(+�j�_ݵ[���t
3�e�|���G�
�X[z�+�O���6��^�����INN����Wm�
7�Lꈈ�䒤Q��/+P��Ѩ���E��N�JK�3���,��r%"""��!l�0ymI��������������I:Ez��):peE��{
�f&tQ��:"""""�0�JQ��N�";Y+�0�����z�=�"l�s&uDDQ,?#�{�C'�P�������>�j>���.f��#J�|�0Fu:�l�)���f��A�j_������>cn]��#���hX�#�pm��A[�i����T�sASg�c�Ym�+��(/�s�Z����f��n���z0`����e��'i�0��mJ[w��������&��z�8+uDDU���c߱�rCTLꈢ��x5�t���/��S���0��03�~�|�𸡾�ou>nܽ	�ݛP�QO�e�o��
��Iա��� ��=� 8:�5u� 'U��M��a9J��` ��F�������Z��#"���5uD�rRu��Q���� ��\AҜxT�_��k�����U0^h���U��1�2�Q�~�W퓫�\AyA��P��i��03U�FSg ���C}#��l��A��7���A��ADDD~bRGe�֯D�F��ӗ=�|��I5�4j�z^�Zx��>�o�5�03��騻ڂ$����:�4'ާcE#&uDQ�$/f+Z:<�|�l������-(��Bݞmh��P�,'U���Y��03 �������LꈢLҜx�X|���<����F)��b���&)3%h���z�I��xEz������IDDD��Ѭ�VG�w?vLߜ��Y�~�Ǧ(��bʊ����T�3�ބ�Tݔ�~DDDD��:�(30b	h�����Q^��槜�T\;UΖ�yb(+FyA�����?"""�h'߮�D$��k���Q��77YyA�s����+1�7?r�ss;��/4;��4;�qwoB����x�c�}��hfLꈢL���0[QU����'o.4T)/���|��I��v��S�����?@��l�TaBGDDD�#N�$�2f+�><���{�6��SeŨZ�-Ω�M�=�>sŹ����9Ͳj�JT���EN�ι�x��G9咢Nv���Zd�$�m �67�c�\�e2[q��>���k_A�F���4�g̃N����A|��=9��u��:�(Tw�%�&GW���xSg��'��h�5�� m��q>����H��RYQ�G�F�8��8\�Y���~�(�g��L�ks3�� ����_��`ڟ5�v�\k'�o�z�=��*�F�|���f"+9q��)���i�2��8w��[�"�=��������BZF���'��t�,š�Өa��#��_]����4Ծ�Yɉhl�¾cgq��ޔ�w��d�bד˰c������w���[��6>o�k¾cg �6���uO  j/}�|�u���~��'/N;v�F��[��U���?�'/8��؂����®w��z�=d�hQ��)�O�Z�)X��~#b�J��V�|���������O�?��R�@���_��ɏ��DRQ��Ԕ(��3r !!�k�N�P���~�t7�r�(�}�5j�,r{lB��X�bUP)��o�u|jK+���bhb|O[>~���H��u�(��Κ��k�2���V�w�ηvJCj��\�-�\l^�X��w������5Ed�L���[׹%X�V-Á��ܞ����q����P�q�����p�'/�%э�](�����E�s���7p��E\��
�c<y��oLy|�����}�+�q{|��  ��������_!?c�Ǳ��c���n�����7��s��9��"��o���-n�TG���δ�����
���a��_���]n1�q�o~�L<;�����Y�7G��e���/)f��X�#""�'����p{,sI.�sf��x-!6�w����o&�P�%�ZŐ�6>ϭZ6�z�t5*�b�'$KxYɉxqm!^\[����8|x���ӨQ�s��=��������Q:n�L>W�s`Mn��&;y�X�1m�|k��Ǘdz��c ���X� ��؅�ɳ�G�5��Sn���k���@JB<�-��X,w^*�O��ޫ(Ê�#��>&uDD��AF|U� ������^��B��~��I�t��q��8��i���9�$�8f�d�}�<~v�o,
�ؕ0��d�����p������xs딤�d��d�N���*�k�s���8�ډA˨������?5q9���qJ�[���}�㞎8�E��V�c��}oʴda<��p�鷍�]n�����Z&�6�}J��쭎)cl�?�-��)�g'k����޹�N�tR")��lْ�P(*�@\\�)>>>I����}� �-�r�HU�W�_��?�el���}�G�M�&���%A�Pa|�
�Ō����A��>� �`��c�{�F�W���f�~�v<S����Á:F�?xl!��q�����_�!p$��/�������O��{�!��dMn&�� u�
:���B�~��wܞ�x���"I�ƪ��`�2��?:�������7���Y�����͆�w7���|k6<��F���.�?E��.}������څ�N�gh���X�$�[����;�L����:ׄ�'/:�ҝ�:}׻ﻍ���˨�|�ۿ�8�K���;�S����|�|kηv��>��-:�����_��?���������9�������}/t=C#h�@Y�b(
��@�q���.����Y�P(�34�m_�F�5�*�����q��&H)Z���t�����?����#.��Q��:�dU�W�PV��fﮞH�\gw{,1)���n�����I�Z@��a^�b�'L��;_��2�r�G��	SߤZ&���F�S�5w��HC���g̓%�7��%����۸zʚ2!i���63!�6g����MY;(�ף��5uDDRF'�KY�R��Xb����p��-$ν���ˠP�_��K~F��n�m��/6/_��?y�GN����D$�.��Wv��MGX��ӨQ{�\��ų���n��4�pg2[�$k�SovonŮ'���U� ޻�?+7'""�R�e#!1s��	 �զaђ����t\�R1���8�Ņ~b#�]O.ùW���N����{e�ٹa�'� ;E���
��N �G'u^�Cv���݀��Dh�����B���x�e��[皘 ������>���.��5���m�s���L�$
+uDD䗌��ߊo:�����FO����ڧ���V-s�W�dS����n�͋k����uʪ��[��(��ȹ���}�κ}>�nj��]�ۏPhb�����6���`6[1<t�c#r'(�=��3���O^�8],P�k�^EY�&t�����r��v�R��HCv��c2y<D����<u����'��X�#"��d-�.���u�:t����=$�H��]���e�}��kr8��J񼷗?��q�߻e�?�uk��!�{d2[q�ս5���,L�B�-�    IDAT�Q#?c�3�DM���P_�]Ҫ�������{���P޿|��9�2��^���������?CaSw6�!10�#""�`||f`�L`��M����3f(�\[(j�r���o��ý������5��آ_�2�d�J��N�.�׻��K7P����_�b�G��y�ٹ��9�f�k�2�=՞[�Ǜo#��oI��Wy�*�����\���Jvq�ܺ��s"0�#""�%$$  t:Gu�61�ί?C�|xL�l���mA����8 B���A�^���.}�S�⪣�_���/߀6>{�=�]��T�4��iԨ��.�vR�G��|{������qp�:Iײy�0�g��N�$���4����I�F������jo¼�Q�5)��a���m `��)F�)ڀ�E����ɋ�iWb����ɋ8x�"^\[��W�=�0�Į�bK�	����[��ֹ&<�j�o\�wr���B�k�,�:�b���'l*��1k'u�l���}�7<������{���%v\cG�bRGDDS(Uq��O��wU1j<�Y�{�����;�Q١��nj������lE͹&<yQ�QM�hm����k�:�?�]��nS}e2[q��E�6�Ry��c*��uO���B��X��=�6(�i�صj��sq�������w�\��qn]���f߱����t�cp$%�T,'�^{��hS�3�ܶ��vL3Y�����
g�B\�o��A�(j/}���8���#�pp�:d%'���7�wg?þ���{�*|��%""�hS�C��sal\<2�W  ���a}��v&�h�e��B��������~O!�Ǡe������V�<�����6>5;7x�$Ц(�ͭ�<r
��Q���+��y���[|�lj��pp�:���ܺ���.���oL����in窘�b���~}&�^1�x�mQ*�:�:��	�����	{���O^D͹&����7�:߇5��h|e��gϯzܯs���4 "� ��b�͏<�W����q�����ohԌ���qv��C��6%���KG�Qc�������K7������йjl�7j���Ϙ�ڊ-3>'��1B��yc}P:W��]���;~U�6/��)�a$l�1�����E�L*���+�� �۸�����"d�:��zq�I����J��0��Q���z��;��>�l������ߙ�L��G��;�T�o\�״�}��e*�l-��R�+~vv=�{� t��4�mד��n��7�]��hvٚ@.��Q���{}�?�u�(��k��Jr�E��W����bo��Ϙ�׺T]|�$�������3WP}�J���f��ɉ��I]��N��E?֥U9%z��@������ZC�1�c���~��z�=��(�!�;��.���f%'bד�^����'8���?G���x�m�+�bp������o8��:�2;E�5�����=V��Y�z�\�۱�����:""�Iv�q���ҍ�K�B����Pvx׻�!?#�{��U�ńN0h�.�q�Wn�ij���E~'ukr3�������T��P�,����uX�F�,�����޴9��m�;vv�ϡ�o�}�f&kr3Q�s��ݞ�˺T���nKͯ�&wLf+�:�aMnfT�8��#""�d�'|z���N�� �7>x�_	�p�*l�i	����>�إ4+9ѯ�ukr3q���۸�6��?���z�x5Á>c��]Z�Ө�ݢd�����^�[;��Z�S���߇�(�[;q��E�X�����v�|�_�ŵuaH��F9�2�#""r���e>%.Bӏp���S~��g�õ���k/:���[ס�r�����1<����)����^qͤi{��8����f�9���Em[�y�~����_7=Lf+�j>�ؽ����)Z�)���8���[o�|��H�����c���ɋ�u��G�SA[�c2[E�н�p{	O����q:�&蛗/�����]+�pv��gn����I���ǣ�S�����y�K��S�6Q	Or$vLꈈ��i�3n<<Y{�`Ht��Še�GNy����f��e�C>_���?g ��������>�o�t�pt��k��E��!f�)����yڭ'&��c���V-�Zw��ޔ��q:��<���1�#""zhMn�O��bP���%�2���ِض�N^����VwMf+�s��yc=�7�c���'١�Se���uAٻ�S�x������K7<V�}�Z[V��������N�&�n��`&vLꈈ�Z����}�!���'>���)�P�ꍎ�!���r3`ד���k{���#ܺ.��� BE�}����D��)��L�;e-ݠeT�
��)� ����{��&�O^Ĺ[�x~�㨯��J&I#X��:""��|�8��<�����s&�}����{>�/��8���4j�=鲒��F}s+NL�����P�N��n��7��^!��p3#+9ѧ�)e�\غιf�����7�!q#�cRGDD��/�߻�#	�}�>�qJ���n�''>�������OIK�6¨<2�<�n�1x�as\�u�&�����Og����2��Rh�:����DDD�|�=���A�׋��n�&����Lh����۞�^���֮���7�M~F��]=Ϸvz=�-;y�J���Nt��mV}��-"��lŁ��.�/���XG�醍��Wx�xs�xޜO7�K��{��a���*�>6�:"""������rm��E���7����h����ـ*%�u��V��͹W���g����+Q8���uR�671��]���﯆.^�s7��V5皰E��b�*������ۢ�5�tS��H��4��S����8�p��/o�k
�6$$=�;N�$""��)Oӹ�g�N���ߓ�/��r���ـ�]J���{l).�u5�u����Vv6�c��+)�����K٠��/�}+��@V�܈M��)�e(�I1�I|����w���x�N�ӹ����M#�2}.�W>�}W���u�����"B{���je0�����J]�ߚ���sq��]���lG�{Q�&2$�;&uDDD>2Y"sO����~U0"uj�/�G�ur�ٻ������y�X����5�b�]�I��k=}�&o�0��[�9G'i�����:"""r�Te����Q��Gܧac�P6�&�/�y)����1�#"""')׶E�Ó��5�vEl��W׻��I�X{�I�EJ���N�׏"���:"""��s��\�ʛ���ͭX�s#�����BY�GAY�8p�":�ݛ��1��S%y�[����]��8��m4�v���7�T2)���qK"""�g���������� �"l��c�_��&7��/��0�{����u�ZG�д��}o�Y''�J~F��s�Ө�����-&3���<r
�+�q>&��uR���[�0Y��o���F�] �0�#""�o��z��Г��V����Zq��zr�߿_�s���������4j|�ڞ���_�z�����WQ��󾍫a2[�*a����N���66/_�|,н���F�씩7|i��Өq�'/8�4��������E	;N�$""�o�n"m��6>5�6�M�Qc������ƛ�F�^_��y�`&;yj��E����|�V9�vs н��F)v�.X�a��/۠T�-t떩Ϙ�]����B�ǟ��Lꈈ� �6���H�Ey(�ٹA��ʵ�(�db�2��ٟ���^T�<%��C�r+'�ي}�>q{,н�<M���ٻ���;��H���e!"8�Xp�d0�f�T�2"����=A�dfrj5�����`������cMrƐ��(g-r	V0Nl.��E�`ld���ڒ��R_��;�����[?���r�~��<�H����<�'Q�wK�_P!ъ6��  �"�bf�y�g������+�,��mј�#X+y������ӽ:`Ц��X�t��e,�^D���'��x��We4��Eya���F�;9c���P�/��h�� �+����;k�~�"��Ƶz���*��灻�g*<r��:?ҭ	��P�7��;^xY�O�;��������|v��dT��<sf<{�S,����7|�p�$;�����=�Ԗh��Ǵ��c������"v�:  �8�L3O5�)+�k��BvݺV�xP^F�v�yh������*~�a=s�����zC>�Gό*���3򔌑:i*ܼ��3�źw�ۧυ����|5��=q����w�=֕�ЁǶ�ÿo�-�Wh��"
v�:  ����}�����0Wm���Ѝ��<pg�ih�Z��f�7��ĝ_��o�ᕤ'f��3 X�蝹f+/#ݐѺ���z��>l����9k=Z�{ׅWO���
��.p"M}mF3���c�C�?��zC����p�`G� ���'��ւ���I^F�<�=��N��h��%���myံ��i�?[^8`�3�����Ϳ�k̺�x��4'�>�A�g�q�'"�jj��oה��4�y��9}oe͠ue+�Nen�<�(�����k�`G� `�h@�����*��{]o���L�ڞ0&�u:���sa�9=m�C�Dx{�F�9����!��}�v����F�֕��3�6�,�軤����/��3��̙��W<#b���ٜ�	=3�0N$fO5�kK�|��P �4m�����i�� /}垘*]:��ㅗc�s]�
Â]����Q.	�f����HK���~L���-}�7�nH���_?6�㼌th�mT6���j�H��_?�����;��>o\S�[W�b�F��=�ˣQk���hb��hԡ�C�`G� `��_?���n]kȺ�D��;j�+��x��ԉ�K��r0����6W��z^�륦k�<=�n��~����������״��A��������"��W��{oW�_�3���N��hǈ�3gf��ٵ�`��޸Vo?�+������S���#�{�o��b!�5Uj��%=���k���*������I��
��l۷o��X,�jPzz�HFFFA�������1����n 9�ׯGn�|T?`�}ӵ:;�S�a1xx�Z5��ӵO���P�ק�O�j�>'���}�����7]�W?�X�/��$JMY�~��;��f�꺽o��_��l���u�Z=��u��Ks�tq����>�=��>�{n�TinV��nS}M������ڕ�.-TEQ��33��ժ���#�~^�޻I����-U�s>�=C���r0��ݖ����{'㪜�=�ԵEya���F�/�^V��3�uin�vݺV�k��۔�f׈�#�קue+t뵫����ڻs���s׆�{��ׯ/���G�W[�����>���<U�j׭kuནQ��a��H��?��:���Gkt�z �L<��Q����c�o�lІ�Fx�+��<B���:0k�ቾKz�翉�o�?���~�E~k�Jb��tOD5N~��g�[�f��Q��Wն�Ks���e������z=��=�]�.������R}MUܣ�������k�J�|T:��U��ը�jK��Q�o�>�/,WF�~	 @8�=��}ݳ(�h��H�+�9�;�z��Ԟ�V�+[���_ZU�btRl�fk��̜j�oP#좩�:�ξ~տ�ꢙh�4Li��x����%�k��:�I
{~���|X��a�%�<�_�Չ�~}m���Hm��REa��>����5e%:��v�}ӵ1]����O��;�j2����nԺ���gS�Go\���ᾘ]g_����1�~����L��ghT�>���rm��ڶQEyq<�קW;>�ۧ{U��PuiaT���������z��.�^��FO�:uqHwT�Ϩ����麇����;��y�1W���?����~,��-U����Θ2��{'����bj�/˾}��V�T5 ;;�l~~~l�u�<��N�R� &�̽���*SS�JjY�x�+MM����bL�,9#.����[I������g�rS�{�9�	�j��%m�6���;�~���Ж�r�++�-�W���y���:���^C�_EQ�*
��N�]ZS8�SQ��'�U}M՜"1�t����̙��-U�:��v�e�����W���[,��0B�<B�x��a;Z�=��_?jHI��l�Z�}_�'�}�b	,�M�g�ߊV��SϿ~,��Έ>z��o��C|$����3>v�'T���'�YXغ�Z��dF(
��x�xlFp�պ���|?�B)  \Ů��z��]��>������h��I�t�C�����z����W�-���
sD��(O��G��{�^:ܡ��ް�N��V��{o���^~�d�]8��> S�e�1��oI��� A��a�c����k�D�%�u�����1��U����J�7_רS�S
������v��ۧ�E=ʹ�0�J���1������^��{5��,d׭kC���	}󧇴��
U�{ȩg~�֢�����+[��L�N�]ҁ��3F�������P�%�P\�#�tך?�������望�R�����ŢQϤʬ�����������d��D�����=8��!��]�᪢0O��)?ӡue%q�6�f���L��<pgB�v:������#ij{�[V�PEa��T�6$��R�>V�uh'�.i�C��X����5}���=���?���z��	�0�/$��;!��`���4����nB��Z���2?}l�IW_��5.�<�H�J�sT�]���옟c�Xd�X�i��б��9���co{2�軤��^5<�m�*��pF�����vEy�(��at"%3�IS�58�rv�x�u"u*��f/��H����v�?��g��7�r��ict��H֬r���d�Ŀ����gҫ4�'�j�ߍ����?�G��0��A��x=��H�O�����jo|(�s;�]T]�+j}�A�U�QS�5���
2jo|HY�k~E]����}���˞�#) �,�H�W�#�u~�1�R%Q�.�^��v��FB���W�����bڠ|1y���)A��SL��(O��{�*
��o��>�k�����:�w)l��p�G5��U�r�������{����g���{���W,�=c���@@���# O�P��b�U@u��'�-�: 0������oPS�fu����S=3^o����,�W�Oތ9Ѕ��9tV�.�QFf��)�)�[|ۦՋI0�xl�)<���pGB�q�ݓ:��o�>2r;�X=���{Be���[j���Pn�Z��¼�7�Gb�^���7���?c�����ڦIϰ���~`O�UzF�����R�q���X���5�c��O���O�z�Ԝ��7�q��?���"�=[�O;�W���u�����KW���-�/<��EO�-ȵ�,�@�EJȲ3B �Hǹ�*���f~��Ӱ�35J�s���7�����k�[7��z��O���h�!m�Xm��3%I%�*��9tV}���▘��L\Y�d:�wI[^80���b��ׯݯ���}��}4{m�b�!���t�����Ӫ��im�*׉�KZW�bN@���\{tL�n]Z���]j�y����e�k�w�~߫�փ���K��&<����I��ǆ���#�4��{2d:����g���뫵c}�Z�ר�'o��~��j�'�%C ���,����j������%5�>���b�6�u `2-G;UW�F;�W�y�65��MՖ���~��F����yNN���^5�xኛ�;ߩ�K��h�u�<ˬ���w�Q���3��YО׏�dDg��Ѯ�U_S�=ܹ�G�9%5o_�������ۣ=ܩ�����-e+B����:�}�o����GN�jW��9Ӳ��{�Zo�
�W����5��jxxX��.�ᰫxE���	oC0�u���h�%�[7�q�F5l���x�`�t�����n'�k9 ������l��F_x�EO�mͳ[�,ғF�S"��)�\æ�?���͡���fW|�Z]�=���ߑ=-]EJw��n��bY>�)����ۧ{��;ݨ�����K��gm�����s�}G�����j=b������E0:���A�^~�d���=��yL��~x�ywG���،-&��	�{n�F\�P��ٕ�?|����Ј�3c����B�XW�B������p�{|�����*=q% �t�#������d�    IDATu�Z=���q{��/��F����v�QU>���!g�k>?ӡ�wԆ��{��A�=����O]��������Lӛ�Vk�Ƶ:r�wƿ/����S�?]o���3U�����\Ymv�9/�\��UPP���jY,���,;�W��zMh}�l͇ޟ�~�?�Pæ��3[��T�Ԛ����>�:��.�)c�V_|j�)5�|co�U��w�&��	�<jz�jy�>�>����o����%��b���Z��z䛼�1���̑�jU 0w���D�%��{U�n]�g�ݔ���>:������,#.���~L�wLMI��Ji�s�'��[�jM��W��Kou��;qy�tO��G�{B�5��XÕ����w�N��N�vb������{u�T��U�umQ��T�Y����_dL/��j�F\�}t&��	�軤k��gs�jm��SI�s���ܢue+f��RU�-/P���Ϩ$���\�ۯ�wԆ�o����ޫV+?ӡ]���V� �1����{�O�5��j{�Ka�W޲z�v��S-�`�
K箅��[������wy�Z���Ӧ���z���{~�8I�����ڱ�zN�kj;��G��23���w��uz�᫟��~�5�[{��~k{��.��� ��h=~*���k`DMmG�ކ��J]�N�I��^�vISB�=�_O����7̎��=���;�[�s�v�?���t���=�_{^?��~��?~C����]Љ�Kz����tʗ��`��/�����go71=��>o�u|��V�	��k�TQ�7��#��ծ0[\l�Z�-aF�wm\��53�`�e���0O�gmi����ue+tǬ���j]ي9[`��^�k>�aij�qKUy(�Mn�鰇�|^v������E8�7�5���]�=�Iψ�3.j�K�50r�"&�~"Ia��I
��;�ھ�B��������}��k������� ��*��UwcE����	M��e������}���'C0�m��ӄN�
�GZ�T���k�+o�|�e��#w��)Q/�Ow���=�I���1m����m�茜�ۇ��u8�����>����u|�J��3��{/���+����<a��=�Ԉ;�}f�]��.�uI���z��M�}��՞׏���j����[uy삡�-�t� ӡ��]�Ѱˣ����V�B`����eFH#�G2]���>�ᗿ!�{0� L��������Tæ�P��. ��Z��e~}�{R�%��ͻ&imX��>}nj-�+o���JwTMM�="���Q�軤{/��ӽ�v4.Z�~���#�u��aG�"�tO�����a�%�u�IZ��T������-/���u�	��[%L}���g��qy�ďߘq<�����;Bk�z�FC�ئ�������{d��C#d�}����ȭ��}8r�W�=���33�����I�軤�_?�-U塯���P��S��r�x�==��7B#fӧ�N�{�k�v�릿�g~�������N=�ũ_���/���J��^�k1���U$�?���)+w��3c�w*��ڎ��z��nP��݆O�����y�.Co��~�5�/�k�B �PS�fՖ������t��M5j�����%�~�?��m��Hekn��s�9��V��V�#[nט|^��F�~���p%�}��� ו���Iq��3�O��m�EX*�jN�]҉�K3ʾ�*�_���<:����S��{�vzi[�i�{�\hs�`_x���:τ=���^U��8�����K�;TQ�7�ks�+o��׏�9^��U�+[!I3B���9>��h��������R�=�{n��\)|�'�.����{|�s��~�O����zo�{ZJ�N��is���3���SZUPF����;��L���݄}���B�4��)���O��f셧Z�a��^S�����:B �L�7�]#�@��YW�&T9,�i9Z]�Qc�^��=!ɮ@�+�-���IҤU�u�O�ե�C������42�*#.Oد���wΝ����FL�;>�ߍh�'��.��ْ����K��>�Ν�@��(�`�q��ר��t��\Fp�ѷ���z�ڱ�Z�[7�ն�<���@��ŧ�O�m�X�����5u `"�������4�o�w=B2X,6��W���MZ��Z�y9r��]y�*i�my  fc��U~�t�����+��5֫��Sr|����l�E���;��`�Y	�׆G��x�Oޜ*f���@@?OŴ��F_x�%��)�: 0����?�@��Ȝ�d���Q��g�TKs�++�L9y�dO�Qzf�` H���1]g�ٵb�M��s]�kt�3y'���M\��i�[Ԗ����9�k�[7���!U�ݣ.�a�'��ymyiT�	�o��}�D{�/�$�nm��F6[pyp��|�E�b��]�:#�$t/�ͦ�K��
 �Q^����^���Y�Z]�^�44����S�P_��}v��gj}�����WN_'���������F��9uk�f�Z�-i~kTSu ��4��w���C�G�bY4��e�Q8s���>Y'G��d���2r�W^�_���r����'$���� �����ʟ��V����r��S�K���l�Z��R��oC��?Sæ�9A���)�~�ID�.gk��k����y�uF$���/6���>Ց��G�)�B� 蛿����v  ���Pqh��O�d���ҭ�Ϻ�d�ov�+���ۡ��٣���W��Ψ�y-��Nijf��A��'P���J���e���N�   ��o�98��')i�Y����T�a�@@B  @d�wnU�j9ک��|Ֆ�������8w1��A��P�  ,k�?yS��^h�W�7�*�P��Ў�Ւ����k��Eiܻ��_F;zH�  �Gp�dI���"�R� �l�:  "P����?}]���uu}���T燞o�nij�)x?D�����H]æ����Xܲ�Muf���uQ���f  ��L_s5}J��a�G]#j�߬���<�n �A�  ��~�g��f�~�G���
���T7�T�O��q�F�%*�Q�d�X�=$� p�奪-/���~Iu�kTY�0�`�z KK�*),���t�4  �*��r��O���Eu�����R5l�YpS\�K��g|<}ۂ��fǹ�Qm���P����������!� �G��5顏�'s4�cW��snN K9ʊ�A�F=�*��:q��y$��%Ip=]p���������M5j޹M�z��vD�;��F�Z��RÏ~1�܆M5��;�]T��筴���y�R�^k9�*�_W�F��?8����FT����q�5l�	�D�<j~�9�g���HS!)�`��H�9�ػc쟟jMu[$��6D}M� 0��֤���B[s��W�y��*�,����Ue��(-;��X,Y,}�y4t�du��e���r;�WOU�tyB��Z?�DM��U����d:���}3�Nנ3���6��-/Uˣ��dD����T�,�t��~��n����v��ᦢ6n�0��'o2�`Q���E�����: �~߄��㲧�H
�/�2����5��f��$I�w�*v���T���h���Kp���G���G���Q������7�	{�VY����|��TS��<�,�W��m��^z��p;=��<jj;���ҩ X�F�;��� ��X,z����JϋOu���O�m�(����R  ���:����х�?�u��ώԨě�uA뇟�x-P")���v$t~pM^A�C��6J�褩i�;~�3u$Zjp��� ����BO�ӧ[����f�ێs��?M�l��ϓ�  &��%�xro��bm��RB �X{�C����io|hΈMp�g�f�M��n��?}=��*�M���;rUZ�N�׮Sz����a���N��|m��=�(S��S��s��pU�n�}��|o���.OJ�,�{��
gӿނ���h���a��8F ���b�]9�ػ#U�ϳ[�b��u ��Ֆ��Yw�~�G͇ޟ�*����\���q�b�HF�r
oP~�-�)�VNA���t��*\q��ӭ��i���,���٦����p#n�Ey��F����:%��g��CA�#�j���f�����*kKַ�&}���o��a����z���"Q��~���`�kܺaF�hj;Z�4�XGA�#4:��r��׬Յ�:{����UPT�tG��v�,KB��l�������
����N�,9��^K������_v/xn��{�0��o�Y[���:���p2������V|S?��E��'o��TO�����$��~s���TY����#	�XlZY^��kV)?7Sc����Z�η��(]�� ,N���٬�zroA�������v��=�i�A���	̷n���E5�QS�f5�ܦ�㧴c}uhzf���W�f��y갼^��m��iF�R��T�Y�[7�
�DZ�$x�|�۫�v5��>:7}�n��,�G �.����p��Ou$�9�ػ�귶��$F� `Q���-/U��H��ܤzz������v�,�����^�ˋ{�H���¯��n���lAܫ���t��Ia�x�����)������0�E��~k{���k4��O�-��Ƌ�6YfD��u �ht}��9�/���xhZ�BO�����{I	
rd�PY�M���I�:/$�ىڛ�T�UGނ{�Iх���B�nm0�|����)\x�Jiz���BdS�fISm&�0��o���=�b{�7���{�ܧ�6�٭�E	�P �\���5������a"�k��~�&''599)[Z����,�P�z�vh�3.Ir�����}Ѕ�?�;�pQ�T��7]��eO/RM�N�mܺA�;���Xmy�Zp�)��+f7jܺA-��q��r�30[p�{��`�kz�Ii $�Ţ���{���ܧ�6D�������ܧ�ט�����~�t���cM ,ӫ_�X_ڬy�=���@װ�&�~]������5u���rTV�gs��|�	Ym��y'd���3��j�Hz�����t�i=~J�WBَ���/�r�S�5�o}�k>�~�Ѻa�G�o�*�����3^�0F0c1���G�Pˣ���8_�;���q��� `f���zW�]�O���@@����uM?���Z,�JTg�h����}�: X��S�ZP-�ާ��aGꂁ@���9����u����b�)7�B����h��#��s�5��Ž���Q�h��CV�`J��z_]�N5l�	��u��Z+9��p�u���h���צ���8wQ�����nPæ�ｩ�Z?�$��1 `&��Xt�d�;�1��$}˳�۷��j�J������>���o�$�\�g:9�Ju3�����Z��z���4��}5���Rmyi�}��nPS�fu�����9��>���F�mGB#s�jԼs�T��W"j��}�Jݔ�ٌc���O٫bzO�M�����^������ׄ{0�z�d�������  �+���"�|���u���`�����T��Ֆ��=Zc�Xd�Z����U��5�/�I�E7�jK��M  `&�_�"���7����6ը�T�Z�����2�n�������oPæ�?u�i�N_��kg;?�urT�Mv�-����z���eM_)Gza�kpBҙ�� �rE��E�k`$�^���?W��ݡ���~v�װ�35%�J�pS7���/Å�?�  @��Kk�R�5u   �ǚ:    01B    ��    L�P    &f/))Y��������8��=K_q�D�   ,Q��   ���    ��u    `b�:    01B    ��    L�P    &f�t����1U���^��>UϏDFFFaFff��?�����⾧;@�N�7�M    ���/�גnJuC��>���������z�����O�    0\    &fOu ,]��"��ޛ�f   ,i�: 	㷧�U�2��   XҘ~	    &F�    #�   ����   ��T��@C�o3�*=_�P�j��G�   `g?PqW����Oߑt�a���    ��q�u}��[
�.���wT8h�h#�   @�4nݠ�m��n)� ���   @�d:����*��P���Q]�]���P    �wn��e��ڎDu�RtA�;
�    H����j?��5e�-�@T��;�H�S�9�Q_�H]��Ҿ��6    fm������d����:B]n���Wz/|��v    �lL��P���5����:9�Nus    \�V��U���7n�G�'���>5�E����f����T��^��qѰ��F������댮R   ����1�S+W(=}n����ٳ�
������46��ʕE�?�T�~��ϝ�P   `	����a��:k���w���+Q��ΟTaav�����$���    ,~������y���|��~6湉t�R    ���   �T?�E����0R    &�H   �%��%τwƱ4�_��i�}���<�3�kKK�s%B   �%⓮:qp�q�զ��I�	X�t}����<ע�Ң�<s�s�    H ��:I��}�8,�w2��1?�2��zn@}���O    �����#8�'����3#�>���:    01B    ��    L�P   `Q�_q}���4~�M#��b��P   `Q*Z���nKu3�o����wk"=+��	u    ����t�   �"�T���N"�   0���
t�   �I,�`gd��$�!w   �$*Z-�6�\:�����ut�   ���^T�k$�͈Y�ؐ&�u    �������+�͈K��H��ʨc�XS   ��B�����r/B   �Eo)� ���   ���]���P   `�Zʁ.(�`G�   �(��~��]P��({l �k	u    ���T7!��Ƈc��P    &�>u    L�s7��]��d��o�n�:O�׻|j���F�   `j��4�tj����ύ8�=:{�W���S���u    � �ΟVaQ����!��w���+1��R��?!�   X"���;/��?��?��f�
�    ���    ��u    `b��   �d�����8�f�+==mI>W"�   X">麠���Zm*+-������熞�л   @�Y�7XI���S��ay��K⹳1R   ��>>}>��|RO�x�l��   ��1R    a��7�aS�
2�Q뇟���H����0R    !�wnS�����sU���ƭԼs[�[��0R   �p�5l�Q��Sj��/B�ZP�j��vD�.ς��_q�r����ܔ�[m)\ӵ��   0\ݍ���?	vy�z�Ԍ�2T�Z]�ݖ�."~�M'o�[�Y1]O�   �4]�Ψ�_��.�@'�    ,rK5��$B    Xj�Ψ@'Q(   @U�i����;.I�w/X<e�h���T��;	ik��$B   �j�����"THe>�`Wr��K���m0,�I�:    	�q��5���h�V~�Gu_���G�   `���5�1��g?Pq���M���.y���[}�!��P
    SX
�.���p�א{1R    a
2j�T��?Q��H�X㶍��^�a�G-G;���n)����/�]Y';B   ���-/U��� ӡ�Ag(Ե>��j�KC��U�QSQ޼k�b�2"�1�   @B�<z�$����?�$5nݠ��R��T������W�q��mTA�c�=�r�������b�    n��jU�����|����su7VH�������P���4���z?Z�.���w�=6ӵ�:    �N�l9�:V��P]�u����))4�W��1��c�Ih��5>�u�:    Iz�zRܒ��B)    7|�-I�,�m*�c}��?�������nX��6W�f�?޸�u�<�w?�4�g,���F�   `��h\��jz�*�th��ju������.�<@s:�re����F����=۫@�؉��z�l�:    ��8wQ-G;հ�&4'MU�j޹Mu�kTY��+CL    IDAT��������u���
��e��Q��[~�_�Y}����	�   @B4��Mu�h��j�<j=~*T8%8B7�����3�^����;/��?��?��FI�s��    $L���n*>���G�P��S)h��B�K    	S��PS�f�U���Z��j޹-��#u    ���T-�ާ��|Is�T競�T;�Wk�~皺勑:    	Ѽs�*��`��ޜ�+����vD�5��f�3�]�pi|Ɵ��IC��+1R    �ר����EP�����5nݠ��5qmL�I���88��jSYi������zNB�   `Y���B�B�.,��&Z�V�����wqX^��#g�z�l��   H����50�3>>}>��|ROo\�Y,ϝ��:    ���`���ω$ b.B    ����X_}�s��P�26�:    ��8wQ��O�q�5n�0�y���O��U$e9cM   ��h�ɛ�,�WS�f5l�Qǹ��tJ�*��T[^���|u�����6����m�ڏ~%�ߗ�'�Ǒ�K�T�t���,Y���[g��P��   �IA�C��6j�-7�Y_�50��?Q��i��	{}���%�<�l���ޘ�'�E�P   �'82'M�H��-�`o���~	    I:�]���Dz�N�|��vF:�P    
2Qo&��q���0�Z�3*�I�:    	Pwc�Z�/�k~��?5��K%��$B   ��8wQ͇ޏ���	����bmZ��Z�r>J��R    ,Fl>    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01{� s����5=�RZz��2?�_#���T�   0�q�8�У���T7e^�/_V mT"�  `	b�%�666����T7#�˗/���?��    ��:bllL�������������@��   $��SZZZ��2::��&    	G�ò�ZT�e�l�,G�N��   +B���4�ʍ��YRR�����a�   bE�    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &fOu��
3��ސ���C���ci�����|�c��n  �]y��+�R݌��,�zzc�k��
=���X
c�����f  `W��T7!*�:,�>cC���   bŚ:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� �P�f�Ck��_Ia���/v?    V�:,�t}�q�%9��   ă�    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� ���Kg\~����v/    �:,�~}�g¸�\2�^   @�~	    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���S�  rm�Zlܗ{aN��߳#��   ��n�������F\~C��?i��%�n�=����\B   B�2qflB����o֐O��   @�XS    &F�    #�   ���    ��u    `bT��i�|>��n��~�l6eff�b���Y   @R�`J>�O���
�$��+�׫��\�   ��_�nw(��|>MLL��E   @j�`J~�?��   �RE��)�l���   K�����)�u�oZZ����S�"    5(�S�X,������D��%�   ���e�X�p8":�������۸�|θ{   q`�%    �#u0����R݌�ݮ���T7   H(B1>>����T7c�ϧ���T7   H�_"n�5�I���S�    a�C\&���-(UAIy��2��_�Y��n   ��:�er�u����W5��    	��K    01B    ��    L�5u �����A����n  �p\��&D�P ��seU��  ����K    01B    ��    L�P    &F�    #�   ���    ��u    `bl> �jJ��o�ָ�:����g:�t/p%¡? X~u R*7=M5��r��c��e�m)l�yџ  ,?L�    #�   ��1�@T�\�*�՘˘�YΡl��������\.��*��D���ONhrx@���2�{%B�k\�?9��˗��Ŏ4��o[���CǼ^�F�n����}�I�Kc�C�>�x��  ư���r��VZ�����+*��\Y�7�\s��ۍz<�(���u�~-��-��<E7����ؤ���T7e�  a)��:��~(�m����T>0���n���oVVV�$���L�C.�K����$��ŋq?o��d�gFF�._��,� ��lY����<���'�===��'�a��7���v�r�-��?�3�p�*//Waa�$͘&8��������&&&��ե���9sF��c
&�%�,������ٳg�D ��-�PW\\����<��?�?�KA�$##Cw�}�n��v�|��r8��H�|>���kddD:y�~�����O?���"�'  0��`�C�xV�������l|��SFA���Mx������!MK�XȪU����k�ƍ��Ϗ;x,dhhH###�����~�;���Gt]���	  �Pg����r��p�je���z�r�\���]�����٣_�V2��4��U�V�G��͛����@ ��VNq�\�������~��_GF�Db��G}T_��Sڟǎ����z� ��Y�.Uk���Ҕ��-#u���x4::�����s��r:�S%�P��&�dggk���)	s��\.}��gr:�:x�;����
"�'  H�e�R���D���JKKKe3�˥��A�^�z��������'�۽dB]��n�����׾�5egg'tZ`��N�z{{500����/X$�A$��|�ǔ��C ��-�!���C���EVV�#u&�~�����y�������D��$�.q" ���z��'��C�f��t4)�á�������v[(��SPP ����ߖj�4�����	  �[�i�P�x,�Pi ������|G��r�|>_[�ժ��Y,]{�*++����Þ�� B�  H�%�6u��ru����K�>������h�|������)�á�7�>�����"�'� �d�,#��E@�mۦ��~ZYYY�	 A999���T~~��y�egg�=���R��O���b~��'F�'  �:B��E@�|�ISoϑ���믿^iii	"��\;  ��	���������T61p���ʕ+<���������Ą�_.� 2���ҙ3g499�={�h||<�y�Vq�?��O  9B]�|>edd��΄&''5>>����ϛ�������7U��4��]�V��������$�.�Ad``@���w�=/� BN����VSSӼ��  H���b Q�$���g�UVVV[����*++Sqq�{�y�N�����9՟��'  ��X�2�� z��'URRb�"�*,,T^^�jjj�iӦy�+..�Ĩs�{џS�YXXhH ��� �q�}���n[������L��k׮y}a���5�\#)��	  f"�����Z?�pؽǖ�ͦ��2����'�H�3�[�Y�&��	  �"�����򗿬���T7%irrrTRR���r�[���{/�����LX ��u B6nܨ��k�O��k����Z��G,�Oc�  �G�K �Ͷ$�X,Kv'�e-##C;w���MuS��f����D^�W�a�=�Oc�  ̏]��b�hrrrɭ��Z��X,���,��V�|>ߒ�����jݺu���HuSR���D������ׯ���G۟  `~��
Kr��|��n�+==]�E�@@~�?�-C��v��o߾,G����K###ڴi��=��Oc�  ,��0�����˗5>>.��#��*�����5�\�[n�e��"��n�q�q݇��bT ���>�/�$��jbq����+�����)������<]w�u*--��>����  ,�P��
r��r�\��wX\���USS�$�
�"??_N�S_��c����)��  W�O�H
��/�˥��IF����UWWS�押�<�|>�_�>���ϙ��O  pu�:$���._����ȝw޹��~Mg�ٔ���իW+;;;���ϙ��O  pu�:$] ��c:fj��v]{��Y����v��nݺ���?�������X��	  "CiB�������f3������:+oKQk"������J���Ѳ��u��]��Q_G�k ���R�gI;�ͦ�˃�nF�


�f͚e�A�|rrr$I7�pCT�џ��ڟ   2�:��R	vf�j�*
z�#--M���Q]C�/��  �aA�ǣ@ @�$#����p(///�k����ҟ   2�:,���<�iq�+--M>�/�>�?�K ��갨�\.��K"*5�/==]n�;�u`���b�O  ��aQ	r��
)�����jrrRn�{��&''�!   )E�â������NA   ,Z��~�=`�w���Y��X��
��b��D��P�EirrRiii���LuS   ����7�����w���?��X��m$�ٚF��,v%j��P*vQG�W�΋�焯jܽ�(�!,��=lv��E�[���L���oþp�C�2��]j_%G�nD'e,%��&��-r�^P3�(��ΐ�~���4���cZ���{� l&r���Ƃ�~�踽�b�
���Cz��I�;�Y�2�eɿza,\�/�ŗ� �@ۙq� �~��;&udZ�t��:"�K�����n�0��,�?�����x��/����u2��u�_���Ů����,��?h{��X��v���Q-�`�K2�Z:��j����Қ��Y}��E���Ç��Ԅ۷o��1���ʙ�z������.ڛ�����8��gB�Nf�g_�_�y�,c:-Jn�:�ű���Q_�	Hh�� S�d25q���ں�k��L�ϬVVV��imll�b��4G���ʙ�zu�DU�?w�/!��2z �^'s{��S�1�����WǦ�����PZ��Z$v\~I��N����Oj"i6B*�*yo'糰r�^��_�k�o����Bu���y�4I��dV���+3������X��EI�:6�rn�m�İ t��<L�X<G*���e�Ւ�d����d2Y��8�;+w>�ٕ����P��ש��@"��<�H��WǦ���Z �U�s�#e2�ZY�Y���8��鬭e�A��Ζ�8���ʝO""�j� ySǢՎ�r~,$�}<���2�,��èK�D�h�Is���U�۷��~I��|���$""�&YƵ��c!��/�%���x�A����_��IH���U������|����<�̧����=""��TF�:��cqY�|�<�wT�GI?��կx`�L&���|��Ge=�����|�t>��v� pr�β��Q�e�̈e���/�˩�1�#jp������e�iii	{��){�W<�|�t>����A���c�,��~I5A�$��P�VWW1==�g�y�t���.�H������/�z<�s�T4�fao���œ눛��<=��ن�_���{��|�'��}������� G��� 89��cO�  x.mm`:}ng\���h���'�կ{���:^ṕ�7�r��u���W�cj�����ف��_B|-�_\�������9������?r���7��Kptv�s�-�#s[����q�?�v�^Ͽ��焫�K�Z��M&n�<u�#��R��ւ$��K�/-J�=�8Z�c��QM��V��������6|uiccKKK���X]]-�y8�YXYY���|E�Y�o��#��@;:;��4k%�{�����\���y\җ��w����7�:}����������7��<�^��$wv��:  <{��mq\�]����9z��7կ��=�n�w���I�u�f�/>���|/����aDc	�[���-�,N�xsW��v�d���x����W����z�����\���Ww�#��� w�͒?�*�ukFF���K�:6�~�b��s���j�,�쀩�{��arr�����/���}��������|fi5��8:;��߮��;ث~R�5����]�(����w5�I�_K!89O�S�R�G���l�;��0p�&����V) `j~!{��G��;؋xr���G�_wtv�7�Z���:�[��(�����$��������]=��ȅ�#��QJy��d���ϏB[ө�x_[MZKQ��֊,c��w��D�I!�N�ʕ+��d2<x� ���wiT��jm��ZΧ�n�Fpr���7@T��k)����-����!����a���M���ݥ���~���A|-��{GIDɼr+j����|�X��7���U�>'³w�u�f[Y]{Ky�+�'gv\�,-ͭL�F��[+�(��l�JM4�� ࣏>���߰��!�"���I���裏��{�5l���|U�����^�g� �ހۛmE���g�l��M�/l�u;{05��pdnK��݅����b::;�Pc�9y����jUMY������E�Z����lC��mDc���BJ}�k]iε��M[5���TSA�:��������7�7�,��`qq�dR�$d}}?��Op��Q�g��_@pr���C!O�n��$ `oi*�9ów�*���)7��X��.�#sp;{v�KUh�f~����S���yy��L� ��f)	X�����u�N��o���5��K�b����Nv��A���BU��_����������uki5m�嗒(�E��u��3�������D"����w��d2��S5��9�����D���|j;�;��4!pr ��H�^%1+�r�U��H���7���F)��I�J���CM�����Dpr�`���F)J�{����եQi#���MG89�Vn�#sN��7<��q
een2�u[��۟K����L��N<u��%��zݴ]c����ӨKت-�N�ҥKX\\l�����
���055���/Χ�{颱��u��=�})���%�?+�U��(��q{�S/��ei��d�ꏲG�X�����rM�1�����-I���N醩�2��Z*۔�ن�<?�Gm���K������J[.�<�xr]�v�sn.��V�s�����J}�Gc	��b�[k�V�tR"Qݥ\�J�.���X,����A,3z8������O?��������|�'p�fիc��&8:;ؐ��'gԆ��	僃��������V�$N�����Z
���E��q�G�mk;O�S*j�+׷��
�:���E��|�':}b[�47�*�� ����RI+t]9˗�zݴ�:�	�R�0�p8���Y�����O>1z8��x<�믿��9j
�'Q��_��M�N�@���-gw���|M15��=�+����=Ww���J+��BG�7ԏ�t������a�Ȍ|���N����Y����t)	���+{v�G�($=}�]�J}����.1����䌚�z����n[Z��^�6�ba��AJ�2�#�mdY�ݻw��3�`qqKKKFIs.�}}}�Z��/̝�D"Q��jΧs�؞(�P���\  BIDAT�)���\z+[�x�Y�#_82���;7;��t�������#�N
5J�M�	��	��4��f*JI�vJL�%������<�_��]R�YS:izLh:�����;>�����^���|C�p9��1�끫7�<����׭�R���.��:u��!��j�j�8�r� @Ū6�H��X[[C[[[��666 I��կ���s����E��{wnWl�o����G^��ֆ��&���u��9���Kx����o�vyy�}�[XO����p>����
�����+�������������/!�+��b�`o���+�!Kd�[��|�'���qQm�����Q���P��w��_��V���,����hH���hii�7��M������0zH{�'��/����ʾ�\���ػw/�S'�f[v�[K���t�;jz����� "�mб��g��X�� �U��>��/�����X���Ckk+�}�Y�ٳ���T�'����Eww7~�ӟ��+�q>kH|-���f4��c������Sy%"jD�\z"�#o�`��L�	�9ܻw���>[�&3% �������B��7��>rP�6:5��{#b��߷��;RǢF���̸W J>��I���j��ޝ�����~�ݻ�������n��	s�\�����'�|�4	Ƚ{����Y�����i��ԛ��R��WΦS����g�N����v|���|�'tI���ID�a���JkP���q� ��rʤ�L�V*u+++��ں����yҠ������hjj������֭[�����\���nA�$�A���E,þ}�jv>�|���z��&�`Z����o����y�Spr��j�o �'������59H������}�`��{N�@��'{.���\zK�$ˈ�Dd.����[�n��T� &udb{��a�Z__������o���|��)��v��N����x���ҎVVV�L&100��,Q4�@<���g��r�O�WTEs;{�9�=�|�\1�ȱl��Ko!��B��	�G����F\�]�N�;Ҽپ}�Ͻ��V|��1�ȜD���s���cSՌ���G F�}<�:2-A I��àH��h4�'�|_��W��_��Tg���v�����~�3�/�$	w���|�(p��p���D4�P�y�7����BprF��g��?r��.�Ԁ��5t���ߏ����lI�k1&�� tX3b��n\�W#f˹q�(��J��I���je��ܽ{�(��v�Ν;����L&������׿�u|����/~a�X���ԇ����%s�{����;�״>>����%�k���*$v-��]VI���R���Licc��q7J�LX__/z]:���b�Ҩ�I�ڵ��bdd�H���UMF����tbqq����*��,���	�P6��;d\�����X����<G#��ڒ$���_K!�,��B��ē�L,��4�$v�s�^��b�;;�%1XiB0�#E���D#Hg2�WCWWW��'�����'�O>�sss�{��f1r555�駟�7��M<��Sx�����Q�8kkk��Tr>wo7�[ng����-�=}N ����b��U�D3t�6|��>�ݯ��H#������`/<}�-�5���ݲ�3x긚P&n����|ϥׁ�F�$"��Y%1�v����~XVW����7�����.�:2Q��5��$�i�^]�������������a�Z��"�U��455��p����~�iX,ܸq�n��h����q�=t�f�Z�900���fD"ܽ{�n�s��Gf�g�K�#��������	'g*��4D�S*e�/4ѽy��|C����9�Mb�Rj7N��1 ���.���b�<�݈�DT�C���3=A�W�|mgƽ� ���FC �F��2:t�m�Z�=�=A�N�M��/�� �J�����u��˶�6����������9Ċ������!<xP�f4� �w~�w��҂��%ܽ{���H&�XZZ����n��n��'�@WWzzz��ގ��ܾ}��_^^�.�����c_)x�Q���c��/����l���`�����a��=p���l%+pr���o��{�Ww���SO�f��ܫ&�J��WA�:<u��v�A�>'��?�������VFDD��2�ɐ���v���6:��k�xA�i��)X�#S1CB��<�;�{�H$tODdY����YEtuu���v� ��������b�ǿ������}�>��3]ǘ/�L"��m��!]$���OeNͧ�b���>|�>��ABWL��M�:GgGv��?e_�w��f�nU2{K��6�5�#sۖ*�A��Dc��؛mjsV	��A� �+~,��xM�� E%���D���nA@ �:.&ud
� `mm��a4����o�z26����ê!������qUc���C,..b5��M@�������AI���:�sS��Y	-����=�F82�m��lC���o���t@�b�v���Ec	u�`82��tD�`˾�z`D���jY�F>�c���<"2� �9A�s�q�77��*��dRG�cBg�ŧ~�O����֍5H��t&S�18���G��e?���~��}�6���#����@ =��.y���S��Ep>���n�[�89 [U�7���_�xo]n<GgGիb�+�|�yO߲����D��0����߈ʕ��e����VM�}?
��C"z$&ud�zI�������o=��-xʰ���_��aߖ�#��8���(V�W��많j�4��M�g!�X�����;5���bGg���������*B�x7��^Q�2K��7���@��k�臈�:2� �$���ՊL&����F����ެ��T1ng�#�Ԋc�A�z%t���-q�J��\U;���Tٿ�r�!��7�`oiR�\��S�LIGgG�^�Qg[*��Wy5�Y�L��,R��.�߉�1�.������S7�ă�3�7���s"x�8��?�M�n���FШ����\U;�����lSv刊\�X�n>����;ػm)s4�@pr�n^�"x�8<}N�g�����I���z�5��]��=��9�f���}�M������D��_|C���;7��*����	�8z�hL�j!�S4�LB��� D�c��fXͩڮ�&�LWw/Z�h��TZ���*�ĵ�x�����9���8�Z�J�����s�7< �� ³w����X��Q�2�ZO�#�\�~8Q଼hgG]$;��~�G�!�C`�Ɩ9v;{����K�#�gD!Z'�~��TϷ��"�{�������c6϶T��*�� x���:}���۾noi��ϩ���~���^�瑲�AY�`o�m���^1���`u�
�YH���F�n4�|O���A&n �S[�+7��Ύ���t(u4��c���j����_�6E��O�3{�����MGt��f\#*WFV���;eI�N�.��3�*,��=z�>�#�S:�j�;؋���}�u�x89�k�LIr<��R���7���^�c�ów�9�mń�ϩv�՛+?�����f&u�+�ł�����;GD�|�}��m#%		��<|C�e߈���[Yf���;���@��M�JN��Q�j�j��r�\,v���I�J�� �U�Bϭ����X�X�����v�Ճc��s14�.OL�4��� L�y\�������͹��_���S�!�֢���oX��k&L�Hs��$1�#"]){E
-G�7G�~#�v���P<�bdoڪ�߬q�H��L�]�]��>�z�S�u;���P�Z]Wx��w�S��$W��٥�:�+�/�SϑT~F(U�����ȏ�z�5�{ng|C���sh:���F��	&��z�;ث~ �,�MG�+66_�s3&uT1Q��(�2��4R�����r�����rtv pr����_���zc���ܛ&=؛m�A��.u9dprF�O����/�8�ju��FLGgǮޣ�R%�_���q�i����4�k)�.OTe�Bٓ:}b����t����^/��_|��
��]{�������h,ϥ��9�.�ԓ�G!��=puw��ݕ=Sts�|��[��}�m]�`�*�q^}�r[�֫F�A�$X,�AH��l�,�2$IB&���$.�� �J�����u�t��(b�?�����vS������>�]N�s`w)��6L��7�\�u���O�7<�h,���}⮴�w9 �7)1:�"prX���	RDc	]MSI빂��܎�
e?[�+�
=�*U�|��l��Ko�����<}N�g����U�yV�{T:�V��7w�`�_�QX�����2��٣V���H;��|�o�Om+Y���tz.��pd�����g;�uv�]��v�d+�U����N�����}Z��3"&��B3��ԃҡV�_֣��N�7��5?�^{��6ڛmp�oG���sh:�=Ba��g5��V&��z� �1�#"������P��ܮs�P�JwKe����U��[pr��5=.Wi6�׍��g/�S ��<e���/�Sa�� �����+��_���wt�˸�B^[:?�eRGDD5���;�޶?G��f���;؛Mb7�f�S����B|-���͓{�m�YO��3�:(���Q�J(dj~�>'��ܤ3�Q�I�R��=���O��~v�2n�Q:��/�����.O�庺T2�|$=T��?r��~� �h,��郒�j�`�[��N�S���g�s�<0Z��s�'�y��LUc���i�9�������Ҕݧ��Z��p�e�Z�k�܄`RGDD5J�\�$����W����-V��(�l7��	\�	���j�,����ϩ�M�!�@v��w�WӤ.K��YT^_4�@0�:���P?��՘�u�����S[�+���
θ�k��F�O� &uDDT������r�Զc�����vـ����-M[lG�%��^B]���+���[�##�#s������Mh�D24��x#bc�9�z��89�P?B��޻�˸�h�����J$�~Y�x���r|C�r@�w���c��!ttv`�� |��[����&s���e�o�_������j�é��TZ�m3"f���T��z\>���P�V���.O�t�q��J� &u�bRW�����(	�rV�B阨Wg7�X�l� ���%L�����|C��l��=�[��4�<@3P�*���qT�2n�)��L�t5??Q����F �22����+�eYF[[���ˤ��teo�e�gy]7j��r��;��٦&����S�SL�`����^�r��ۆ^�3.��j\-=*������?62<U��?��Ƥ���H�0.��z�J�&� �$""""�0�ƛq�lv���~IT3d�daRT���([\� ; �-�3h�DDDD��R:�I���2�ɐ���pq,^�Ұ�l�㎽�Gd� ��DDDD��R:�I�)�2�eɿza,\�cSǢ)   �vf�+��������L�LE�,��/�0���-_bt<�n�0��s�QG����O�����G_ȸ�˸��5J��3��w\����������x��AU�~�k_S�<�9u5��s�V�&���2��ɛ|ul��'*`��q�1( z<?Շ}ˋp����� �2���D�c���#�U������f��f�1��A�t�,�����u�$��x��饌�ƅ���*�r~,�rn�m��0;""""s�4����j���Ts+���ș4�)$�[�_�� d��XJBW��&���M1�#"""2-:�I��$�3���CF����2�H[$���|�WǦ���Z �U��DDDD��V	� Iݣ��E�~{�Y9?j?{�"���nH��t:���	��={�0.�2n����q�;��L�J�ؑ��2��\)-�ۭ���0�QdY�Ç)$�Ɋ�KE8�2�G���q��Fi�yf����5�:����O?�4�{��w[!^����R�k� .���3�>Al�8��A��bEKKKE�H�_�V�uW�D�q��Fi�yf����%=: `[F"�2~��85z�Ƃ2�0zT�_����ʸ�˸Տk�F�gƭ︕�+���B���c�4z T;��E��/P�e\ƭ��N�h�̸��\z&t@/�$2+H��7n/]��(�H"�ЮY,V,..buuuW�>���(�2.���m[��3��w�R��LꈪOF��!�J�:6�~�b�S���)���n?����q�v5�<3n}�ݭj$t �_U�,��G<��M"""�ZW��`RGTu�(��C>S&�DDDD5��	��������H3�N� &uDU��6_Ǔ�C"""�ZcDB0�#"""""҄	�����Z�p=�|�$����IQcRGTef��	����DDDD�;Lꈪ̔	� ��C """��X� Q�1Y�rn�%H�0zT[�v;���vumkk+�2.�(�Qm�����:�*��}g�=+��BF� ���5zT[Z[[q�ر��J����ʸ�˸�5J��3��w\3��K"���)������ڊ��8��V�'��˸�[y\�4�<3n}�5+&uD|�6:�0zmgƽ���v��_��r�2.�2n�q��h�̸��̸��� 6�L���u��vA�ŧ�!Bſ@6�@v��2.���(�6ό[�qk�:"��3ro]�U��JG�!�"�V+b��2.��X\�4�<3n}ǭL�$B��w'_��f�}g�=0Z͘T�dY�Ç�q�����q�;n-��:"	@�5#1:n�V̖s�.b�Z񈈈�H_L�&�k���j$v-��]VIs�%Q�`RGdJb�rnܥW�}g�=L興���`� jE��q��U��A�M�,��/�P������ͦ(�CG�����7��O����v�e\�58�Qm�����8?jH~Ťn���Q5�2�eɿz~,\���
���C�����
0*�c�K"<g�x����k2��r!\��汶�q�^��#���Q�cRGdb�����uX�c���k��0)*	��^'�� ��p� ٠Q�1�#�������G�f��DDDD��/w�ҽMDDDDDT�d׌�ͤ���i��@DDDDD&$`ʨ�L�J C="""""2��(��ͤ�˙LPF��������C�q-��+u5��X\��ݡ�DDDDDT�2��72>{啡��ũl�x"""""jd2pq�����1�RW����f�""""��&���L��sq,���ֶ��������Y��=��/+�v��|� ������d��$��αfR���q{���L�������|
 ,A
��=�|�����I
    IEND�B`�PK
     �]�[$7h�!  �!  /   images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     �]�[��n GV GV /   images/5a738b76-89aa-4728-b8e5-f09c859dbb14.png�PNG

   IHDR  �  "   �?��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���|w���������j�dɲ,˽�v�$!q��;:� �H.wGr$��B�����s)$�@(C��;.�w˖l�����&�Ųg������gƊ�7kiFZ�|������LB                 d�]                 � �                ��@�                ��                rw                @N �                �	�                9��;                 'p                ��                ��@�                ��                rw                @N �                �	�                9��;                 'pϲ�Sgj�vړ�&���{�����4��oxL���E               ��s9l��n�ץ|�C�M���>'����"�Dc�h`$�a��	!�����"�^՗jz�PUE>�#���B��������7���aI.ۺ����_{���w($               `���/�kz�@5e���nE�/���8�?2�=8����ݎޑ��j�$��&�Mf�-5�j�-֜䲱�/��a�~v�����2��֖=�z�[;���               �Dg4�6��sj�S���ӊT�e_����0�����}ښ���h���T'���	2:�7V��tf��55;y�oWv��\Z�\��P$�W�Ն7�j����               �(�|��Ơ�5�k�2x�Y}=F��Y�E�q��7?ftvqg�6�qD��w+�A�� �~��:��Jo[P��"�r��a��Ը�]���~��~��ں�               �#ľ��\�ϩ���rٲ݅�/�,H��:u���"z~{{*�k�	�;��P���;���u�*��DU[V��i�fm;أ�lث�li�X8&                [�������u�P{�g���<�Cg/�I���~��~���T�j�y܏���]��A+�+e��gɟ0{ZQj|��yzr�A���]j뢫;               2'��҅�R����ݚL
}.]rrcjl�߭G^ح��R,��/���c?mN��&���&;�ۡ�'���e�S�!<��.m��%                ]j�
t��3���5rح�����Ƒ�=��.���}G��A��X-��R���E�J�4����+S�xB�_�ܦM{;               ���4_�9�IgͯI5��j�~�>~�<��Yz��z�]��ϊY���-�++�|B�+9U/�qD��|��t�               8^�]vv�޶`j��P�ש�٬w-��������{�'4�pO2:���y:if��-kjɌ2�j�A���f��               +�ݪ�V��{Ϙ%���*�w��w-Ѕ�g�'^�;:4UM���鲷�$��x�ϲZ,:{AM�����E�oث��~8               ��ȟ^w��z�?�h�}��W�����oT�����)p�_W�.\���A�c��v�,�����ˏ����               �����Gϙ�j���Y�\�Ee��u��g�P|
u��rw�Ӯ�ϛ�s�	�oNm������Γ[��s���              ��9}N�>q�x���q;m��s���\�{�%��T0��M��|�RUӵ�N�M;g��7U$O��               �.�æ��>G�h�1��D߾�,}���䦃��D��b�.Y٨��1Gv�E0���R�w�Y�����Ү#              ��3=X��w/Wu	ͨ��s;tӥK���L_{|��&�Ip�8�q�"�1�ZH�B�K������3;��_lU<�               ��U�uㅋ�vڄ�9gq�+���|A�#��&u��<���_���!��N�}�LU�鮇6h,<y�              �d�Xt�;��ғ�̘Q�׷>v�>���ڸ�S�ͤ�Ϫ.���[�@�KȬSfW��W�����9u�
               ���a�?\�Xg̭2�����?x����+�ū4�Lʀ��͕�ǵK�r0�A�ԗ꟯<]7��s�t@               �<�>��x��TSjd��f��_�D����ׯk��t�3�M�'/Y"��"dW���?_a�ܟ��{              ���(߭/~�Օ�e�H<�Y�<����M�'��&U���%u��ꅲZr?�>4I��;24���{b1�`4�*֙�[{��j���[��-�|��Z���k�y�������v��|�C���)��ߞՖ��              ��e4@��GNUE��\���50����	�ĎF��X<�O$�c�x_"a�U"^�t�J���mV[�Ӯ"��Y��9+�
�~�˪w��z٭V}��W'|�}�܍o�u�/P.f���Q�92���;��p�H�w]{����ښ����v���@��꒼y��y�ֽ����<E��g�              LPF���.?Me�e.:�=j���=0���ѱ_������GN��w?:��?3��:���s��`ae�י[�ݤs���f��?|I9�>)��XT�kϟ�S���]�c{����	=��}׌����Z���so�ۍ��|��*<��U���k���s�Ż�iӝ8Y7~�)�<�'               L%}�ç�T�}$M�~�g���������������|��&�{k�u�:{�՞��|���N�Q^Phɑ �;�h4��ߤ�j��O�S��,V.4-��7��ڲ����_������k��w�'��0N��k+��5O+��rز�U2:��'���<��G              ��W�s�:YU�y�~)�'��m�ݻ;�w`���Z�ӕ��кjU4���[C��?��$�w[Su��r�ש,�py��"1���-��&t�}nm�>yq�����z{�'�?�v(r׃�k��o�<_5���?8�wͫ/~oe�����w�V��{���1               w96����-+���	�_z�ȓG�F�.]�ڏW���\�=��͇/����2zi�5�]���ԙ��գ/��D3a�E>}��S'M�lo���v�����r���qw^��HrqY�uW:7��ܚ��낅�l���߫;޿R��)���              @�1��7^�Hsj�������v�����|���wk�֏_���������O�-��������;_}�|��s��k"���|�C����*�R�-��;^?��mW�~P�[]�oimM|zcՏn]�P������L���J�n�t�n���H      &0z�x�	y�q��	���.krݦ�H���O}�1+����vKBV�  8nƵ�p���蛿n�K�B�aU8&�Ƭ���,�u��"�Ԕ�      �M>k�Κ?-+���m�u�?��?�z��!M0w\s�S�ł�o>�����;Kggg���q?���^w�o���_ń��؛�_�⼌ﻳ4����w�r��VMp���;��������+=�zZK�{�.{FϚ��z����      �ƪ�
�	�b*�Ǖ���Hȗ\7�5{3] 0nF�}4j�pĢ!c�����V����&��     �-+�+���ge|��xB/�hߴ�;|�;��&�֏_�Br�r�=�����냅��ܿ�i���[��~��	k"�p��٬�f�gt��x\vtlڹ��_����jy����o����8�6�Ȣ��zK��`���ơ>���!      �>�5�wLW\~gL���#� �4ޜ}$�R�b���F,�[���7����B�      H���<}�%�p�q�?:8�򮎫?}�E��$s�G/�Akk��u?��)�+/��82v�+���Sk���{fB̨8��g��g4et�:G��Кۯ�������%�%���#7��Ss{�ϙ�����o� ��O�k`L      SY�=�2OTE��J=��2&�� ��+�|�1���Q�z�6��sԦ��z,.      ��鰩�=��se.f�ƴn�����׭��I{�筿�U7}���Λ^��9�%�L���a�թ3�_O�T��0�|�C7�Y�
Dg�˻��ٴ�{�WoXۣ)����u��xlac����L�����k����<�xb<     `�cm�7�
cxbrڸ6 �_�'Te����f�=���sԪ��'���]<"     pܮ8�EӃ�_��h����W�z���q׵�lomMT�}���V�q�2����ok�ƽ]z�`nG�'L���ՋTV��ȾFB�ĺ����_p�����[�-yҔ�y��Us����C��Jt��3��3o     `��Z��'�
�Wzc*t�  N�͒Py���1*����wa��Q�B1��      ����fŌ��o���/�?���׼w������_t�}�����U�)-�8ҽO�բ�/]�������V�������9U�WG�p���G�q�ի�i
{�9���~�w,���㴧���eok�;:t�sP      ��E	���ɋhzAT.뤝U ���'�PI�D�7qרU���7��aw     �?����/Z��EV<�Я7|���w���ۮ\��#_����/Ϭ
ҽ��"�.;�E�x|�rU��}.}��y�����#�nm[jt0Rn�|�]�{9�΅5�+�:�:���nM�`\����m�     �Detj7����EU��i�Z  ِz��K�E%!���t`ȡ�a:�     ��+�1W%��'��|�>t��Bʗ�]����jFñm�LK��V�T��lnӖ���E9p��y*�:Ӿ���z{_��?����~�g?��?��x�����O�޴N�<�H$O�G_�-     ����WCA89�r��� @.�*�*o45�	���ƀS#F��     `j�=�H�-�K�~��Q��}��rŚ�
����C��>0#�5z������ܗ�b��^�HW��+E��wO+���t漴?��M{��v�u6ߑ<0�?�k.~*q�#�N�]�|uI^Z�1�=0�
�	      �٬R�7�Ƃ�ʽ���׭�n������~v�M��^O~�� ��y5�����n�XF����y��Z�͋��pԪ}�v��w��     ��բ�]�(zN���p◯��ȧ?zѿ
ԃ�k�J-���'�>}N�)��WMi�.Z1C?xz�rM�܍i�?~�ܴ�g{[oϮ��-��n�K�z�ƛ����3L�T�O_[}�ˮ��6[_y�U     �<G\�
ê/��iͽP�Vw�\�x<�3�n9���p8�a�[,D� '��G"��cccM�����rddD�P�5����j	����mخ�}.�	     `�8Y���
Һ�p4�'_;x��csͻ�9��~����%����Θ�'7P���rI��ߵ�^��i��ގ��W�zg�y����u�%�w?�γW=�������%uz|�^�<�'     �\R슩�V]^$դ!ی�yyy���W�ϧ��2?�g�;��� �{l6[j���?�D"tJ�Ac98����Tg�l2~���ES�g̪��N�t(�\&     `��8�U�Һ�h<�������+�|S8f��>�eǯw,�Q6#]�����Y���G_Q.�ɀ��i��jN�>����zx�>���0.�]�z�힇���%���<��rUט��#oo�?|�Y     d�q�&/���Z�e�u����B��#� ��d L Ƭ!>�/5����>�������7G��z/rǵ�=�E�T����"q��     `�y�iM*���V߸�����+�|F��VK��{<�����<��4]�y��Z=��.�;�;��s2�~�I��d�����/|b��|����r�#��W4|ޚ�)���jnm�6��     @v$T�iAј���N����U\T$�ߟ��n�� L>�;�^UU��X,S����z{��ӣ��0>�I^GB�JB�����t     �GQ�[.oH�>~����7]v��q���G
���9�}_]Y�'�0r�F�۾��rE��=N�֞:3m�㉄�m9𩻮�d�pBn�j����w�>�zU��atq���O	      ����/
�ȕ� �ѡ=�����D%�ũn�  LU��Ţ@ 5���Sݾ��ݭ�.���f�ûӖм����°vt     �ĻO�)�Ö����t��qι�	���]t�{�c�z�u��rQ괖jͨة]�}�9p_��A�^g��?���3�\��.�]�oo�=2�:P���skK4��D��u	      ��Q-(	)��L���p���Le��*M�=�.� ��.���_�h��W$QWW��vv�ȑ#�F�i����3#�����~��	     L8�<�޵tz��w��6�m?�VK�ȝ�n�z�:����[:��t�7&~�M���F��[�[�:�����/��8[0M�Uћ����A�gs �mM�>.=���;     H�GL�KC��{���n�A�'GQQQ*�  ��xH���"5b�:;�q�HF��n[\KJ�4� �M=.�r     `"��9�Խ=O���_w�5�S0�'/�����~�����g���)�+UU��C�Cʶ�
��9�Z�����$^|���~xL0�]׭�����.\���t܌]�T���|�     �ٜF'�@HM��,J_V�՚
�WUV�:�j �<��~�#n�ݻ�t���T���s�8�:�|T3G#z�˭�PZz     ��i���e������CO�z���L�vp��꒡���<��V�E�h��ߤl˩��%'7���s�ۿ���Y��^��������JM��g��5���<��      �bUB́��BrX�l���Ju���s�r  ���PYYYYj�B!�wt�P[��ҶϠ'�s�iπC�t��t     ���5*���R��k0�y0�ZH�����}���n�,�}3͔�Y\���j�G#ʦ����RS���´��tp����j�������\v�Ϙ3�U�'^�H(�S�    �ɯ����2� �h�^W���< ��p�\���M���~8xP�JKWw��HCADվ�6v��ƀ㭏     ��է�n"��K��n��F�����ߚ�ȯnX<�l�ٵ]��6�F���[ٔ3��g��x�dyew���iu��\���������]��댹���K�     p��ք�B���"��|>��֦:�ӭ ��RXX���1��Qm�i���3}?.[B'���.?�;=���     䎙�~5&G:���s�-�_�U!�v�=7�}�Q�u��a��tpO��:cNUZj���c�W��!#��=���ʁ���
<f�>oIw     pܪ�ZZ2*���`{iI����U\\,  �ی������L+G�h���4}?AOL�N��^���8��;     ��jH=�&v�PȈ�?z���=��w,�}�ٵ��<�H��Q��D��Ԗ�TK{��#1�=2�>!c�N����ue�6����"Ք��@���    ���&��$��s'��X,*+-UCC����t:  �c�ZUYQ�]��ڹs����L݇͒Ђ�1��E�L�[}a��     +�բ��Ԑz���uw��E[��Y�w�C�_R�9̮}��i��u�����;�^�QȨ[�Xݺ�W��X[��3��i�c�?�m     ��(q�trpT���i5�`{Ey�f̘���< �����X%+V���v�RO��7��ΘΙ6�W�]��g�o��;     ȼ%�A�{���	E���.2�hJ}R�O�_���ڧ�T�?٤��#����=-j(3�n4W[��Ǆ��r��[�e�7�]��9��    �_dUBs���w���577+??_  `�Iݓ���رC�����6��/)S�7��z4%�     2봖�4�~e���_�v�^!�v��?���ݥ�S3�E�nͭ+զ��ʆ��W6W�n��^w�Ν�W^������?y���k���\f֝,PuI�ں�     ��8�:58��˼��~�_���TTT$  0�!��+��ѡ;wjddĴ�ިΫ�sn���:     0Eج�Tf�l�hL����⾫����?z���K̮}jK���/k�^3�Hh�ၿ�f�ZK����W�>�q�p     L�/���Q9��tm��|�5k��e��@  r��bQEE����<�7v�R86���ת�Qm�uhc�K	��     ���i���8L����[��K^��`��U����=NS;��#�}��p�Z��3̿9������/���UG�oG?�q�M�*�$y�����     �o%4�(�yEF�����6�U���jhh��j��  `�0���֪��2r߿��҉K�%V�;��;<��     �ϲ��	+����U_�amO�COn>�)8�̺U�y�,��pϰ2-����� N��������u_��=]syrϒ�3�.�^*�æp$&      ���*��s����>{�ly<  �7�á��ͪ����m����kJݠ'�s������l     H��i��}�{(�ُ��!�u|U
~���f���2ߔ:����KL�i��;�?%䄃�C�,����5]��*�ڼ�[     `j+v�tz���������2{�JJ̿f  &����X�\Ԏ;�DN��/�^��U�Z�����
     S���PC�������Z�	����-��*>S;�ϫ+�z���b�k�~����׼w��⍅��50�����-G�&O�     Lm��:�lD6�	��MKud���
  ����!j�֭���8�zV���lTgL/w�u��     �i���Ե3�	����3v����2�;�̚sk��z���-�7O�<:�_B�h]�*z��x�����̺-5�;     `��kqɘN�Z���ռ�sUTĵ  0~N�S�.T{{��nۦp8|�5��9^{\��*     �	KGC���w]s�z!gt�ޞ\�p/�w�"�S{�2)k���<xM킟z�{$�-!�t��(�05��\�Mg     �"��Ȓ�1�,<��]� �Y***T\\lZ7����|�a��ݫѨ���     ��3�:`z�C]/9�k.~�̧�G��^��u��M��{Cy��5v�|�ڵ{��2*�}�x�6�Մ���R�s������1    ���nM��QUz�'T��vk��*
�1  L]��ͽ��-��=��P�bWL�֯y51�     �zґ���<(�}��{���&3k�'��_�vP����{}:��C[��s���,��3����f֭/��k�Ļ�     ���&��bD�����4w�<9�6�   ����j��q�N����ۍ��a�zC��    ��z�*�w�Zs,U<�!�t��>�\�p/P�e-�>=h�_���'BNj���P^x��5��Ћ;	�    0�����FR]L���bь�566
   �|>�V�X��;vh߾}'T�mK��a�;�U�M      㑎��{�t�^�vH�9�C�{���ƽ1�L��%Y�W�Z/���X��m!'�FO.L�W�|    ����S�v�3~�5�^�.X����_|  S��j���f�~m޲E�h��k����o;�j!�     �ݴ�|�k���*��^{��S�Z�x�f�,-���)9����#k���gj�����;�����##�6�fy�+     0y�9�:�jD>��ۋ-\�P.�K   �PQQ�������>�:vkB�*���G���v�     L0�4d-��"/9�k`��"�0���>���@�2%+W�y.���v���r���^�lJ�6��<(���     �>{Bo;�p��i��2{v�{*  @6��|Z�b�^ݸQ]]]�]�jI���=��U!w     pґ��<#䬁����´���"yM�������Ccto�a�����Ӟ�)�7�Q�2�WV�E�DB     `�p��:�rDy�n7�F���  �
�á�K�h�Νڽg�qױZ�S�G��ݫ�sJ    ��'X�1�^,���J�Y��m��r3k�3)+w���)����;���=8�US�_cV=��"�ۡ�Ѱ     ����uvը
��n7�cK/V   @��X,jjj���Ֆ�[�8�&>6KB�ʇ���^��;     �ӊ�ݦ�����^�vH�Y�c����̬��3?���d�W��az͑Pl����G�{���B���;     ��Ӛ�Y�#�nw�\Z�t����  �ˌ�f<�^y�UE���a�JgT���C^u���     ��<���ݞ�P����:�kx�ʤ��������~!�E"�n�k�Nӫ    �LKu!�Q�����F�}�%r���B  �.%%%:i�2mx�%������a< X5������
     ��۬�������Bnk�1f4f4K:��NV�y�;�+�.!�E�	ӟ�1��"     �yƥ����*uǎk��߯�K����:  �X
�r�
��a�FFF���1Ϊ���ͫ�!w     �?|.�L�8����㻈��i]�*z�+n�ʹ�~Z��FV��!fKX�BNK(nz��ag�M     &��%c�ɋ׶eeeZ�p��V�\  `b�z�Z�|�^X�^����U#�ת�Q��ͫh���     `�r:��X��㻀��EL�;���攕��#���G����z̮�s�    ����֬�8�� �d�r�R!��/�������ө��m�W�      Ғ׍��CB�E�Fw)�Y�2ݐ:;w�CɉDB;��v
9-�v�]�I�    �	�6/�E%cǵ-�v  0�8�N��l�	�ܫ�Q-)ӋG�     ��!�����
�L�g��\V��ۦ�hBѢK�
9-;����&�    `b�;cZQ6z\�������y�� �I��/?�$��a�������̂�zǬzc����     `��X�OY&d�	9/��ͬ��c���J�=3�k&k�6�{�$�zT�Y���욑sl    0Ѹl	�^1*�u����Z0~�/�  d����ҥK�~����侴,���MGG3;u4     �-1s3�)6�
���v�f֋D3�\CV�ј�'��/��f�)w�%     �>F,}epT��������X, �  &=�áeK������踷�*�S�#z�ͧ�(��     0U���g,�6K���\���h���������i)r��j�]3�O�     �3�8�*ot��j�E�Z	h ����r�e���/(
�{{�=���G��C^�<     �T�����n#�>x�vSo���a�?'+����ob�%q��T�iv�������     H�i���������j��Ų۳r)   k��AF'�֯W$��%�����-     0����z�_b�Y�BNkmMX��ͦv<e6������#㿑��8�r!�9l��F�?�     �����V��&�����\����RK  ��(???5���_T"1��R�&X�cv��      S��u;��尙V�e����	>^a�ԙZs`d�3��,���K���BN��8�̮�74&     �ی�+�F崍/�e��Ra.����  `j+**�ܹs��k���+JG��P�F"�6�     �є���cZ=��H�i6K�4�k�d�!uV���K�������L�O$4���3     ��Z!�{c���b��B\~�_   ����448�={��{[�-����z�ͣ��    0���L��^w�u��U��BN�l+̮�?�G�GM�Y�uLrZ�ߛgf���1��㟊     dN�;�y�����بʊ
  �̚5K���:r�踷��j	����%     0ut����Ҽ�BN�Mz�Yr�9!'�sͮy�oD����{W�����V�:D�zB��Խ�o(�:Mm	��;,     ���քN	�ʪ�=�^YY���z  ���?�^X�^���x�}Į�M     `jHG��fM�.�9���nv͎�)p7�nI��"�i5K�ߍֻ�k�z퐐s���f����     �gAQH���������ܹse����<  ��a�۵x�"=�쳊D"���x�pEpL?=���    05t���v�˵T�Y��R�kf�)uV��=C��mV�������9'�k��5���    �\U⎩�?����Z�p�lV�   �y<͛7O�����%��ΘZ�!m�u	     L~����Z�9��{VQY��Ys`$������;QY���ВASk�;/��TU����{:�     r�ՒЊ�QY4��U��٩�   �˂ee���վ}�ƽ�ܢ����	     Ln{�����V��&�����M勴�XCW�Mn&���n���8a�~�"!�|��_�u�����=2      �{��U���̚�UUU	   �nVS����ԛ�a�H+����6��     L^G�GRݷ���jx��h��$WrJi��<�kN������l����'��x�sW��3��?�q�M�::�����i3     ��	8c��k����nn   ��j�j�z�g��o��wLM����9     &�D�ͦ�sk��S\��_�sNU����{�f�!u����'K(��a�ԇ�d-�#rYr��B�()�\bv͝�{O�o�s     �~K�B�����n���ϛ�Z  `�<nw�a�M��6�m���Ю���     ��v���p�(�rʧ�y���4�cv]��ɴ�ܣ����:sO���C"��S����Cl�.    ��R�Q��6������   �_UU��vv���}\�9�	-(������     9d�]r��5gV��o���i_��BN�{=�X-Sk��� 2-kw���ݦ�[j�[Z��ӂ����|?|������5%�?�%y�     ��a�$��$4�m~��O   N\������Q(4��d���w�;dެ�      �l�o~Sa�æ
��3��˄��P^x��5��V��'o6MV��R��8-������O
YWQ���f�4N�m{     r��@X>{��?�f�j������E  `�r:���Ң�_ye\��Ɩ���gm޷�     &�ޡ�u��8�Ժ�kD�='����S�
ͮ�y��G���7�9�p4.��jj��҂���{ֵ�[gov�-2����     ��#�f��:�655���
   �	��������qmW�iz^D{��     ��K���p�Q^���o<|��\���U%�����X�7�(�p7���vjic�Ժ��*[�����+/�)d�}���/+1}>�Y:Y     ���hL�q�/���Wmm�   `���fuvu)_����!�v(���;     �ы;�h�I���4��E�O'W����5am�^��u��C��ޯl�j����GL�;lV���O��.dMS��o�Qw�.�     �BgLu��O͙3G��    ��r���Q۶m�vƬ<3"��Ow     &��{�*��aGעc��>x��_y��7����U��;��f�5R�	eC���l;���3Of��\�Pv�w?:�+W_xPȸ��{�YՁ"��v��C}     �aAQH㹬SSS���/   �O]m�>�����S�[֮��tq    `�����#Z�Taj�B��Z]�wOru��sj��IG�g_oW�d=�~�oD��z�<��,��e�����&W�2�����t����CY{     ��bWL��b���N�C3  ��k�=[�=��㸯����hk/]�    ��~����wâ���Z�~ ���CBF}��Gn��̮;�j��)p7�fK��w���w������7��KȘ[�}�Җ��`:j���&     �����=��TӬYr:	K  dBaa����t�m|�VZ�T�P�.�     L6Ͼ~X�h\N��Ժ%����Zr�2!��Ԕܘ���ooO+ْw�+�U�'����
�NkMy���w	�\U�5������{���P�     @���c��F���}>_*`  �̙9s���+Ǭ;ք�
�z��%     0�]�_�Ѯ�Z̿g�xF��Z����ׯ�2���������t���k�mH��΁Qmx�C'�,7��ɳ+�k��ѕ�W^���v��2����od�/��8f�     i4'��7Ϛ�t<  �?��ri���ڵk׸���k[�S���     �l�xi_ZGI�����*!�Z�~ oYc����=8��ugSN�?ٰ/-w�æ�?H�N����<P����5�c�~��    ��+p�U�;���EEE*++   2�~�t<xP�б?�htq�Q��~�     ���Ү�:�7���kz핳*��������/���VŁ��*޴\�1�0r�ٔ3wcʃ��Q�xL�=�����o?��[/_}��6��Oण����     d_�?�c��itmojj   ��n����A۶m�v́�v8gv]     &�x"�'^ާ�5����Ms���_r�TH�۾���+�+�LG�����>e[�܍��c���#g�������[������k{�Oܬ�Y~Z��?�����     ���U�9��7:��~   {j�MӾ}�422r����qMK���?���F      �߰W�9�IN���ڳk�J�����r��� �ESM��v�w��^oWG�_CJ��	�~�����&y�濬��1�6�lr�Y0U��~Z����H:~�v�զ��     �7�0,���?FC�   �]V�UӧO�֭[ǵݜ@X���v�:     �z�B����$ga��TU��yf�vWie!��tD�!�lc����}��w��x�À�H��L0>��AY"!$��rZI�����U�uuO�TW�U�V������SM����ݳ�����y���ޏ7���)�������憛��+�i(��?���F���7��,Z��
��%����}xӅ�1>_z�ة����>��?z��@ƺ1�W���;�����Uk�a!�B!�B�:V���>�����!����B!��<�6n�޽{�J����17p,ٜ�#B!�B!��V6�u�m��4���]��r���o�s�c{��r�!|��o���]�ڬ���$�?�V���V����ۆp(@X ^}֖�&����x�[R7���?{�i�w7������!�B!�BV�-�YDTS��;v�B!�����[��SOz܎�,�B!�BHr��<~��!\�{cS��Xo�ቅ�����G�����O�Z$�<��_~�$Z����N�����+.<�)�k��v��������WN���Ǯ��+/?c�����'���9!�B!�B�ǎތ���}}��!�Bi6oތ��?�LF��nKW���"�7�͍B!�B!+�W�.ݵ�)-����O~�����ǿ��={Lu�������4�5�80�{�=�V���_��Sxݹ[mҧ6u�/<e��w����y��}I���S/9cӏ:�����/���!�B!�BV������!}����A!�BZMӰu�<��ҏQۺ�xj�i�)!�B!�BV�bN�^qFsZ�E�k������w�/����Ajb��[�:s����OZ�K�=�V�%�s)�t�^���On�k��y`d!�}l���={yw��#�ݲ�=4� ���8���B!�BH+pro6�U��靝�!�Bi=�����a��c;{2xj:��ŝB!�Bi7����q����My~����gm�6��7���\yH ���?���]�/h�k<��8z~�DK�-�v�Sx�ٛ1�k�k��st{&wۯ�×�H���n�8sS��-#��|�ʯ�>B!�B!��<�b⤞���Vh�B!��&�Hc��8|Dއ��8�l�ݗ	!�B!��r�\���~�wi�J���a���m��r����o�D����͟�|�Ʒ4�5���A�Ѳ�d&W����7���׹��u���~�����=�'V���뻞>}��P3_G��i��~B!�B!��;s��r�횪b� �B!�˖-[�-N��2�N!�B!��)_���x�Y�1��Rꡞ���]n�?�p����'@<�䗾��ל������;�}���x��,Z���[���~���m8}�@S_�glz�5߼������u�:H��M#/����i����Z߹{/�o�?,�B!�B�Zek�|{����A!�BZ���~���bffF�1�:��W�Z�!�B!��^,���¿?�?�yM}��C]�W���a�s�zͧ?��A�|��?��Ugn~��67�>��ƿ��I�"-p7L���|�W"R��Z/ߵ�������_w�K���I����u��~�I#m��n�k�N�+?�s!�B!��V!��X�)��e�fB!���gs����G�>?��X��P���EB!�B!���m��+�܄�w�6�u��;�o8�O#�~����o�7�
��_t�8s㛚��nq��l"�V�����s��O�_qZ�_��#'E��w����Co?��y�����-?]��Y�����=�d&B!�B!��VS����t������韏'�B!`���x�q�!�����B!�B!��?|�!|��F,�5�u�:����;�ڵ������s س�T���ދN]w�r��=���9�VeU(P_��i\|�zl�m�k��28��>�^���~��o��0����>|��G�[��ȏx�={�B!�Bi�t�}Æ �B!��P(���Q>rD�1~�B7�� F!�B!�����T���(>��g5��:�!�?^��:���W�?��+��Q�?��f���M'���;O۴nx9^o.�-R�2�"������õ�{"��g�7�D�����C_��������Xc�sϗc�2v��wm�l9nq`qxr���# �B!�BH�QM�������@!�BV�������9�_�B!�B!����y��Ņ��k�k�4�={��<6��C�|�=��k��_{ӻ.ݵ��=�e�t���a|&�VfU�-���u�X�
9sY^/֔ן�������k{n�e���7��ϯ��������z��5u��'�uiyÜB!�B!�gCG��g߇����@!�BV�5\4E:��~��.�wB!�B!��1M�o�� ����@��x?�����w<���������:���1վ�?��36�)�6����-���9�Vg��-�w�^��u��޸l�y�6u���M��ػ���Ц�����g�l��y;���#Z��JZ\x��$!��V��YLwT��vɏ;�*4�D<\�p�,zw�)D��;#�J~��B�z~/��Rƨ�H���J���
���T~�0̧��q"k"�3A!��6t���_B!���P�p�}��I?fCg��DE�B!�Bi_f|������D��^�z�7^����n}��ǒ��7x�a�)����{ֶ_]����|��������Up�>�Ė�l]��q��u�����������ؾ�o�����m�_\��w�����z;����O�|���@!�ԋL�pzwDAGȺ#���j ��)4E�f�����0��>��f����T�@)\���+ӥ��Y瓕W�R}�4����gߕ��fB����
�k��f,>G8����P!��B�Aՠ����o��5dMYCA*��uV@>mb6�ͤudx3B!��P�W5�;�.TU���(!�B��c��u��Q��@L�DJ!�BH;�)
zb
b!a� +� �Z�f� +�X��eW��g@-�^�뭔����gК3ET-q�j�P��3U~�0����P�-�l~�[�2Yʳ���n(Hdd�ߚU�5�2���x"!���<��8�t�c�ϯٽl���߃/>m�٧oJ���9����=��6��|wө��/8uݙ���]�H�s��7�Ar��VU�����Z?��s9:c�{���[Gw�������ѭ����g���Ǳ����ι;7u�#�,������} �B����J_\�`\A_�j&:4QE�j�Fz�L
�\�T� �(�%�_����f�5���tyV
����Z��i,/����� �(Ў����k-KJq�t�W��mk��\����f��������3��o.>W؄2��H!,�E�0�H!�15$ti]�t
�H���A7����B!��P�@D�3�
�:��B!�����G4E:��~̆��Bi)�2��}q�!a�k��������/�Ӻer.�_z.�l��2��`)���7"Y|��Oh)f����A0]��y+5z�&
6�U�ee�#f�T�0�P�P�e9���"gj�ME&��TNE"�gML%ML&�	B�Z盿|�n�%�/�|��b������F�֏^���|⪷܈U�;�|9v���/:u�]}�Qˌu������9�V��h��?q�}��;^V���r����37�fvg��o���}'����\�V{��݋���?���3#��g����~�TF�V�B�M11��o
�"@WHGT�A320s��z:��aŐz��������Ei�ƪ�����=��1.�܎�Uӂ9ט�C��ޝ�v�q�}�q���o����X~�o��m�jB�U�E�D�����2f9�'�7���A!��V6tȷ7����B!��^���q��A��;�<2!�BH3��������S�1�X1EG9(��z�t�t
��%_1��Z*���j���*K�*�n����|y(�k�p�$
��sn�Y�y=��L*Yy�Y슏���ͣ-?p�,d��,ܽ1��B�
�`���-op.�ê7���7H!��v��o݇��/-ݗ�S7��o���;&a��y�[���=�������go~�X_Gd�����1����&Ve����g����>x�9+��=���/K�s{�~��w:>��O��O�����7�~���:���!u�? R&������&�A!�=�*��c5���3�bj!33���I"�J��SjQ\RX�P��uk�D��t���qI(�;�����\y�q\>�8���w� �`��8�;+� �^5���t2��2�(?�
Z��b��n�X�_�B�!��0�u�I�Ь��d��E�Bi;�u�ܭ��	!�BV5���cVa����r~!�BV7a�q��x'���3d��a�*�JCϦ�XX(��+P�-Y��;7g�
1���
���Y����qŜ`M�B,ۚ�o�Q�U�o���\�l�2o�5:�uX�`���c&"=D���ݢu-V§�׌�i��M�ӑ�=H!�+�i_���1�ױ"��b���]����O�����˛�-̇>s������9g���c+z���b����j��}��o���:�!�]/Νf<��柏�=2�oG&�?�>�Sh>z��F;��r�H�[G{zW����о������B�������jAp�	�Ur����$���ֺ�Y����%��P��s��֪�ν[���<��׸�h�b�c��`�m�)\��c�\�����¼�h%r7���������x��Z%�kC�D�+�H�j8��ł��������!!��DTQ����tw#��B!��^���
͜�e�����p'�B����`c���.�/b n��s:�T*U8OɪPf�����~"�c�2,�W(
��=��.�
�ʔb��nEYw}v-�r�ߝk�ݢ���ߙ�q(��!���=@4G$ڑ�MFN� i�0��pl������ҢL̥��ޅ�/��;^��������_v�=�ؾ�><�����+�`����8{պ�����ypg̺ Za�Y,_��ꀻ�o{�
������a5���uh8��>���S~�����N���o?��������M'G��{7�t��i�ևC+��2F�b�o�}?�z�0!���a'��� �CYD���M!��G:���Q��T�V�-�^��6g��j^6��f�lmw	���cѱ�\ðO�)��X4v���Ea��̱m�j�c�$06���`��^2�!��5_��p,�bߌ��\��B!�1�!{���vB!��Տ�i�����c�c9�_�V#!�B���l��R1ҥ` j�S�6��&��X���Ղ�f�E~�t)�WI�_��/��c�oh�w���Ex�����7t�Wy�h�o(����YR������[�i`g��X<�XgW�>m�0�a"�60�a��BV�����_��杗r�+�XGx������_v�3{�L�<=�������>޹�˱m���h_��N�v�?x�Pkv�������_��W#m�:]��� 	��قV�+V^�s�t�ħ�9�������{hb6}�����?~�l#_��|w�P\������8�}ڦ������]Xװ�t����o�BH�a�O[��Fv}V��������\!Įd�TzYPR-����z��]78�kp;v���u��v�)H��-��Ƞ�3��5�p�{߅��c�@�mξ�ލEa�~O%aZ�������X�@�3R��p'�`<�bߴ���	!��F0�I�k�!�B��gp` X�=N�BY+��	as03G��B&�D*�(�s���R칠�X~�!<J��ʰ||� �X���ߚ,n��hͯKt����c	��*�B�w(�&�f�����Jw��7�#뀡ő4#8��p`���9^�B�r��I|�_�§�y	"��������s]oo~{G��������g_�I�6����'�z�Í|���!r�X�-����_��y�����x$�Z�],���V���"�n]���w(�[%�^�jO_��sy��r�4�����dO̦����s��Sɔ�h��)9�X�B���O�緎X����n�Vԑp8<�ARUm[wG�̮h����躑�x�@W�e>�!�
�]�����{_ !���%���>��N]�,¹$��y$�I@W��C��E��b/m�av�M���ã��)<�hw����cѱ�\-�Xx�Sn�E+T�S�9�@�h���O�����^��Җ�Zߍ9(��P~m0d :/�����S���a6�:?�J!��#�a%5����B!���	��E��5���-��B!�Fƺ5l�Q07Сd��)��g�Ng�.�@BAjџ�t�*/Q�3���R,�P:�� ��k��\?�ЎlIV-�a��X�w�0;$�C7�P7��w�M��k�s�C��;�F:�DS�̘84k@7�BH����?��_���Hk�W�{���vr~hmW���s��ɹ�љD�d:�H:�}.��'̜q"m�Љ��#_��ԟ~��C�Hh$�P6�5e �����l���uD�\p+c�ۭ��DZ�Ъi����ՠ���<��To�hZ+8���o��Ck;Wt��?�(�����}�A���} ���tGU�P1�Y��L�3�@ƀ�U�Q�-
��.8��.��k��#��l�{����kα̱�|��;��	�;�A�,�h�J P��9�81?��OCˏG��CQ�����H��X��ϰɁB��/o�r�V�ݺ~$�B!�����B!�rr�C1Gmc7B!k��'�����) �@ra.�CM�P�
�6O�d�W��~�X���h!�'z���A���q;����z����Z�� �wi߰�M���Kw�N&a&߰'|�1*�:eFp<�s�:����͖BZ�����t������Z�����ߺO�����o����oi�̮����}���-�Jq���>��G������
��d�:>y�����@!����Ul�+�ٻ��������T��U��H$�`��PNAJp\d�m^����~c�9���8�X�6'��WCCа{#��}-c/+ж(J	��ǆ# �����'���0�]0�]��E�xa�-�B�n�$3� �B!큥m���c||\�1��B!-��ʾ�?�>�!�̒����L��;;[����
��ʰD��L9V#|D��לh�7�5�9�?4%<*/��y�h���Q~�W��7\�����x0?71�Y*ǚ΅px����\�ޝ�B����)�ٗ�ħ��b�wEAV���<��}ý��n;Ж�ӗ~�O.�_qB*/<V��d��ƣ�&@!��Xa�S�4�F���H-X�LAM��0{rQD*��W�݂�vAJ2Ю
�-dB�ݽ�d���E�ns�&h��~,+X5#�$��6_��yA��jl?�1�N��\�C4�=��2B��z�'�<;i��\{\�B!�����p'�Bi+�0	�Ũ�B!�D)�>�!j$���A:��:��P�av���(��vg����Z�e���ߜ�Xt�7�܂��n/�z�A|C�p��7���B��r,s�%�p�j{�f9!����Ӹ�ڟ�Sx���?��E����n���V[�-nyp&�R���}):ca�����<>�ջp(�'�R�bb[�қ���Zfr�Ш��)�.����X,^`�
���U�vQ�]-Vy�#N�"P5"��*J'lk�Y��'@�0�;S�V5o�1������d�)�\=�w{K{�p��O����3�����x��R���d�7��򶅄Bڗ��\Hɺ����!�Bi��@�G��B!+�h���*�#���X�����0��.5��b1�B,�2,������9�2�N�	����փ���k���m��G��7t�c�ܯ����P'���xvR����	!�ɱ����_`��_��NY>�<��?~߾�9�mp����cxߵ?���~!��!�¯�>�O�x�YB	��U!f�c~z�n@�ѐ��P� �_��)H�lo�8�'P5F�*|��[Zp��ƕ_���Ae�����).��5gؽ�xI���ī� !�ZĪz+_�E�r������}���`L`(?���DGg�xf���Qx�BB!m�l�������B!��=��]�/TU"��i&R:uB!���U��!��@R0Rs����:�!����߿C�����w�=��z<D���eB(uY[Zw�����*��[a��cY~��Z-��Ҿ�`���aw�oXC)Vi���͟?����9!��r��ځC!<9�C*BY�X����+w�^��w�� �g6��_�p��ڑ��[<1��_{;>��sq�� ������;��o}�pH!D��!l�3Ы$���F*��VhUА(QjQh��{�=�)��%VY4C�*�����$���Ħ��űR��l�9kns���a#L<�Z�2�sf����̥y����岗�jia�Z���֜B�0�.���[6���:��ޠ�ԡ���XP:�oN�S�Y��BY�����ވ\Qoo/!�BH{��*:::��� ������ɶ�	!��eeK�{��P
Jf��@F�2�")�ó�OT�%Q�%p���7t�#Z��+|��;ז\��R�X��+�2�:#�U%Y���X���p,(�rY��+t���~���"��^�U�oX*�͏Ǻ���>��.Le#xvJ��&�	!k�0q��?��L�CW��X�EI�������_��T�ʚP�����7��=goƟ����C�`��$����o^!�o6�j8u�D��Bva�D
ꔊ�b(=��"�@��0����#<5��=P��x��/�
�b]fw�P��zU�]�IKU�AEH]�KM���y�LM���e�tQ��ۃ�n�w�9���iz�a��5�\3Zj�K�T�}�|�X�:�o��)���F]��v��}Hk�8��c9d�cBYt�h�ܹ=�� �B!�GoOO��{�wB!�^,q�@�}UKC/x��;</�w�H��;��C�����_�ݹf?.�����[���K�*�����EEY�	;uW�;b�",ۼ�,{�+� �;�P�+�j�w(��b���+�y�s��ǻ��B�{?���U��x�4!d-��Gb�|�m�c��>��a�e~��{�ٜ\i�jeM�M�>�O�������o���B�DSLl�^�J��	d3Yh�V�]+�H�XLf����#N���P\p��u�r�(�s�y�u��5{�])����|�u׹��ŧ�Ƭ�">G�n.-���Ax����ι��{�~I��U	Y�q=A�~P���ǂ�{�897�?��P~���^�H���1ު�BHk�ѥ����!�Bi?���G�H��5A!�y4E����!�g'��d�N��@���9�٥�C�^���z��^/����v���/>��_��/�U�<��}-e��|F�c��8�.�z�a�k���B���/��E>a�k��l�o'G��CR���!<5�C�y��Ҏ���U����T��?�Z�>!�15��gnz �<sk�5p���м������N��_~
�!�Z2R��B����� �����0N���e�ca���mZ��*p)��l���R2A�z�,*�C�Ő�G�� P�C�g-�����B����&?9.�����#�k�9��!�5�6�7����5W��e�|�
�/>�,b-�ŮF�1x�=� !��c���N�Ø�-�/�����
�`�\O�@gk!���/"��`]?1�N!�Ҟt����!IB!d-b�b�:��]f��	d
�Xb���=B�A|��5�[�z�c�B,�",_ѧ0��R,�1��Eٵ�ؽ=��Zʱ����{e��7�n�	]�l~a��z<CO�P�7��m������I��Bx츎���;!�����'�������`�0�\�{��õ�<����)�^sw��n��?4�x��􊳱k� �k�
!��1ءb׈��P
����$0a5��д�a�*��)L9ũ �� A��*{ �z�,49��kp�+��z�}���5�q�׼��������qNuнJԪ8�<_|w��ͪ���U%j���P�[��|������k�42ip�
�/�Ǝ��H�rΥ������ul��XON���D�B�J�%p�F��k�0!�BH����l����	!��Z�ܫ���bC{bz��eR��/��������n�bE^��G���>�Ǹ�3��W{��u�|C[Hݻ��x�9���P�	z�y{�e߯xP9��/N��Aw���
��л�Oq��������+4%���ݠ�0�xu�Wh5�?~���&�����{>�3���O��]v
B* e9<�����C�	�5�d��ľ�������ڀ���K0���γ��q�S�ˆB�*��;���6ųP3Ә���:c�]`�U`w�KRA��T^�v�|Yh�X�Mh���"��x��J��s��c����W�U� 8^���V�9���A�KbW�\Y|*	Q�/�9��*�+��� �h+=�Q�hd4��%\U�6�D�������9��\�50��QL!dy�
ɽ�ttPC!�BiW"�4U�n�]FT��e�ӄB�.*v�J�&�L$�Ni�R,U����=DE�����
������%�rNX�e�+��j�����Bqٕ3�.w\9W9_�&>�6�����
�� Ǖk���⋉}B�\E���:K��J��B�~�w����X˰ܼ���Fb���x��^!!�m�du|��O�����j.۽ĝt���o�|߸�idrk�}`M�-�����g��헝��\�Ѱ�ĉ�$�������_��"�����C!�ܫ#n�bnjX�_D$�"R�%�^�ك�"��C���dE*�P;��$C�KBՒ�T����}�k�^t���׸�c���s�GD+� �����|I4�r�
��E�ҾB���_�D����{U��?�^�`U�pe�D"�s���\٩���u\5�52�\�/΅�رt��1!������w'�B!m���utvbnnN�1�!��5B!k��
�2�����R,)U[,Ŋ�U��l����7��s+����v��l>�T!�(��]�%���z��Kߓ�� �Nm�X����q����U����p���R,Q��'t��Ω�����%zy���d%���Ӱ�B]#�0"}8��c9dX�NY�<1����{�ғ��������%����<| _��1��Ma-���%��w�/��8n�ճ��ғ���@���ff!��|7��ܚ�!dmb������vf��sЭ[jZ��H*��f�%�^�HU!N���Łw��Q�&
�/���Seؽx�x��<�s�sn�n������Տ3�.��jw�,q��z�+ /ދD��^�w���w�<6cQd�	��d��^�Uզ�Us��<��Y���6��Ąى��I�BH#�1M.�g��B!�����$�n}Pr*B!���ҧ��!]�,�'af�&5V)V4Z� 5M�˯K&�^O9V��Q���5T̋����?(�Ek��Z����)�p1VsB�2�X~Y�X�`՜�V�%��
�aw/�P�����	��2t��GCW� �n<vB����	!��{�9���=�Kw�ǻ^����������y����'�ܑiܫ�Idp��?��޽o�d'^w�VtD�֏i|6���z߿�y�2LB��*�U0�. 1}zRG:�n�+lX��$��JcUN�r���<Ghw�{�ճ��778ϩ^�>��w#��n؛j=�9_ٞP��fV�S9�
�{�Tr�����K��xe��o����F����RM�.BVb�"�1\1�5<�t�ON���D�BH�X��^����	!�Bښx<���0��!��V����rK���40�!���B�$�B%��������p{ �j�sNT�%������j����2�~��>�������潎k�y��by����/(S���\
��۳��X�oX�u��)(�N7u���j� �'��͑��4'��"����!���a���M�򒓱m�5�����;�?�o��4��Ybm%�`��?��G�՟=��>�x�v��V֧>n��s��#�3��u��Z�1���~��榧�N�A����T�]��D��F5�WRj��f�|D)���6.��T�0�S����v��Z��=W�f��������߽,��.f�"R�߽�~�l�]J�4��5��]���C�K��QY��t�B��˿ot��[#!�BY��@c'�Bڄ���������G&�.����q�7��^�P����;��}=CQ�]^�	�׶�����m.��r��)��+}��W�5�`�h�~�����=C�B,�&.�*yx��XA��A�n���;�e�0&��_;�;ABV'V��և�㶇���x��;q�����n�YHeq˃���ñ�H5��0��M��_>��|g�4\�_|�z������H��'�rxp�qBH;V��ׅ�)�@f�2�4�I)u񶁚V)Jل(-�H4�.'J	��a�B����E*g(�)L��J㒈�?W�&�w�����YrN��݃��e�dB��q���h�t��D,	���Ʌ�����+��%
��r�����>}#8�w��:2�B�&����b �B!�K<��^\��@!d���Wîa]��&��(H�E/0s	��q��F�ܫ�C�2,A����h��ʗ`y���(ƪ���y���y!�8Y_0����݂���{�Y��d��
C��z��B7�0�_�V��8g�	:j�NЄ�Չ�W�}�+l��37��݊���)^z��4~p����#���@�a�]�B�
�[�`w��ސ�6b���U�)�l���p?� �~�(��BښH����6w���9��BɤVhi�B9%Jl��Tv����Cx�;o��T�t��m��I�W�L�c�9�9��ZƵ�:��F!#f��ڝǵ�+*��{�л��%��HUja���D,�<o�ۛnw[��Z�EA���5=��(.� �7c�����̦i:B�&�ʷnZ%�B!�K$��^�wB!�E1�k$���Y��H&�	IMC$���P����B�OP�K�K���b=�X�>�!��(f_�p{=~bа{#B�~�bP�Pf/xt�op���b�*��:6�������wQ	�K�]�͕��=|Ɔ.��A<3��v'��>�&��/?{_��)��s��׵ʩ;��/��|�?z��ٵ�D������Kᦻ����8.>m=���:k�0b���B�?{�<s�<}i��	!�K,��v���EHN���#�ZlY��
�va����.ѼPk���ցN1�~�ڃꮡv�M��&H��굼�n�ZE�Z�%�n�OȒ�d����㠂�нz�v��W����ұ|нV���X�]E+]tl'f&5�񲘁��$"���0��[�B)�T�B�Њ]B!���!�:?�R_ ���h��3�4l�B�'
��t���bq�",��k�ӳ�]���-����b-��⠻��Y�b��
��6*��H�,H�=h�=�_�<�u,�����B����y�~�X�A���v/o�*�������tF�6��v�Ơ���(9�� ��!d��������G[�{*��1�����v�a��������80�{�)~���	�u2>��w����C*vo�[��{� N�4�xde~�V���}xt�	<��	<wd�p!E!�J<��uj!Ԟ�<c�(�,X�O8�nZp��۽B��!w[��j��&Q�]u����X�Z�*[��B�[��*H��Ya�Z��+���c	 �N�=侜��hι&'\Ʌ��,�ycQ��WF�q���.b�,GkC��z	ZU��v�%�^�怹��ѵ�v蘂�s:!��]��ܕ��	!�Bڟp8��(�	!�� �b⌱0�u���G*�F:]y�g��������9���"��j��ay{�~>��S���m܌@����M�e��A�B�|3��Z��Aw�?(�����r,g��t_Zw����g��j��
�-;q#��7��ƑL�=�C��]%��0ٜ���:R�,6uᬓ��{s1��R�w+���)<���x?�%���b��y����f�����y��F{�}]_a�~�c}�0|#H���Z��sx��la�>�qxr���tET�t��e�'�YB�Z(�HIp���{�۽�)�US��.Fم(�XdW=Z��T��TK�]r��]�w,s\�+.���J�p{�d���������A�P|���f�Es�8�^)f�D,�he~{#�Sв�9T�5�R�{���oC�Gнj\�l�&���g�:.�2��P?8�`|�awBYk�49�"0�D!�BV���Ȇ�bZQoqQ�!��e�j��G&�F**x�V���;��A��@ޡ_)� ��ӳ�����z��Av� {-�ߜ�8�Zй���IhY�����?��fz�A�B��{�r,Q�������s�a--�n�a���ŽU"�m�x�`�R�������BZ�'�����P8�a�X/N�oV^���Zy���Ɣ7Y��'f�8<1��[��<���N#��'��M���\
��쑃�y�w�;���8z:��?<t���G���R���h�,�Kf
�LV�\*�م4fL��Ǧ�1!��%,Q���al�/6�O����HYd*�QU��8e��ك
U"TU��.<�ϭ��	O� ��ze��W��"�>�Z-c�qa�� �=�V��pCZ��E�r�G.��+X���_<�tY3������U�w��X�����97{˻g�]$^��*E���g�]6��K.�Cї���B���P��4��B�Z@�u3�wB!������"�������U��BȊ`��箏`sləcГ:ҙP�g����ޡ�Xk!V�R,a��Q����^[1��g�,�o�����m��V<^T��b�]���kz.�x_�����;�ޘr,�gh���6��ݱVtX���:�n=�������8>�?הӏ	!d%��K���=V1��0�ׁ��z:"�툢+F<Z�PwD��Lgr��F��`>��L"S���&��Mb|&Y�������o}���!�����A~ƘVhZ��Cv!�d�x�@�d��L�P�W��k*TI��]D)�0�� UZ�Zs�������mέm�w^�V���F@��{��%p��=�ͪ)����Jv/���W�w7��&b�ir�γ�W�M����SsЌi\���ً����Bڙ����6OB!���X�}�w��ƀ;!���eǠ�����Ez>�D���b�@�X��w([���.��]K��a��yR>����oݯK����	�{�؋�U��^�Ң���z�9�{�������������
»y����B/O�o�o�+�9�?ق,�]�EEY%�*�����@�9���+���zh���(��so�"�;��x�h6��-�aB� ����㳅���HBiY,Q��~��1$���
���
U�*�2�^��`�\�\�,����
�����(���9�X��{��[���B,r���y	\vAH0/z.�����լ����K��W!`���M�}�F�@[����0;��^ӧ"�?Z�-�d�S�"���BU�4U����B!kK��VP�x�H!��la�@Zb���'��v�?��;t�E�`M�v��t��+Ū�+x�=Hx���{��8)7�5�&��s~�2jG������J����)Ò���A<C�sd�����s��dU������b�*�0X�]f=P9�c��8�����c1(��xx"��r �B��BZ�����I����r�!�(%���{	UKk�bT�%�;ŨF��D)�F	R5ڋ�c��TS��-��p_\��d�[!�����ye)�M�����B���p��"��9�V�W4�L�*	J� ���aq���
�;[ݭ�u[®\o�C���<=N�B�U��G	t"�B!���w�LB!AY׭�Q��)�MO�C�T�%��[���!�B�Qx�+����<���X��s����K'+������^>���c|���as�kz>��'�?��ceʰ�ޠ�M�kI��^k�
���2����X
�W��;A��>�X΂�z��@~��>��?f� N6r8k}7�C�暴c�:!��F;!��'�7�pc��,f'�C�P�)����@�� Uoc�S�*�-1Gu�+�[
���T�[�����%H��~Ⓦ UK���@�St	N"��)z�͋ϭ�V�v�"����y�g{�Z"1Kz�[~�w���~���
Y�Zjog��+���K{�hUo�]Z�ͅ���HO�V=��ū���H�^��Z�$/�4�	!�B�A��4u�il�BZ�Ψ��֫�3�0;=LhHi��x�=J��Qޡ�oh��˱ľa3J�*���{��Z�Uw�����e�+��LY��9N��k������f�Esr�aP�Х$�����c-�_((�ҍ0��4��~�����6�	���&�Y���B�wB!+Ʈ�N�M#3}���(�
)QȽѡ�ʦ�@{EÂH�rIբT��
V�-j�)D��Pu��+�6��$�rZE��KdQʿ6��$��� K�xQ0�3��<�	�;���,���}��Jf,�� ތ��E�kȽ ^�x��~�m��wWUs�������!3{q��rԮ!dU!۸�ɓB!��N7�C�z�B���O�I!9yƔ��J��Y�;���EX���7���C�2ޡA�E�Y2k��A��~��<���9)���C�-ê�c���0뼴�`�e�J�dʰDs�����ߧϾ��XA���EX�aw�b,{�=h���gX����Uw���FD��+zT��G�b��濏���BY)p'�����T�t=Н=���Y�&�����ea�qJV�Z�J"�(��#R	D���vQ3�E�P{�w�qq��x�%@9%/�IF|�<%���3���&�M�*=����K�x�s+E��H#�;C�N��X(f	ּ�+���w���л�^!8�����"�3�^KSC�s�x^bv
�	�a8�{O���d�BZM2��0�N!��&zݧ1�N!�Fƺ5�7�#�p�DɩP�ۋD"�eXn>b�@����+PS{�R�꠻ES����.ǁ
��u?�P6�n���3��F��~�[_�=XQ���Y����Uޠ���A�t��g��Xr��`A� a��V���-��K��Ɖ����pź.�Cxp\���BHp'��t4����������Q(S*ҋ�v��v{Ƚ$>9(/A�O���D*qۂ]���WTn���U�
ԮP<p�&��Ϛ����4",=L�Y�Z	x��s����b���ʊ^�w����,vy�.������Dw7˹oD��y,v�U���W5��45�v݅c����<�����ԇ�� ~u��B�f7!��*��9��!�BY��0K�$�Bd����ׇ�>\��I9��?�
�{b�|���K���:�����9����W��Ƌǵ�k�m/U:
pn�*dh�W����~�l��z����}+�r����cA�}��cy���=�V�*��t�~�g���+�
��B�@�m��p�)vcB��wB!McK��s����Cv!�D�jZ���+�)�`{��5,D�%1�[���d���E3�����`,j�M"��Kp�
��E!E�Z�����J��Ur�v��T�O��	Ż�S���b��Jl�
���i��6J�jdؽR�2<����%�Z�rXU��R[C#�e��zy!�L@���e�
:6��Ssx�X�BZ���h?���	!�BH����i'�"ÎA/��!7s��,��?\�`���U���;~��/��}��ڽB����縟+��y����}�{z�~�wн��ޡLA��?�r��.7*�^�7�˫�=�.��Z���tw��3��xU��h�������	!��À;!������1y�z���>{�(ғE�)j�-8)Q��!Hɶ���U� ��(U�*Ũ�}��$
���-�p/��s��*��� ���,��x�9���V����7��ڊ��U)B��Ĭ�k�V!�6����pwWT^!�+W
X>�U��/��K�r�V��P(T�&�bC~��B��]������
��2 S�i0�N!��&z�g0�N!ąΨ�K6(�L�ca~��P�۳�څ�v�b�Z�����^�%�!z��[�K2��^j/?s��������~^XU����eY2���<:��,�f`�PQ|��`>aб�_������VwY��t��V~�3��;����#ؤ�p��>L���&�Y�΄B*a��BHC��p�:��1�����h4Z�dC�v�I&�.��C�Ά��H����dw��6��Ū�|\�/ι�P�S�Av?A�/�.+5>�n��~��H���D���J?/w�M,���.�|��c}�����`,�7�s�$�.+X��J⑟��r/W�-�.hk(�[ZdCg��!^Y����.�V��c31<=��B�JbH�]�|E!�B�pיG!��`�@gd��>}*��B4��{�ڝ��A<Ċ5E�������;<;<�z��V���;����<(7_�-��`������]��ׇd'`�<O� ��tԋ=��\鑐��ʌ�����C�>~aɇ�)Ʋ���	�;ׄ�"�Pv/̇�J&�����u�	!�T��;!���Q����&���T����m�@�W�H������r�}�i�l��}��XtA�p{�gԘ�{a_<�
�{�M�(�,'<y�N�b�L������g�������[X�o��d�Y�\�������)rn�V����A�u����/`���e��)`�ޥ�*A����](^-�4l�sص����~�~)jW����������wB!�����o�@�>��BH{	naT����r[{4�*�
z�g��vg���7��ٽ��ܘb,�F�K���t�]�#V���U̕G.�kb�I&�����Z�e<?ْ,�c-ޡ[����U���w�7X���.w��pWUk_�_�����rн��|����
��tq-D��B��	!��/���Lt��#�0�D*�H$�f�im�	�ˉS���8�liث������W��!��av7�?�4�^k�}����$h��� 'A~���k�BU�yq�J�r
W�9W�'�^��p��w668E,���]��hxw�ݗ����{�!w{��+�^��Vwun����_���G�&��N!�v�� �	!�B�F@�L7V��F!��l���,����L�-��J�d�����|C�B,�b,wqJ�dC�>~bc}�ʵ�^��kʲ���V�������0|��skg��;tΕ~�}B,O9V#
���� �a��ݯ˴a��	Z�'|h�_��0B=���x�~!!��Qp'�"ͩ�!��I`~��)Gۂ�0�Ӹ\�r�P��
B�b��0U�(T���B�W��O���{�O�
�7ShZK"V#~��� B� ��P������A���fq�K�r�J{��{i_o�]�� ��\���{i�5��U���л]�
��-���8:^�m�3}��p&�kh�:!�T�K���ks!�B����}��N!kMQp�z�p���G��,���X��/t�e<C��h���m�b�P.�^z���b�b�+����y���%Z,��׎c�ʲd6b0x ^�#,�U��nw����"�z�����z����*��z=C�b,��
�!w���.�"�0=y��^�m��~ܵ?��W!d���;!�O,a��M�kS���@bJC8^�B���v7�JV��;C��R��`Ws�P��],JY42��/��E�T�|�������yy��]�r�H��Ĥ��~%:y����	�~�Z��	Z�߃k�C��}Ѐ�ۚ��%���W��+��.�� -�^��-�[rv
��q\����QܾHf�\BH3�%/	ҙ!�BH��	x�g��:!��֠'���M
"s��^H#��J���J�Dޠl��������ڽ}Cg���ؖ(�jH����{�^�E�<�V�W�Z�[�%�Z~�_�c��;\���	������?εJP�����R�%*�r��aw�B,/�01;�}���߄�ᎃ*�S�	!��a��B��NK�ڠ�3u��$��@�x����R2��^b�(��lmwګ��m�BTu���M���Jc�x<؎j��[p�MA�4Bj�����f|����e����z���{#Rq��x1�n�<��X<�tN-���w���p�lg0�D�JQʴ	V�	W^awQ��K�*�4d-S=�"^ѫ ڿ�>��Y6BH#��;�M��B!m���n��=i�wBiw��p�`ɉ���	]��˔b����fw��v�v��>{o�V���!����j;.IΉ�ۋFy]+�����ѥY+Q�����]|��kP9�^�U�K�K�z��=Cw����S�U�ݟ����^lu�'������t{OdA!�=a��BH�{5�;�Cf� �)YK���7&�nkd(�P�x�J��	����)�@�ŉ�����
Q�"���P�h�h�g5H�NПaPA��f��i��l�T���:�,�Ɔ�~��Z�+籼xe���X�r���~��2�Uy��\���a�D�q�a<���o�0�N!� �˽�gp'�Bi{��`!���@g�"!��-g�aG|s�Ǒ����9�w�G���J��C�2���$ˢV?ѾV�Ń&{�K�ιz����w���֊�؈_g�!�Fd�[�U�O�<��8X9V����q�й.�	�<Cw�P�˫���@{����#ؑߟ�m��~�u �����[Bi'p'�R� Lu�c��Q�'�BS8$L�����.X{�&:��^"�P����nXO��|^qЀ`{�k���r��k>V[��Z�,���(QJ��j�=�%������/�Q,jW��]��ڣZ�
"\��5�	W^��"�J,bم+�`��p
���Sˍc��^L����}:�4�	!�fd7�����!�Bi?��t��u^BH�)�x����1$��Ȅ�D�
�/�`)~�a0�P��"��X�+Z��Z�ܝ�J)V+z}����K��khdAV�ʱd�K&��5WU�UK�=�W(�s[��	��CgA�o9�O1V-���f�������	\����QܾH�0$����wBYÄU��-��Ǳ07W�*n#(�B�����[\�م��]��R�	��V�y�~���fo���V�Z�ZF���<��8%�J����!��_���aq�+f��n���ܗD��vww��?��'^�-2�v_�$X9���|&�@$�<^?A�s=n?,���!�%����=#�!�BH{��]�Ò�BZ��.��0fB�֑����54���>>�"nk�mm��-��S+^�UK�}%K�����F�Y�s=��Fd5�����y��� ���2��2Aw���Wh˄�E>ae�U���Fc���z���G�/�=*��q��0��1�N!��	!d�Q���
"s���J#�����b��@Z\�%��u;A�G������	��	V���@��
�W�_��_���;̾��+!,�F1KD�d��d����{��{Q�Z
��ķ;�ޥE����	�{�ޅ���@�@��VÂ{.�i����>\�	�6o�]G#8:��B�� ��T:̀;!�BH�J���wBY��:��y�OEn�n�~�X2�v��v7�P����u�g�Zi\�+�1�.p�d�K�X��:�٭DA�j,�*=u=��Z��^kK^a����+�����X��a1���8��B&.޾O����BBY�0�N!k����7���x��b�bh�'��lnw�j��o#轷Q��9�^�p��
���'o!j9���
E��(`-_c���ts{���_�h����m
{{��K�j|�=�he�t��e@�+E,?�JZ�r��C�!w�}�4��8��4];�၉�0�!�o���L&���!�BiO��{A`��BV/g�aG|s�Ǒ���D����vY�P����n��o��b,���Zq�R�:���h��Z)Q���Y��ˍ���3�n���+%j��Q�dz���qgq��m�_�5]⿪��E_�=���.}Ӟ�N���b7q;v��E��$J	�  ���3�w�ޙ;��|���w@B0x�����x�}��p�
����u���w�=�KU�e����Aw�kKs�`��3WO���靻� `�@�  � ���S۴�x�����^�B�B�h P�	�+ũB�+0�����ٝ�!bQ���i�Vq�&q�a}|�Z�EL~N�Ǐ��%N�	��BV�<c�Ƕ�͏)����ʦ��Y�]&`���>�J�lo/��uZ�����*��]"^9���=�Ӥg����G����  @E���kx     ���Ɔ��Zw  &
�}�B��P��W���]l�;>a�P7�^�x�A����]��^�{�}G�#����;J�Ϊ�w^ܹi�sTH�$�FA��r��y6˱��^�{��.�����W����0�f1�q�����ame��4����ct��_ߪ��g|� ����;  �0=P�'��h}�.mV��QQ��"�B�
����xT��@�	�A��e(H�P~1�}<H|�܍;6���sl�Թ���-jP^���63�|�:���Z7��=_o�(b��v����c�'`��������V1�t��:�TA�����umu��7�ӣ�;�կft  ?�u����     #M�Z5or-	  `p�
9z�b��n�Qm�J[�"�۷��;�l/��}C��!�S���
ǈd��y�}Pb�9q�%u��?�-l�e�>�
���U�.�

���B��eeX]ϰ3Y�������+@�n��mA��n�KtB��w�Y���:j,�_�;D˥����&�w  @FA�  F�''��pw)An\(��%�L�
�z��^�]ּ o[��l�-��t)1���ڶ�U�*��$�eߛM�I����{�#L�OK�
%��;��K�_	�{�js��U���A���UAw1�n;��R� �J��pU]���%��ţ4G'�׷Z�2��  i­�;�w�<��.��    `��6��7
   �,����D��Y�Zڢ�bg�g�;�B�wh^�lW��lhO��ݽ�=�Οݿ����@�(b��a�?��ų�U��c�r,��s�����>�J�B�����V�(�6���|C�,x�ۛ������S�i����M�$�  s �  #�g&�4��V+�=K	��)�(ſ�jW�=bT�(�p�	Rq�)�jW6�+�)�Ͼ��c��)ہvS�b��I�L� b%�=�	����ΕD+C��x"V?�8�}��]lfh��;�����y��{��agG������}�R���R�f[�����p%��=o��N����si�t�~9��� {��;��9:X
�!�    0�l��Tom&T�L  Y��x��?�CͥjVv}���p7-���ll�)Ʋ���Gt���V��B�l<�HR�Y�?�0de���8�+t��
��,�.���q3�p�������+��,�b,��
dpw�� -�c�_�h�>�T��GDG��+w��$   � w  ����}�<b�N��$Ԯ���BC�+P��RњLE*&H����P{2:���40�{�$�ϙMQJ�|Q�)ռ�Ĭ8�w�u���kOؽ���лJ������PO�r�)7���k	WRъ�gv�!wӀ�+\5D�J"Z:�������h���;  �;��q����:    F���u��6�u$  �����/�ݡ��m/�8!�����o�K��b��G��IR؍|D������!�R��b���h�g���rAV�>a�83������{��.�<Ü���<C��s����,KA��b,~�i�y�Z��b�r,a%�F�&}i��Ν���.��&� `� �  C�l[�ե�l�6.��S|?A��
S}��8N7�.����1�n��bwǑ�C���~���Yl`Ⱥp5��J���lSa��YI��b�L��!��,E[C_�]|����֠�����6=�U���������įEA�E��?�.�����\E�  ��|����~m_[[��G�     -VWW���9��gh  ��`��5Y[-Ri��܃B�E���b��,��<Ġ�{X�]�Cdb�����
��B)
��0�m�{QH�{TAVZ>�jlt����~W��� ��	�߀v�=�3�����,����
�?�.�e�Xn��q1�`C�w(	�oVnї�s4vAw  4� �l��}�~qJ�u�'L��Rg\�$F����ıLX�J�R����C�s/@��7,"О��$��a��&�sE8KR�
�o*h���6�/�Un3�j���A%\Q��՝k(^�	W�vwؽ���=�*�mj���f@�]�����;┧�]����n���g�Sm����5�[ ��und��]]E�    `Y3����  `�����e��v��r`���]/�./���,�����2�I>ԎR,s�8GÔ���8A��d�
���M�B=+AG��ߣ{_�������7�r�������лS�%�|�����/��[zk�6=w�h��Yzu�D�U�  �6� ����ǖh�l[<�T�r�z���=H����D�(B�
Q}�f�=\�JW�t�=�8�:O�3.6�l�Ra�~�)h�mZ�2N��%��vw����$\��X�����n�Q���Ղ�/��C�`o�B�,X5i��w�Vw퀻0�#`����;ݨ�)�q��sAw ��byK?��b|     Á�u��V�   ������M�Z���b��>�����C���a�3Tb�<Ĩ�Xq������XL�3Ho�X{��*kY�V����y�6���vUa�n�>��*t�_P���wz��a1V�k�����B�����fe���G4v���e�����
  �� ���](����2m��e�TX[�l)�>q�n�SrA*<�֬����Ѹ�F�=�@{RB� ��������MB��=o��-A+����qQ�v����b�]G�����L�R���;����~�muϻ���"^�P�����b�]lg(�o���wό�Jy�~y�ul���  �K���U�    F�L���n4giw  H1ؾ�ۋ]_PY��hm��kb��bp�ݼ�]+��ON�}Reyuy����3��Q)��K�X��1��V���0긨^a��Ӽ/�+V�]�o��v}��r,y!V�#l�o*=�N�{��|��fw�Pluw���G�Aw  H�  �|�t�ۿD�K�,��UAv�8%�Kĩ>a*X�R�R�!w�O����v�P�y˂���AV�c�̉3/�s��`C|R��(v�4[L�'x������&��A|,_�]%bQ�x%�u+w[z�U�x��:"UG�r�+���ٗntW��VY�]�׷��\���=@�3���z��L��%  �Z#O[��¯8���    ��`�u�ǟ�M0Y  @<���:m-�h�U�v��vo�]]�^���y�q�CYѕ�Ku_r����c=ԎR,���:���H� K��Q<Bռ$|B��$�����m�m���{��>a�z!Q�_���/K�da�v�V�����\��Y:��x��+A���MY�}�hl�<��N��6�4  $�  �A<^�����Ze�j�Bp�]jkj�������(F���U�������(��R&����Qm`�!%)2���e��B���
S:�+N�d�=��%����M���c�"U.@���u�^SC�/��ks���
��l��v[޻��Fw�pp�w����{k��ڢ��}��Q�n��7��	  F������ǯ���~��     �����x��,���  Is����]ܡ�e��X	����(��x�����աv��vm�Ђ����cj�Z�=�0�^-�&��fEYq�I�c��m�QO%��>~�_(����2�0(�.�Uc��ݒ��*��G��W��5��A���[���9;w�^�U��-� �6� @�8{�H_<�IՅi�-�\.�E)� l
����L�*x�{�)aJ&>	U���P��A��m�M���%Zŝ������_��T�9l�S&��ld�#`������9��+�64�
V���������/`��{��v;�O�r�"t�uĪ�L�R��1��:�/ыW�k��9� ���V�N��[�Tp    !���Ưn�Z��	  @B�
9z�R���ߡz�������a���j�P��n\�m��Hw~Rb���}�=Zw�bٛcs~���"q�(�4
�P�|\���0�.)����ð2,=��-Ē����^QV��]��+�W�n��M��d>�t����4�ߢ�.����m5��k  $�  �����g���봱��ry�`��h]�k\(�ۃB�wF*N�UM�J�e!�����(��I�Yx����!aJ���V\1+�U��(a��e$^���)(����V�:��kto�m���U[��os���*���sE�B��'�VW�\�B�]y���~��8�x  Y��p �*    �Q�?�/6���?   �S���K:�5K[K��[,��ؘ�7T4�������C�2,U1�Vȝ���w�h�a�P{Z�XIy��X��%�/��%�����b� +��Xi��g�J ����J�r�}�]�:�_(�{�BwL_��t��7�CW~�d5+3��cT������z7���  �@�  ȁ��p�uy�,'�K�RIj�5-D	�w��6�{*'
N*�*L����a N�>���G9Ԟ��{�96�y�Q#�sd*��=FR�j���{����zawy�O�2��U�}=�*���e{"�(\y���f�^����.���{a_���ͽ�	�_nT��W���4��$  V���"@���     `��V����e4g~w  �I.�K�_*��wis�F�B;��������?���ڃ��@��j�&�X^?д����s���B�&�kc����>�����hz�
��Z��;6ʸ$ʳ��{�a�4jtw�������c�}�p/��4�;�@����ms�	���X���� ��hP~�}��Z(��Wo�[�/�s  �
�  0 Ɗ9�ƥ֝�[����,N��A��_��)�@���֮/L��R�v����~��a��վ0���,d��.�%J�϶8��c[��9_�U��{?A�U�{1����9Ab�L���z�J�����BC���=ls��\K��.�ݫ���'�9���y�ŝ-m`�v �𱺝��f��¯X�_[[�Ç     n*������  `�g��Ra��˫Tw��E*��mm�{��~���ҳ��$�Τ�"ԞU�tl�96�&y����sg� k��c%���vW��x��{.�K�/������r,�ս�6�^������
�
��}y{k�ƫS������Iz�N�   ���;  ��ۺpls��7��r����S��v�h�i^��Q���aJK�j?���)��� C�iVI��3�����9lD}��nf�)N��7�l�IG��.��D��}� �/L��*��\��73��+��R�).C��-G��M���T��b�,��aϭ�Y��x�9:w�~:���^�  �D�i�p��5z�RA�    `Xl]י�����6�  ��O��EZ[Z��R�il���~�|�R�V��.�2.��'C�*�D";�!�#̚?8��Xix{�_�[�e� k�ʱ�'F)�
:v�y��>���zz����W�v��c�W�V����X|�������F�g�Q����2�x���v�>Z@�  L@�  R��%zd��//S��XN0D�
���z�#H	+X)���X��.FyC�Ο��*���!M���ci�c2�tl��q�%}�ax\�
P~L~V��β8%?�U�񠰻)�����U�h�
��,�x%of�	W�x�w����6����h��F�{|�U�šѠFe���D������O7� �n���߿��^�B     `x����w�f�ɮ|  �g�P��tz��Ӵ�,Ҿ}�����=�=D_V��,Ԯ
�{���X���ۃ
�\F�?�9&�q�ؘ���F�(Ϗ���Y.���	Uc�P�/쾫�/'�/��>��:~��/��ʱ�ޡw�f�+�Ӥ�|��S���ͦ�g(��*ϰ�p��k��t��@O\=C�U��&  w  H�����ܩ�-�t�)�u!��u�]���_JP�q����	k^�Ѷ��(��*�qQ�G�cs~���
6~���f�T�y����2�nS�ҝ$^��'����zc���,YK�(Z�3���m���� kgؕ�V��{-�Aw�ͽ����ѽ�t�Y�pj��}W/0
  ���&KF[Zc���h�^�r�D     `8�k�zݬM��&��  
�9�����X�A�9*����b1V�՞������d�C�՞�Y��8�;�d���(��γ}�,?^�*��}.���:�H�˶���Wv�^1�*�����%�9��k���b��ap9֮�G����KZݻ�Y|,�
��0�3l4
T]��O���&/����Suk�_k   Ip ��8�?O_;פ���T[�S�����He#���� ۽-���q!Rk;?	*q�dm���ڇ[��;7���$��ɖ����n�=������DmZ��%�J<O�����D+OP='oi��X�&Y�=�c*�����V��v7���,Ch������xI#C��~���N�����S�z�͠� �a�Z�m;�z}˯�tvb�     �p2w����M،  `B!���^����mj,֩P(z}C��XZ�={V}�y�F�=�=D�kk�Z�=p��X(����,Ȋ~O�'���x��7��vw}@�����G�e�a�׽r,�{�O�b7����cyW�nݛ��Q�F��w�*��/n-ޢ�-�Ɓs��7Z�4  H��  �)�^���}k�[�M*�K�0�J�r/f�E*Y�BP�]���\��%N�!	���T�T�%o�5Q*�@{RBԠ����I�J�{������63�|�16L|��%�*�ٿyK�R9�h����d�Tp�]�����+7��ig�6�Wn��7�p��
�����"=�_�g:G?�]��� �c���~o�H���V��?7��;    �3??o4����y4� �6Ϝ+���}�X^��b��ڮ�[�ի={}�0�0Jk;��u
���C���5�P��1I��;'μ��3l���vq���h� +j�=���F��?n�Y����@����u7��0ms��cy}����+@{��n��^����<C�ݽr��t��w� �͟��nah  ���;  X�+��@c�6�6i�X���1�p��P�6*�S=�J-D�B���s�hI��+L���ݯ��D�#P��-@��v�M�'�R�1}�L�$�)��q�)��6�'�1��T���m
Xz�7���N�{N�����	Y&��NWp��"�.S���x�5}��v�����fw^�p�2K�,R��9z��5v  2�ݪA�}~���     ����5�V�Fs�m�W�  ̃'J���eZ[���b����IWyWz�	���P]�%��ʱ��ʱ�	�nw���Ϣ��q�c�g����:� ��sE��ldE��,�������{L����E���\S{�G�zC�U�U+@˂�U�U�a7̮���momё�5z�����1�xAw  pA�  ,p�x��9�LkKTwĩ1O��/P�.��܋eU�=�u���E�\�8r����$�N:�T���a�C� ���FU�r�0�%J��+J�=lޠ�]�
:&{-�'�hi�U758"��L��W��|~�	���W�6����(\�{o�#ri53���Vw7��y?�{n�}�L���7�!Z ���Z�s��X~���S�N     .�ݻg<�N#  q�@��zf�����R��U�a�K����D�����;4^�|~��3�P�p�z�=k��$��(�
f���(�|��P��'4�T���x^�l���}r�WH��2�0(�������\_н}�ݛ�~a�b,�g��1�����ڬ�����eZ��7�  �  ��`9Ozq��뭋ͼ#N�[ڃ���KJ��`%��u�)�@ej�-L��-D��(X�=��L�ƙccn��</6E)���le�1>�F�$�4�+W�j�X���1ꦆ�h�+okjenhP�ܽA�f�ɽ�iro:��w:"Tgi��p����/��U���w�շ��H��x��V9L�Wt ��z�V[�ᒞ�>;;��;    �2{����*,F  �Q�}�j���7����b%��m�OX����J�0�?���j��U~a��H4�����c�u|�9I�c��K��_��|���b9V�^���_��7Z���x���@�{���;{�;J�p�skR���y��W(~�hhc�.}i�5�����ֹv��e  �P�   ��.�p�H����ؠR�$�dK�D)پn�F�=L���S��vY���s�?�����/F%���*��(��γ}�ax̸�lp�����T��gY�
;�䱰��������
L��$�T*�*H�
oh�od���K��+'��iuw���~�{l�r����'���Uk�����H�.T������m5��5	 0Zpp���m��sss���     ����2U�U�9+�y�6�  ��g��Rn�6*Uʳ78���.�Uav{�a��h����p;���kkO�#���2О��wn�eL��,de�'�g���$�%ƙ#�����$~!u����bI�B��u<��{�Q��9i�]������r�G����ϰ��
�-�L�_�?H����u ��G  0�ON����Z[Z��R�ʝ�1�n�����"U�`�q�]7�N*a*,��&�԰�ړ����:���A�7���y������
Z&b�^����Α헷4���Wъ�_�bqjW��.ޏto73t*W��������~���ze��}j?-�'�i�� ǝZ�����������s     ���;w���`/ ��ġ}����O�v�䴶���y�bs���n!خ�!��/���ů�$�Ο��{��a���y<���a2�tl��Q�$q�,>VZ�(��}^�(Ȋb�;6ʸ$ʳlx�6<�x~����G���x�<������{��A��_�#c9^a�7T�bɼC�R,޷��A��8+@�j�0ͮ�3 �-�@ �&G���O/ԩ6�j�BwIA����*W���{�T�68ОD�=�0�� ��=��{�sm�1g:6����:ϰ>>cC��c�s�<~a*h��*��%-P�O��A�_�\�X�\{�+RyD+�pUp���V��<���7;�UG�������p���t�W�m{{��kS������1�Z�h H��Z�����rA�avvw    �!�?�޽w�x���   *r��+9�/MSm)Gc�����m���a_����c
+>Sp�]ԇ���x���H���1�m�1g:6�s�<�����K�=V�aМ8�⠼°�s��e����D��w�#����������0�нt�z���_X��&�f'����,�������A������S�
=3y�~<M�� �G@�  B(�.l�z9O�o�f�A�r9r�=�y���B�^a�_��lW.%nwft�o����6��2Ԟ�`���8s�8G���~��Ay�Ǐ#L��7�d��MbL����9���{����{W`���|�U<�Jv��3������ �J����/����zhg��|�<�d�Hխ�y] d��+)ݬ���z-�J�677i߾}     ��������&��9Z��  �u��X���YڪlR^����~�Prw�A����w�P��o��u���[�O���ˠ�ä���9&�qQ�ǝ��y���Q�Y���s�U�e+�n3Ȯgc���4���M�}�<>�W�������:�.z��q�*Ў7�ms��݃ݍ��+@�+L�k��r �>� @ O�)҃������z�,yZ�*�J#���������.'(��ۥ���B�,�ޙB$]>О05*�TZ���8ӱQ�ۚ�乒$�H�$&ϟ���gN[�2�E�*�M!Jg�nK�?Ԟ�6���{~���ū�>�=�h��ۼ���{W�j�V����:A��"�ݬܡ����9ze�  =��S7�ί�333���     �67[�m�\_/S�/� �hs�X��=�Jk������<ĠP{��(6���u
��Z+>���!���&�����6�$=6����:gV���F�/�S��Q<B�<�X��M�OL��*�1>��/l����X�~��R�+��*�Ck���?t��V���ݝ�i�ѽ�]���t}{��4�ыWO�k����r�  `TA�  $���/6�6?M[�"���)�t��%���b��`$L��������(�+L���IZ�ګ�U㢎�:'�s�����}�	��|�q�)�s����G��&P��M��A�_|?�2�v$Z�[�h���V�foN^&Z9�M�/���	Vݠ����	�V��<v|s�^�z�^���+� �g�V�Z#G�E�뗙[�hrr�y�     ٤V�9��¿�  {�}E��w�h{�:�V�4&x���P�7+�r��!eXւ��v"��:����_��='α4��1g:6����>�0}q|�0t��!n >J�=�Oh2v^a��$�%�z���^<~�?�������{�g��	ۛ�
�'���7�;+C�aX1V�
���{me�>�_��&/�On���k"  �w  ��K
�ؾC��m*����Z��
T�օ��v����ۉT�Tz��dǙ��2���4�7��>G��X\a*���)��I�v�!^����Gb=�Q�xt�V2�J*Z���f'�����۝��f&gS��{D�B����@��
 �0�
3S-ѣG�Zܷ���޽{t��Y     �dzz�X3Z����~� ��xz�H���hs���K��b,�r,���5�����������̘6��I�?L�#L#�>H1���sl�Թ����5,��=�;�G���T�=-�P6��x������sN�VNr'
�y�����'���]������7��cicI�AO�S�ը��wN�۹��Ɲ: �(��;  t�x�@�?�BkKj��K
bT��������v_�n{�J��la*k�����(c���:'�sd�&�%��|��t�a*j��lއ]�����3�d��Oнs�v×"����OW�R��{E�fG�b�jG*\�awU�]��lk��T���_�=@���{hs $��5���3��M�    2
�}��i�� �'�����p��Ţ�;+��.��>�t�g�p�l������(�'��������o����9&�qq�ę�����ϝ�vn�a�96���qQ=G�s�=����_�<��'�3�.z�;;�^��
;�v{;{��^�W���W�չ��ɶ��D}{�h\��ON��f��bm�  `@� ��)剾~�uA�4M��\�8�h`��˖�S*aJr��d���p��?�`� �����G�ccn��6�>Q��q���sD�l��mއY��3�/39�i���rbC�VKC�P����[��{��7;�j�+Q�jݻf�D���ؤ��=49A/��G˛�  ���,��v����^c���iee��9B      [ܙ�u>�����Vp �r�]z�r�VoSm�A�������՞��MJ��}����s�����1I��Y��8nsL�cm̳5?+�����":ϕ�c����E���f�+;�T��̶_���������n�]r�ݕ��M�B�
�j��=G�K(��f�D+�
*�r�k�s�܁<m��@?��t<T  fp �i��(҃�9ڨT)/��K6�|�T�����ڷ���r�{=��*�qQ�ǝ��y��qu�+B����&�t�4ĩ��Q��Q�����_O��of����0�����w�7�s�}g'/���uG��,A(��ogP	V�h���%Z�8G?��$  �͵�2}�Ħ���7n�g�z�     @v�Ͻ�����fkE�6�  �ΕcE�ܑeZ]�Юo�gU1�y�=x�gY1VP�=�`��g��fq�cIε=�d���8sl�M�\�H���ԏ��͏�-����&x79����U�}��tw���D�Aw�Wt����ao�gO9�b�g�b,Y9V��=.ޠ��x��^;NS�X 0� � ؓ�_�?=�M����-[R0��ݸyA��^��t�T�T�@E�P�T��g����S!V16��4��Y��?�q�c�̱9?��f��?_����cfE����+d�-P�O+��?f{��w�� չ�tW	U����������u�n�{�#`���M-�JK�r� l�-/]��_>N�[9F7� Z �1�V���o�^w��߻w�֫U:x�     �lp��]����L�_v �Qf_���/�+ש��o{�
�P��=ĶW������v�R,�@{r�v�R,��A����8�;&�qQ�ǝg�Y|����ʰ���+�G6�v�]w��8����q��(s��e�)d5hw���{P9V�_���՟���>����h����ʱ6�W顝%���Ezi:G۰ C� �=�W.���-ڬ4�\.K�%!�.��6/t�TS���V�ݽO��~A*���x�L�Fw^��C߇-�I���`�}�8e2vU�q��������L���`Et������ɖl6s]!Klgh��bU�+^��Un�])Z��,Z���c�%z���������k' `��n���TKt�P]k<�f^�~�>��     _�]��2����ѝ� ����E:Ӝ���&�d������r��J����3�{��X:�a�`�^s�K�|�4�øs��dL�c���=?�sQ�(�d�c�3�G��g�+��m{��1I{�6��/�?�[���۞a/��{����O�d5]����궹oVnѷO��͝3��]�� �� �=������-L�N�D山^�=D�
�K����v�0�,0�.�ڥ"?v��Y��$X�8ns�ɸ��α9P�N
��s������{n��T�<�Av�qY������NQ�'t��	U�6��������.���Tb��ʠ�İ;�o,N�__<Bo�=�% V��N݀;3;;K�>H���     ������ϛZ+�Eӕ   ����vn��秩Q*yW|ho�/��-���p{X�]�?�`{V��$C�i��Mƙ��2>�3,�DT�O���h�A�����)��
�Ρ{~�c��#��B�O(�$����w�_�:��7����W}�ns�׷��Tc��v��ϭ2�m�  � �_�\�#�[T]l��ؾ�P�I��^����=�}Ad�m]�X�=������x:�m�1g:6�x[s�<�^����%L��f�=� �\�U��$�(�9&��j�AwjU�	�{����wX��_��	U͐Fw_�]�a�X�'Z	b�����6�����z|�"��u�:4+ @�6
��]�#��x~�q�=���     �����sZ�|铕 ���%:�}�6��`{�/,x�a��'���
�=�|���	���^)��H�P{�`�0�����8�l�9�d���8sl�O������%$��:�~7�����
Î�y,K>�lp�]~Wݩ?���ʱ�<�|~����|�X�����.msWc�x�^8Z���E��-�"  � F����:�-�'�A����Z�����8%�%N!���l�9&�6�ٚ���4Q�([�Tй��G��ƚ�O:c!`%9�fx]��Aw���n#�6~��d�UO�R�34���P�#V����B�����'V��Uo��Wf�g҇[���y�� ���r��pJ/���ܺEW�\A�;    � �w����ϛY/R��'  ���ӟ�ߦ�b�gE1V����՞mc)�C�`�M/p��C�c�u���I��I|?q�>L�o��'jx=h~o�f�]5����iK�/T��k-辻���c�x��'�����������kc����׍z��}B/>x�^���4c �� ���im��Pme�/�^*�7/����@�Rk;��T���ܳl�05�U�uǘ�3g���i�o�򜘊da��D�]5/n�]66�U�qSQ)�����s���"�x,�����KE�]uC�i;�Y�{�O�R53���f���%ݷ77�rs���H�u#O�&^; �\_-�Ƿ�@Q����?���z�     @�8�c�|i��e �Q��ã�ڨ4W|.u���u������b,R��͂�=?�I����f�#̊?��7���hc���o����u����u��Q�ŨAv��$�D[~`ǲ���[�S�C�{�A�X�_h��V|�hs-ƒ��|��4O�*��������  �w ��q�`��rj�����r��Pa�f�v_�}��$���߹7�`�����*X%1.����l�#��e�8B��-Q*�|I�m�u�R����%D��?��;u�
AwͰ�_�R����z��f�fG�
hs���V*�J<.63x� ���Y�Eߝ8H�O�{sX� `F�Ռ>^��<��=��{tee��9B      ]xE���u�y�6���Y   vN�����h�2G�A+>_�����&����!��T��s��ilf�p=�Ax��c���57�s�:�ϕ�5�6?)��d� �°�I�_��o:6�ߚ�C�y
��!���{��Ϣ���V�����g��9^_P��S���=��B�ց�)z�����w�i��6w @�@� 02�r����"\���ݶ8l/4/�	��Ĩ��8�T�°���FU�Jb���8sl�M�Y'��%�Xq����&��l|\!k�*�����kt���t����`�mso
�U���/���Ukk�բ�W��2�����~��	=4y�^���6�  |�R�ǏmQ9�=��G�>�y     ����]�i�Kho ?Nk{�Ֆ��+>b��>����J���Ty�}�����^Ϣh�I��:>�$Α��Q�@��F�1�����A�z�q�@���i��ǒ�U���u���x=D�^g2�H��{�����{�&m���a.��Z��X�����U�����@�,�ʩ��4C @v@� 0L*ЗO���R�i^(�K�p�/�Դ ]RP&P��c���@�+N�.Ȃ�D�Ez2��,	S�"J��l��26����:ϰ<������-aJ5?)q�d�	TA���w�Yн;��B��Q�����n؝H�aX��me��W��@���:�ج��<KJ���}���;g�[��y�V  =�׮��=vt[{���"����ɓ'	     �Í7hkk�x��V�fkho /g�����w��;��*خn���{�^�P�!�����ڳlϚO�5�P��1&�L�Fokn�v�<��d�cD�����mޣx���H�/��h��t��	��P��1��sꕟ�-�'���6��v�{�^�0'������r(�����6�_�;@��& ��A� 0�|�R��nRmu�ۼ���=�
�5/x��~AJ��nE��T�u�tnG!�E,�`���8slηu����fw�r�����l���T�׻m�|+3
y���e�������v~��q��ྦ�X��o�>g�q<�Ƕ_o��ƨ!�$�������� ��(Tⱸ�����W��t��%�w�vQJzw���uA�D�_�r�\�`%�7�FO[�����k�՝�N����Z���v� 0�|�\���ԩ�ӿ���'ND�     ���u�ƍHs�[����  �e���pu��+;��vU1VXV��Ϯ�(��c�o��C�/�"
���٠}&c����۞v,��6�$=��<������������>^T�0hn>�j���3&k^b�~�j�iP=���~���f�]��� ��۾�,���~��3t�c�m�__��.ҫ3(� � C˱�y���Z[�I��.�ۃ�)�8Ծ k^�	TV�)�@E$���.���Y� X�3.�8󢜇C�Z����hyyٹϦ�򶾾N�j����֜muu�9��y���t?��r�����?�9r�y���� ��C������[�>���ǝ1�;v��x��{L]�SA�M��6��q�.P����l���Αl�].d���9�N�-��ngP�Y2�*H��uD+1�rw�)�*q|�r�������q�YA3  �Z#O�����5��^�z�     @�|���/Y���]��� ��!z��R�����+>����
/Qj�c���J��H�?0�/؞�'8J�a�sm�1g:6�sm���A�gdo�7���,�u��X��9~x�Z!�6s��������5�=?>��5�~��{~|���q�x?o&D	Ǉ=�Iy��yI�ޓ
��O�K�9ǆ��/4kt繒����B�~0�Cnr�����{�TM�~��љV����N��'��On���� � @� 0�<{�Dg�����߼�ڮng�I��jkl�
��\�"
n]@�=[��a��-Z���?�q(j~~���t�������h�c�J���b��I�j���l[��|a���k��O�<I<��x�ۣG���Ç�[�?~�Μ9����Iq�)��&��l|\!+m�*��cqC�I��M���wG�L��i-C(��BU�~�p%�r���&��z��5B�+�ڣ 	������5z��J�^�L�s!w @0��9y�N���u�'׮��Ąc�    �d`�lnn.�ܷ+c4X  �i{����X�x�~�н���A�=��:�v�j����
��be1�n��tx=Ip�=�(���3=��������'�X�",��7q�f߳�b,?��s~�,���㍿f=�-�r�𼟏�/Ȟ!�[=�$o�#�g;Ȯ;�tL��z��4��c6�B�s�����=��z�F��{���H����/krov
���
�P,�<CeI�F1o��{���e��;Oo��	  �w �P������˻�Y�F;��q�]-VS�`�\��.h7/P�0.J��T̰�^�j�}����(����>n?���ݻw��u6�x���ܹC�o�v�t��
��ysŹ������Z�b֩S��ĉt��9�k�8 �x��&b�ߓ�L�B�
;�V�]gNRb���t���[�`E�̠
����knmq��2�*ߚ���['���U�e�w�������������Յ#toAw ���f���R�O�"]�5��ߧ�=�     �4[�!�z+
��ݩ  ����<}��6�n�NQ���a�������Cu�����څ-�lwoU���ۓ�	��?�{�$Ǚ��3Gg>kK\ru��}gs��n����~|�o]_���x����0 >_����£� /k�w��~�R,wc?�����<�cϐ=B�UAx� |�P5��WL;��o��%��m��6��݃猪��"4�����c�՟E߰�*���&��V�ů����'/�K�y�n  �� ���S���pq�6kT*��"T_�=��]���Z��
T���ym��T�
���FI�ʒ`e��1&㢎W��d��:��YT���u��u떳���
^�n[|Pc<��r��N ��ٳ��,p�>�d�I�SA�GM�29�t��t��{w�lBU�Gw����+q_�~�h%ib�u6�5���]���V������x����  r>X*��G��l���4�޿O�[�     �.�>��666"���v��B  ��wȅ7*����|Cي�E�+�_�Y�+�7�y�ʍ��~/�~�=Ͱ� �☍�cLƙ��2>l���ݻ����Oq`����
5|�oYO��h~.9υc����~�;}����-�ŕ�����k��aߋ�8>�jl�qA���9�z�6|D��%���&��=J����y���W������W��w����0����=CI1o[�w�;g��[���H� �w @�)找u��^�F��R�@Լ.P�� QJּ`n���i]t�=���A	V6ǘ�3���͛7���&�y}ff�	�Cp-����xs��@�-,lq�������;}������-qJ6�f�=��v����qC�Q�S��}ϥ�����%��D+�k�h%��>��|�$T���s��󸃫����g�'��hmk�  @d��:���=u|�h�{�Gǟ^it     sVVW���t��sE��� �}�;���D;��i�Y�;�uJ��0�d�goQ��K��s�p;�t?��::�2��k�Y�#�nv���qQǫ氷��u��Cd���|;ݺ��¬�����N�7��;� ��/^tJ���;���{͊|O*��+���h�X�}Ĥ���T�;$�� ����r�w�P��W��Eo��)�6�g�����2�p{s��6���K���.5w��� �d�J �4W���ZY�Ri���.	���T�@%���`�b�i^0
��\���S���+�>(a
�U8qE+^��C�lf��߸q�����M�,NT�U{�7�M�����c��}��%�z��s��Z���Ç�E�8�j�iP]gL�*�x�@�Μ8���I&c�	����"U ��'�$Z��uD���{���`���}��<m������4M���hf  x�p�L����`I��`�z���ߧ��z�     @|�s�;��ܚ���JoΏ  d���3]��3��!����o�g�K���W{v��ڃVy�n��߆�˲}�����9&�qAs��daa��9���E�#�}��<��j5�~����_�i���~��𻸱G�-�&�����8�wcl��I��h3�n:?hLп��"�
�Dҍ��������]�Ք����y�g����!~a���ze����Q���1���$  H
� ��O/h��ڨ�hll,P��o�*g�Y�]'ܮ/R�O,J�}���{��='α4��1'��8����wC켱 �K�n�v횳��)��փ>贼s����rn��\$��{*�ɱ(������ݻGq*���]J%T�[�u��^r�+Zy��v7��mm�\gS53�VA�_���Ls��r�2�4��f @��K�U�G_9S3�7{�.�>s�&Z     ��?��)���'�%Z�.  d��w�@���Q�K�COQ��7�~��.[�9�?���7�����]�f�S�o{N�c6��cc,}��}�7d?����Od����/ߡ����G�&¯ytg�71�~��	��{�P56	?��� ��cI��Q����a�t�t���w�+@�eY2�P|W��εD�x>���m�����Xk��da��|�~6��;  p d�c9�օ-Z[�Ky�T�!U�}Ik{Q*N�/+n�݀��(ۓ����"X���E��=���O>��i�d�D� *�o�����¯����裏:��'''��s�P�8Av�q�,PKb�������E+7�޾���$�_+�VA-��}ϵH>��Ag���%���v3�M���������5�V �63�E�[+�ĸ��_k?v�	'     �h,.-���t��[�ϖ�Tp- �.�����gk�V����w���l�n����S�U�j��������q\w��8����m����|�>�d�������$x{�W�}�k#���X\�u����-���$z�Wv���A��QǦ��}/&���]���
�=oP�t���}��7Ty�&�X|�F�N���������U��>  �� �L���"=R�K���n�B�#T�(P�S������rq�+L�8a*P�"��G��+NeM�ʚ05��U�q�a�C�~��#>qC;�����*D(�)�����
��������#/a����#�<�Z������v�=��x,��eHW�Ϻp��Ztw��=\���+]�*L���$����(R����o}���zf�U�^�_ߪ  0o.�o_�R���%�}���駟}�     ���?�����?,�9!w  �"O�.�d�U����CU�=,��kn/����E[�Y�!�z�n���ݒd���m�xix�Y�m�#�8n�f���\J��?��>��g��� -\/�������_��{�СC��9���X�'B���sd�+��19>�~��9�������o{?��o�s$h��5�N�=�7l6��1�0��u|����]7��)�ꌩ.�џ/���s�ν �-p d�\n��������N��cc}��[�`{Ѹ�=8خӺ�#R�n���ĩ���m�������cq�&9���b�@;���y�ZXX�,�����Y\����l�v<x�>��O;"/Y�B[�Z�#,�6��,����e26�}j�ʹG��ΐ�h���xz�n��+J)����J�
Z�����k�������}�Q��	 {���<}�R�G�l͛��Y�����     �x���$
|���J�   kr���y%�kT/��v�g��y�����`{���������C�:x��Q�'��h�x�q��.{�b��-����$ ����Z�O��\��� �r9���,ǲ�T�]g�m�0�Yۧ�7B+@wW��c��e�a{���.��=�X�m�Awɭ�#�-���۹A�&/�O5��  ₀; `��<P�N��Z�"oj�50�7�X�k^nmW�.�ǂD��%�"����)BJ�JS�JC�2�6D����w�	���`T������_���ǯ�.\�'�x�{�1G���,p��TQ���H3�WԲ)h��'j������T�D+U�]&X�m��}�zD��
�����9�hU[��o�>H��N��"� ����2F�i��g��|Ժn=r�;v�     ��K�w�܉4���^����ٔ   S�<����^���"�Je�gh���}�@uV|nߏ��}DF�CtI��`���zV=�$<D����������o�M�����x ����_��Սxc�5��ɓN{��rQ��Ą��5��g�+;��|R~���A��|d�tw���u�A�#7ݐ;_s���*߰���X^��N�*��X|NW�LӋW��/���udS  �@� 0P�9W�s�[T]mP�\V�S%�@���_��_ZP-N��v�p�,��1*q�w�Ɩ85,��A��GE��߈�e9���G�k���Q�j�
A
�Y����̌����K��0�۹��g��Gy�>����ѣG�sl��ecvOJԲ!heI��2/L�ᱲ`�J�
�\�J��]lr��=��h����s9�h��Y�G�=������^f��z������	�Q~�{����/?����     ë5~��G���\��� �,���"=�y�j+M��Ͼ�,c�P����������C4/��R�=K>a��a�s��a��]�yjj��z�-����� �;g����_w6�_[yh.�b����w�B~�pI�+;���8(�P�?��A��ecڷ�/�;�]�Y�7l��e�X�1o�{^����Y�U]Y�/\�;G�ӛwP� �� ��Pl]�}�*���5j�>$pxAG�
j`��ڋ���`q�+T�
T:Bӻ%�>�8eS8ڋ��Q����9��R����hii�  ���#��#.Y��C�T�O>�Y�>���=ֆ�eS��r,��g\1�dl����<��{�p�RT^�tB�m�J\~P��.6��r����U���U}��x��|� -m ��^�v�H7�Kt�`�h�Ӱ���٧�6z]    �k�篷�~�h0�V����  �B�H��+M�X�I��Rh1�?Ю�zC�E��vY�]�;T����]�9K!�a�	m��Q�i�_'p��]��׿���!�����_�_������C��SO=�ln������s��
Îۘk3���8(o0ʾ�1��n�]~��d+@�J��0�����o�X�m�9o��p�t�q���x�ɭ)�����^/R��^  ~p ��ġ=w|���O��O����eb��l`W��t�T��&�_�bT"Uĩ���6�4ħ����b/���o�;�C��.mllh�Z �`��������~���v||�;޶@v<!���m�Qq�'j��q�V�Vw��{��=��+Z��D+���J����{�t�./����Ã��<� ث�v~��ߠ}��U^"�ͥ��I     r����V3[1G�7�����_( d�+ǋ����QY�R���U�X���xޡx_�z�wt�0����3I{��ld�}�tǈ��/d�������۴�� M��
����+�8Áw^������}��s�z��16��6Ι��dlZ�L�������C�O�l�v�5tV�*���M����7�
�B,�/��;�W��k����r�  �� ���D��7o��z����zbTH�=�}A��.n*QJ���j�YV�	��D����~[cm�:'�9M��-/��r����^�J�B �����=������g�q������-P��hיg�����|[�vq��hŻ5��h��T|�F
�J|<qs��p՞���p���`�]�0���>U��_��／�]ٹN�'/�_C�; {���k�����3��s?�v�i���      �壏>r~)0*�WK4[�E �_�T���7h���ry��3������E���;4)ƒ�7��0�Ŗ/8ja�4���q�iyu�7�|�	������!��=��������1\�Łw�	��C��~��I�L�XV�B��Y
��橂��Vd����5��%��ۥXM�o�b��=�0�R��'��	�K��[�
е�}��N�.^�_͠ ��+ @*�r���s�X�F;Ţ|Y���es{�0�me���┩@����Vf�]�:�>�}Y�?�c�㋋������ij��o~��!F0x���������'N8aw��_����w����ε9'�~A+������}��V�k��n�VwY�=��]&\�Ʒ���҃��w!�����w�h%�U|�W�/ܠ''�G3cT��{ {��e��ޠ��Dk~��û�:� =z�     @�۷o��7"ϯ6r���> �AS�}��.m,\�|���cI��cx���v��E����[^�0x���۞��q�eϐWyf����_w<E @z��I�������6{�����f��}�st���@o(	?�Ʊ�}Ĩ~��ؤ�����
Y���	�-,��{\y�{{�[��in����]�P��ʱ�V�n��txm������S�� �� ��9�?O_?�F�J/�.6��,+(�D!���L�T5/�*y�]�xA�ʊ0�Q�D�����v�_��W�ҁ� �v ��������^z��������/~�Nk�X�~�"�nS���?�A�������J��w�6�!��kg�q���N^����b�ΐ�tﷶ��}���]��XD3 {����ӷ��i�dv�˿��ޢ��%��     {���%z���#�竱����N�  `�L*�s����괶����+���l���|D-�0g��s�� |���n��0����4�s9�� �����������˗�r��|�3N9��Ç�ー���IK�G4	�g1�n�C���A���|�S���
���{�a�����A�>��/�$��f���ţ���1�[o  ��;  Q?U��
w���E�1G��5����m]A�ؿ��Z��k^�ol��S�J�b�D�Q� X���fA�������,� 1����?v���t��!�җ�DO?�4=��s411�kK��������N��q�+bV�B��J)X�uʮy��J�r�,�`��.Ch"X���`��A���K�.�/n"��^b��������s�֧$��^^E�C�l
xV    �=
k�|]'����ݫ  �3�Jt�1C�M�(��M��D1-�P,y��'��D����O�1��9lωsL<η�����\�š���M d��{��g��輿�Oȁw.�z���r%��.i����U�����Mƴoy��;�!���6w�TY�9����6w��Ϯ_蹶�byW�z��6w�_ع_[[�Ϗ��쑋��x�  5� �ϯ橸|�;��@�X^P��=P��1aJո��]����)ه��ĩ,�س"LeQ�⥃9���;��+���.  F���������c�=�S���x�`��?�����ZI�mݳj���V�[�h�\��s>�6��҃�K��UO��r��UN4�$M��z���L��N����Q�z���^an�@�/��SǶ�箬����|�Y)%��;    � ����F�z�o�R�,�*e �A���ҷ�Qc��J�U�����a�������ü� �Pk�gwe�;�9/�F�o{N�1�8���Ρv�>��й �����������իN�;�\��V�v���4�B��6�%9�F�"R��ܥmR~gGZ�Em���^�н���]��t�y��a�X������)���K��T���� ���; �:�r��󛴾x���r�eA�ܮ#P� ����(N�"��q�T�
�*H�b��g)Ğ%aj�v��6g�x���B� {�`�+6��O��Ot��ez��睶��~�����f�=��i�)dE���Pq���ݑ�:��ab���� l�if�������y����w����[<Fwװ�  {�?,�љ�:�����B�Bx�]z��'	    `/���~��T�V��c�W�����#  ����g��h����l�lnW�����=C3�PԹt�C&kޡ�y&���?��q���+��o���y��/~AKKK mfff��������������}��_�'N8c���G4	�:��<՘0��G�dw7YA�x^�����=��)��o���,]�Y���s=���c�ze����	z��AZڈ�b `4A� `��
�ľ9�.mP�<������۽K�T��vUk����S�~�	��]�J3؞��d#����:������4==������ ����wy���t��G��;����äh���ߦp5�}��b��˾���Ű�x$�s���*�.�w+Yؽ��J�ۿN����  {��������OߺX�r~�L���m�����    ���no��&����8K�^��O��X	 0��(���;T[�SylL��cu|R�D�C�Ȅ��M��$�؜g�/�Q�۞�?v��z��W�@;{���nm��r n�u�W�~�嗝�����B,.���W�BgϞ�E�P���bV<��-�i߲7�+��[��O�
}��&m�=�p��/��cuW�_�_C�
����3\Y��[�?:Gܯ  � � ��/���i�n}w��T���=\�R�f������SY
�gI�JJ�����z�~���:������ �˽{��?����p��qG�z��gk||�cC��#j��oK��j�]ܗ�hE�%�^��_���;�]a�#^u�)��W�`�����x	^^~�;��m� 0ڬ7��ʽq�����+��u3���>o>��C    0��縷�{Z�����R�n�� �oN�*S�,�P�j���W���ڶw(jZ:�!pg�x|{)�>(�0���͛7�P�3n�  loo�k���l��OO>�$}��_v�|�;.�@��~�j��$�z���]��+��u�܃�����r�^)V�z�BUΪ/�.��s�6��v�.�L���W��c�g @(Z ��Z�yp��+�(W,�>�+Z�c
T��3�*(����/V�Mq*�`{�ι�B�w����g?sD����#� ��~���o��lG�q�ݟ{�9'�>66�KR���?�j�l��m�V<�=�c\QJ%VqSu�iTb����to��*��!/�U��&�6w�`%�V����3��7˴�2w F�{���8FOߌ4��kלא��I    E�p;�qp��*� ҧ\$��KuZ_��z�2�0�?W{�}T���w(���+>��C&-�0+~b��m�;�o?��cz����7���S�%�  q������{��y{�ᇻ��zQ��#*��8b���d���ή^���;����t�A�0�Py��ks�b���������?n���D��� �X�ѷ��h�2O�R��v}��]>0L�R],�m^�^T�ɒ85������8��+J���?����t��]�� ����B����lǎ������hיc;�v���&ъ���w��E�J&V�53�!��@�W��k��EcP��Ks��3��'��2� u�[,ѱr�.����ǟ|�Ρ�    �_�p�}nn.�y��<�:7�����   ��8���V����w�J�t���������۳��I��Ohc����s�����_v6�� ���|���������裏�/��x�:a���B�~[~���$C��8ct���� �~�f�{P�]'��^��"�j�g�5VP����]�ޅ#����4_�/���A� �+ǋ���UW6����*G�*���*�p��8%knW7/�E*&-1*+BԠE�4���n߾�R?�я�
�  M�������ߝ�ĉ�o|���~�i�=��z��Eݟ�p��P��/+��qE)�X�ii �Vv�  ��IDAT�'��A'��煦v�A�����[U�Ly�&�]�7�D� ���6�����t�M��&w~]{�G    `��ro����lno�����i��p;  ]��(��۴Qkt�C�K�:R�](�����a�ޡ��ݽl�=+a����:G�9����*ϯ��
���� ���/~���q؝�P.��ַ�E�ϟw�������uΑ�����h�Cl��Dާ��뷹������ð�{^�N2X���-��o���nЍ����9x� �Up D��tb�&mmR/�..%hԾ���Tr��w,H����$�a��j�v����g�(��o:�> ��g�L��(�{�5���	 �'>|����(��SA��G�����9�P$@Y������d���쓙��{f��_uWwUuUuuwUWu��y���j��!�]}����imm�C=��~3gΔ��g�}6����v�WN�Q��[�1/�V�뎴H���L�J�msM����|�lAw���!w��9N7�7���q8�bbo=Ο7OփR��_�^�W��g�Q��n�h�`ȝB!%�n�݂��������h���B�əs�v6a��Wc��ڮ��Y�!�������;tr;�+���Wnkoo�ڵk��/�7ޠH):�ۑ��w�u>��Haw�N�0Aڧ��r��~a�s8y�ۡv+��#_h�A=��ܕM�F>a�����/Pk˱��R���m��%�b�P�̙����K�H�wBHN�@��u~�5�����d[�]ZAe��,8����H����E*����^���0%�`͚5RS���D@!^D�n�ڵK�.��wߍ�?g�u�v;v�����\ǝ��sB �C��ҳ!v�wY�R�U�&w���rL)L%<�ĵPF;CR�ʧ�!��L��._�E�v��yS�ĎJ�|%�x��A?���W��"���o]L�-^���?�B!����������V��i�®����
��pN=�{��H��9�b�ǳ�bi}B����������[�ͼC�1/y�v������
=__֭['c�������g�7�|SZn��v�x�8��Sq�i����Z��K~�Ѹ�Aw����b{�F�����{:�.y��8�*���"�����1�R��O�_}M����u�k�h��z��͛�U�AD��R�P�"�X��sg������q�r�n&E)�H�mZA�p�^�ݯ���LE����y\�c���l\�&��[���ó�>���BH)!^�6m�$-��v�$^�q��x%ޓ��H���C���0����z$-R����(�ܵM�JqJy-��������u3q��E+����q��Qx�k"�t����r�m ���q���k@~�عS�0�/}�K|^$�B)D��[o��C�|�;+�Qg!�XL���ûn�DeeeF)��G4�[+�Jl7���;tr��ٱo!����ￏիW�g�AWW!�����J�K�妛n��e�/��^(�n��h�ioPw�Wt�C�v�g��^���/YP\�������E	�I�PO�K�+z�2�s�5����}?��WZơ%̔;!#�	!��1.�ϏnA�#��V0ש�vՔ��Tb[B��o^�
TzA�l�T�H�/L���mq�k"T������矗D�>� �R(ū3f��sϕ�$�����[�r�E��g_/R�1;E�|E,���9 y��)������ٚ�E�!�v��z������p����)3��@���dO8����¤���q ~�?�a>��Ϣ"�E/B!�/���#��E;l���	ack%!�X̟�Q���=Iy��J��}D�p{01n��۳�����u���k̎}߿��>��hhh0ܟB���RΊ+���#���B�N�6M��_h4^���H��=C9���˾��K�ŵO,]�������g�cY��f�ֽFS����n��>��F��a�tl9Hϐ�� �?%�ٱ����;�.o�nO/ZqJ-T�R�q�0e2��@_���y��Av/�Zv��9�)�D��$��;{����%K����]j�=��p�9砦�FڞK��h�T�+'�s����O�H����+��63��W_3iŪt;C6a*�%c��hӢ�0g^jb�;!�J}W�C8n|$�sttvJ�����gQ]UB!����ny��w���#�����`�R,N�DEg�w��f+�2��ޢ�Y���C�z�N��>^�c_+��/\�f^x��]�V�!	!�\ؾ}���u�]8�䓥��)��"�w�������R�՞�>�d��XT~a� K.ǒϧ��c"̞��!wq�<�Ae�ݤK�W�n���s���AB��	!��2;�Q=M��3��Z��,�^X��xZA���D)�"�aa�v�Qn�S�"B�+L8p@jj_�l��$����x-ܴi���~��8��3�`�w�q�v+�s��R���;-Z��k�;�IY� %�*E��$V)���T
V�qy�AI�RW��V�\E,�*�ш�G���� ��!�ͦ�J���c�zuww�7��g>�i�7�B!^c���x�������h��5�턐"��pA�0�Z2��u|�|�����:�vm��o�?,�whe�b���<�Xcv�ke��?��ڟ{�9����B��Z�E�L�<Y��>�l̟?_�^�_h4^�n�y�C�z��U��[�
��wU�{� K��jW���69ܞ����^w�p�Px�Շq���x�abfkBHy;!D�/�u񋂶F��T��ve��,ܮ/N�:���I�Ȑ��o^pJ�*���S�g�І���W_}UZ���Dmm-� -�\��(�����i�o�������k�;p7����/�h?��7��9��s���{�߽���駟��c�9F�D���ژo �h܋�U�������z⧾H%#�U�v�f$���V��,m�f�I낕��u/ϝ�'wՠ/�!�o�T�?�G��?�>00��o���=3f� !�B����mۆ��F[��1���j��Oq�ʠя����J���ۥP{.����XZ�0�;4���7��x�}�V���/K�����S����Ŀoq�nyW��ǭ�v����/nݿ[�]~}t���}������wn��)����#�<�G}�{�t3A�3t.��sxe�Kb.��|�6w�����BEA���n���K�����mۉ��&�U�g�;!e	$�jv=mt��Z��4ܮ����3��J�J�0���*�(��ҋx���b�On
X�8W1�W�<xPjk_�r%v�ܩ�_�[	��p�����Ŀq���n��倷S=�[���������bq7����\uu5z{{]�!@	�ެ��ߖ�;�C
�_x�8�裥m��rٷء�\��C�*D�R�k��3"[3�hqO��SXv�*����t+��u|�B��}��i�;Zp�Qx�s"�w�xH�>lh�B��)���:N���������ı��f^B!�D�ܻ�6���Ֆ������Z��	!Ea�� �c\+��=��v=��4�nnϥ��?����&����� ��B�v��F㍍�����-�Ο,qK���N�����n�	�~�n޿|�n����w����׻��>�m|���,]�_��q�H%Y���l��ʘ�=D���XMl�I�vQr����BEA����,(�����%�Ik�B���Z9��E�z.�ނ��+���%�b,B��	!*��&�!�ѝ)P�uY��n���)N)E*��9O+(���Lҭ���܉u���w�b�˩��q����{R���'�p-PJ!�����N��E�p��K��VD'�q/��>�n��.KG��wY��^_�V�Vs�*S���'���7�j"������ ���u鍃���o�]����ݻ����O}��v!�22����;7ڦ]vGEs{-�n'�8�ѓ�8&�/��*bc�=�f�˞�<����2�C=�{��Nzy�l�����,ϫV��o��Q#�-��7��[�L��Э�������oír&���Xܺ��ſy�f~v�o^~�s����wss��>���8餓p��J�wYK����e_/�ڕcv��Ny��u��D�=�#J>���mj�䰻�_6�0�B��n���}a���_���)�oc1!����'B{�o�QC�J��̈́)u�]_�Jl7��ە��l�
j/hF�BP��S�w/W��E���?��c�裏�A!$;�5tÆx뭷0m�4,^�Xju?�ä�N�Q��[,A��qN�V��XZ�)!PI[ �����Vy
B�9�D����"2�L/�P��ʢ	�+aF̉5b�̹X��!wBʍ�+#^?X%�|�U��xk[^[����'1i�DB!���{�b˖-�)��%���բ��vBH�Ҭ F�w`0�s(�H���ci�C=��)���>n�K-�ng����R�],���!��_��^���ӧ����1u�Ti{�~_.�s�n�ѩ�z>��3�
�_�hqG,]�%����_#�Ψ��,����k6��z�a�������~�;_d"����/�ab�F�5�n$NIc򔂚p�R�?z"U���B�L�����Eq�+�����'��چ[ZZ@!�>�k�0�o��6�u�]8묳p�E��c����)F岯ۡ�B�qC�R^%�䰻|;-`Ɂu�Vm�]&S�J�_B��o�5/doeP���!�q=��`�l��!�����=P��$`���BH|��n�\u�Q�K�B!v"�A�l�jk���ߏ��``��1��9g�hk@ ��s
��gx���{��b,m�ݨ���C����8'���W���b�
�K�dB)�.Y���sN>�d|�k_�g?�Yi[�~_.�k̮0|�=�\�C_�����м��ωE��5K.�X��aΩ�����A��	!�@k��/d,P�"U���`%�����b��0��RP-L�7/���d��8��0%��[�⩧��O<a�T��B������+W�s�����p�gH��v�Q�_H�]9�h冈�����!ټ ��}x8-^%�k"�л:�'XAլ _n���U�N\4o:V5�fEHY!��׷T!�c��§�mhlDGg'>u�񨪪!�B��tuu��M�l�1��xy"�B&��Do�^�B��Z�P�?��B�o(�ە�X����R�2��:���
�g�H$��_~�?�8�y��}	!�������O}J���ϖ�3K5���q���]W{���ͱ���/�z���!���ʠ�O�J�6��U�a{=CB��	�|1,�Bo�ެ�
Zm_P��+��f"�6�nl�N5���n�BS2� F1��Z�^}�U)`���S�"���o��&6l؀�K�b��Ÿ��P[[+m/DP*��\��fc^�����ar+���XFSʘG�p�|;�8Y��.\!C�R/}��p��xf�tP�"���ack%�)�>��&���v���8v�����B!�"L����uz_Η��p�`��vB������)]�m�DEEeN��LQ��]��R���!Z��B����u'�)�X�}�ϫV���C�0L!�8lڴIZ��n�/<���1~�xi[���BƼ�!�)沮��^��M�,����{�/�Τ�+���2f~V��H�����r,��U���;�<���̾��	)ap'd�R��_0�=m�����Ys{N��S�M+�c��B�2��70�nwB�rr/��f#!J=��صk!���x�&���I�Z�`.��L�2Eڞ���˾�KvWLѪPQ����Ou�]��'��A1�,65ԢR洃CC���J��o�.Xi���9y��O@Kx���bkG�Ըr¤!�t.��&�U��ۇ;�8T�?B!��KOO6�����n'M�!�k��V!�8ʌ�A�0� z��JcUh�J���?4���v�3>�5�gx�b��X��>�бl���ק���}�B�;��-�܂%K���3�ĥ�^�#�<R�Vo��1'��vx�Ny��!T���^H��b��p"쎄_9�	�y��k/m�=3������ϰ�_�4�u]�����!!�@D��W�t"�ѕnn7jp�&Pi�T���i�]n��(��v�8�Ǵ�� >9%`�y��c���X�l{�1�Q�H�"��.mmm���{���㬳��7���b�B�]����dv�B���x���*!@�1u�=��!v�d�d�]y>=�*-<i���6�w3���~SK�����?�D�^�44��R^l�@w4�/M�E�������x��������̙3A!���ScS�o�nkk��t��#�w��%<B��3)�#�{��B�F��ٌωu���d�]n�6�Q��p���P]�0Ҽ�|���\�����aThѯ�?��;$�� >��8�S�}'�p���KAw'�󚇘�zbL��^!�Q�P��:M�F��2�.�N�T0=��I�azh����[�������G���!z���"�2����h_�P�S:B��@��T��n�Bf{���v]q�`jA����
�{E��ul�Νx��ǥ?�p�BJ���~�\�O=��$\���O��ҶB���Ɗ!d�-Z�+b9�.�zj�,9�nu�A=�JtO�.T��:��<ON���h4�c�0f�,����!���� ��S�/O�Cm�� �x�x����b�1Ǡ��
�B!�m�[��]��z��뛫��!�8�	�C8|`��`�;4��9�7�˱�c������v�{�nc�q����b&Hh���q�FB�.�5���^5kp���c�8�����^�C��1����Ct"o�g�����z��XI�P���2�ҷ�o�K��u|�t94��ar������i��q_��ҁwBFGM���D��^�BrL+J
T�i����a��H���'�&���T��v�� ���� �����[��_���~�iD"B)M��/J��I'���.�H
�k��*�c^�����ldP"�Q�􃪰��\�E)`)+e���P2�:t�ԏ�D�R�+r��߈Sg���;r'�������:���^���hin�ܹsQWW'}>%�B�">kl����;̾���a^�W�����!�s�Tv5����|Ck3>����d�]Y��m�g��v�o���q�5&�w�Ԑd��\������x�������>K!�9�k��M��y�f�J�-��ŋ�2m��X���9y�Ӟ���ɞab�gy���e�p89�s,vGRK7���-��{���z��k:���j����}�8e��Bϐ����!#��MaR�}�T�B���L*�i�D*+�٧��8Ԯ�X����S�8}\>co�������_O��!��>�p��oH_��Wq�gJ� n���R����e�J-V�S�`�P��)��T�)*Aw���>aʗnf�*V%O�^�Tj��us�LC�-τo�7����jp��~�eO��P�uN���ߏc���ĉA!�"���ۇ?�ȑΈ��Aw�_�#�8�9��5mM	/0�V�ܳ��,{����nm7.Ʋ�ڮ�U�a�7�ԟ�ޡ2��-o�M��+~�<��ݍ'�x�<�����`;!��0�5���7�t�q�s�9��׿�ѣG%�^��Ӟ���i=Cm�]l�%���ɰ��Ǭ�]q6U�]Y����Ҟ���R�]�J�DPs���;O��3$�`����is��l�_پ���njOߖ��Z�*-T�C��"�f7�ZPG��
TJaJ�0��b�M^��l���{�n�:
S�R��Aw��p�����K/��+���jW�3�nv'֍�VP���b�[�5Aw����h�ܓ���zPޞ��K73����Ī��1(�Gښ���XY��C)+�}x�@5�	��I��ϐ��7c�[oa�ԩ8���PSSB!��\:::�`{gg�#������*�چB�$��aa����6�[����o(ƅfTh1��7T������=�S���>v�m����>���﵄Bʋ���q���htA�q��Iۜ��<�����5��P9��3���٢��.{���U3?�!��w�IԞar�h[͛�"�����x�	)s��!kSjo�
T��v=�J�r�ũ���B���^w�;�3�ƍ����kײ��BF�=࣏>¯�k�N"�p�B�ڢ�Aw���v㶈e�xc�F�Y�}+�úR�2"q?���5�,2%S�F�c��2���sM.}�{��n
V4U":Đ;!���C��SzQ��o|���8x� �O����<��� �B��A|�m���8p��#���Snn��֎
B��T�����֌
m�]��}�g+�>�cYmmW��V�C�Bz���c�q�1l_�b|�AǾ<F!�;����%K���c����7��ɓ'K����<������(y�g��q��(�cP�"��2ʠ{�3����B<C�7T������s'c��j�3$ī0�NH���/����m/B��a�"d>�`�H%R�����d&P�S����t*��R��<N˫��*	S������BF.MMM�����c�IA�s�=W2ќ�{I�*�����K:�.�Ti�JZK�R�r�	�ʟ|���ޒntW62 }��H%�M�S�U���	�K�K�� .�5���FO��Rn4��ԮZ|iJ�����Z���{�n)�>{�,���I��	!�R����c{}=����H�]3�Ԡ5~C!N3�ʏ�L�D��+nO��z�XٽCm�];볱g�-�n��g~�ȼ�]��Wnޡ���˗cٲehnn!���šC���O<!�b}����.m�b�]9榇X�u�ϗFlO�) ���Y�&��F�a��U�=�{S������ �тf�ó���� C�x:q��!A?�hN=m���4lm�2���4��`��@e���hzA���4)2��9n�On�Q�
�oذ��?֭[��C!�4پ};~������D+'�����cgh��9�����C��^P�v��Aw�p5��F���L��K	U>y0-bA����)D/��!�]�8{J/��G{/C�~����v� ��/~lcpp��سw/�Ν�Y�f!�e�
B!��җ�w����l���A�o�����+�b���~|aL3z�����:���w(���g}�c���skn���ڠ�@ֱ���R��u�|���\��=��n����ւB��E�E�D��q�%���/�)�n��h��Xщu+���3�%���>C�jʱ�H�w�3L��H=������g�pO�D�7�=ԅ3&ⵎ�h	;�B�wBʌ����A��--Pi�̦L�Sr��f�JG���g���� h廏ǭ]����?��;�B1cǎR����>*��?�|���K���}�Z�{���'�ԍ	�J=���F9设�3Z�t�Hn���r��@����RjX��p�<ak��p���!��p��js{%������}Sa�YD���?DCC���~�GH��	!�R�����)�YU���d�}(~Y�n{>� !��Yc�L�D�R>a�A�ݒw���YU��1��j�BM!V�w�?�`�{�N��<(��)t���B!J����t�R�}B�b]v�e�Aw;<�\Ε�>N�����ʞ�hlW�JQ��9�jʱ��X��7Ty�r�^3���3����@__Ż����Iϐ/��;!eĘJΚډpg�Z�ʳ�=%N)��	�Jhϯ�={�=S��~��NAȋ���)�}6oތ%K�`�����}I!�����K��<����
�y�������r�-�ʍ�|.��b����ˈ}���Sr�A�h���O��.߇/pGJ�ʼF�^/*N�neH�����I��cchvv�R~����Z���|b\���G"l����0��1{��esB!��"l��؈}��K�m�D\��~��"��R�Oa�o���b,y�F~az,fן���b,S�P�!3�T�ޡ[��w�\�Z[[�f�e˖I��B�"���`�ʕ�袋p��c���ڕcNy�^����!whf|V!��=CM9,� �<�fN?�g���f���o��3��(>U���3��!�0�NH�0�6�S&����G��]!V���n4��_h�G�Jl�Ƽ�]�%ʋW���zܶm�p�}���g�u�ՈBH����������K�v�Jp�%H�c^������%_�%G�hgPW��(�jdPݡ�g~�1[��Zp�E�T�]�x����/� R�G�*��z�L|D����d(���vk����}�
������A�K["'�D���q�@!�����&��8p��Ҏ������+���R�i�B���Oa���12��Y��c��l�ܮ�e�p1	��}�p�t+��iuV������l_[�b��ntvv�B�t���{�/H-^�W]uƌck��b�=E�B�ꂩL��'ƒ�v�c)=C#����ܳx�)��Z�]���#����Ĩ)��� ����RL��G@_�?մ`�ڞ5�����H��E(m�]+Z���:�V�R�ڭ
Tv
F^��&N��;v��C=$	T��B��>���J��?�y|�[��	'� m+� ee�|'�sc��+�� }$�-�FM�]���ވ�lrԁw_J"S�2h�Q�=��!ZE#�ۉ�)��� �m)Wv��8�s>9~ G������x�ۿ���;�f�����s�͂B!N"��&ާ��+"�WZ�x���lm'���f�pXo#|� B��v�+����`��l�Y����:AwA.ޡ�a�R�
������ᩧ������c�BH!:tH
�?���R1�%�\���*GC�ʱbz�v{���y���I�B�3�Y!�2H�lrO�z��r,�P��v������F1cp*������	q�	)q���o�{t���L�ʵ��,�.S0loO`��䤸eǺS�仏<v��A<��cR�]U�B�S���ذa���/��k�����q�)+�"0��X�v��c�@{b�ئ�����>ԭ�6w��Sb=)V)��uE+�f�J�J��&T�8������r%2�hs����1&��LT]]]x?�l۾3�O���F�!�B���L��с={�J��b�D)�;�k��ǝ!��j!��s�� �5����WhWs{�7L��[(Ʋ��5��x�Z�����R�#�^x�,]�MMM �B줹���r������&.\(]�8��c������g��G�Ɣ�r�]��Jݳa�3L]'����}��P�T�6��g8��'Ϛ�Ww�3$�Mp'��9����vb0K�٭TF�z���p{��y��^�����⒗,yLLu�����.Z�!�"ރ֮]+���;�<��}ƌ�6�)+��+0��Éu;.�c�����p����ԃZ�Ji`-ɓ@ne�АR��6�'���@�'^!y��x��7Q�"d����;kp�aQ?~ �95���/hhl��ѣGcڴi�?_R'�B�s���c߾}سg��pQ�{ooo6W�w��턐�r�\?�3>�cYmnW{��cY�b�c���Xwc1��s�=�{������B!v�{�n�x�X�l���J�y�O�9��>v�ԋ����h�3�:�.��1�=Cy��_��ͼBs�0���|e�\<�T�/�B2a������B��!�����*k��Ԙq�L�2��:-�y
Tv�ӽ���1��#B^+W��ZD{;!����hŊx���)���
�;֒ؤ+d�BB�F�(��]/TВ�ݒG���XZ��1m���he��u��~�ޗʸ�����Oq��ٓ�U͡�9w.�k�`EH93����Q��� >3��k��b������m۶a�I�2e
&O�,}N'�BH�Y'��)��;������Nk%���~#������M�,�C�����;Tb��۵��c���~�_����sz������n�:��oÖ-[l'�RT>��#�p�R���W_�N8A�'����Ct�+ۺݡ����Ҙ}�a:ܮ�'�f���|FAw=�Pڧ�	��;��A)>T�)A�03$M��0�n&R�n�M:B�Yk�=�"\�	�	T�$Hy=�.�5k���;�����A!�xѸ'�V�^����
�-�<�W���i��m�PAKO�I�	)ޞlk�L���[m3L�U�kE��ӂ�<(�82�1*Ɣ�&�>�фs���
V��;�"~��W�)5CR���
��"^K67K�x7n�N��)����*B!�:���hniI��;;]	�E�}x��ۺ*�@!EE����uO��]'�n)�����F�X����>g������������w(<D�	!����o�--g�u���N�%�.��O1<E/e��[L�P�/LݿOn�J��~�ǩ���ޣb<�ڄ��ƪzB�'��p���Z����70��Զ/�E���JY�*��iqJ�	.Y�/��2�)B!���������˗���/�9眓�����v�}
	�[=g!��v݉лr��X��!Mz�L�R�G���׍��>�^��L�*�T����H[Ο7OR�"dDp�7��w�b��>=1��@q��"^S;::��>���'N��	��~��>!�22D[{;�Z[�`�����f[gH
���;!�n_\7�޶}R�]p�cYnn��+ƒ��,����@�ޮ�r���J�;��y�%�~{�}���C$!���}�Y)�r��[��&M�d��S���!�qL1֋Q���&Zܡ�p�Pymh6t�ZP�����,����a�m9˷S�'��0�NH	q����4J��(e RY�������)��*�(7�\�ٽ{7|�A),�FA!�x��%��������xu�5��㎓�e���c�1^Y/D಺�Xb1Y�Q62���Z�J�v��Ku���6ܮ����}�~�ί�˷#�;��@�B�5vW`w8�O����"�����yV,����_#�O��	�e��ц_�!�Bʕ��!tuu���M
�w�o�]�!Zڛ�Cx��=Q�ۄw����Ds���gh�ޮ;۳%�P��=�Y�Sޡ�oX�wX��u���屾�>�\�w�u���A!�x���<��#x�p饗��_�:jjj,���C�3��g���{�"؎<C��'� {��kH��)�к�.=��H����{pѼiX��B���a������ATjHNaJ+RY�ZP�����*U�ݧ�2o�f���d�8���H��M!���l�ڵx��7�x�b\y啘2e�'D+7֋�Ġ�&��#�+����S��<�,ZeG�ϐB�J,CCzb����=��m���ۢm;�p�l�dȝ�Ct�'�>��Qc��?n��Aw�P�5R4�E ^+G���;cǌ�رc1j�(B!�'�]Gg�l��pqfVɆ�����Jb���"n�;�����B,�`{^�a2��K1�a{��o(֡l��*��ipz��;��>��e�=��lojj!�R
������oǪU���o�w�#3@�b7;G�x�z���S�0���ɭ�x���I{��V�t�=��Y�T�]�˔ڟ�;�����.����!e	�B
�wBJ�S���K��CYE����S���օL�*o�J'�nE�*��� �A�h��Y���z+v��B!����<���R;�W��U)�^YY�x���rib�g���xZ��i	E�{2����Ҥ^ =q��(�S_��B��\{jϭZ��*��i���X��84O)?D�}kG���C~�Dk��)�d����Q�0j�h�gm|?�@!�xd���AOw����� �F������Q�C�	!���-�A��`�7̘�9��ڬϙ�a K1�ٌ��|��v�L�ʱ�;,�w(ظq�ܼy��q�B����_���җ����j|򓟔Ƴy}V�)$�nt�z�V�5���3�}}�=C#�0��/��#M����<�wʵp�>,�7��+r'�ap'��|Y��5"J��h`�>�`����˜V�	��+��ħBαm�6����k��Fq�BHY!f#���;�������SO��R])6/d[/�(e�ob,&	S��	�J�"��)e�J�bג:���U�X��*�J�|��a�V��zp79˷3�B�Hc`ȇ�����uc�8f\�Ao4Ɋp�XZ��T�"�.�⭮�BUu���Z��/r�����BH��W�Ed���ߏ޾>�ŗ��O�.�{������a���vB����sD��9~M_a:복p��w���V�enW��3��)��ɰ���|�)�8p ��s�/_��/�B!���[oI_�:묳p�5�uh�=E7B�����������J0�������ˬҧ�~�����X�X�AoX��%��aΜ@��	��~k{���jZA�Ԃ�)��
i_(u��Iqˎ�B�S�>�����?�)�K�BH9"������ӟ���~:���:̙3�v��.��f7C�`�)���u�p|!R�53���LO=�^���
V��2���[��yӰ�! �q����ht���Ǘi��8�L�����&�(�Yg������!������Pb�o�|�VW.�>�Jߠ�UH���a�B�A(�Å�{�h�hm�m�gec�v�g�R,+3>붶k
�|I�F�Z����Q����������$!�Rz�Ϧ+V������*\r�%	�3�h7=E'C�vy��mNz���H{�iIZ|>�b�\��d��g_:]4wV4V!ʐ;!���;!�̹~)ܞ���ۍ2�4�Z�xzA�p{	
TnNn	Z�iᩧ�½�ދ�;w�B)���X�n���
\v�e����Ip�Ǌݼ�m��M�u���)��آ�R�:�9Zt��P����C�]�ʅ޶}��n�7�8� !#�7���UC8z\3k㟉K�5A|V�h�%�B��}~l;T�]���g�	!�A����EOgk�3�!ܮnn�ll������b�5��9ﰜ��Ny�bٰan��6|�� �Bʙ��6�|��x���?��ϫ
�����}��;�^�л]��2�;i�0�ص� �(�p{.�3	+�r'�	p'ă�57��ܱCՠf$R�O/�hoW�TÀ{b���<*P���U�9��}�����͛Q%���/n V4:������s��_��_YY������n���wYXw7����/�[���7p�o^���^��뭛�]6Դ�߅�������o�s�Q�V�C�V��d3C1E)���z�	�im�r=�\z��*��0�}P��>���}XĐ;!$Ns ��Q�a��(�����n�%�BF��}gO��B�@!^�*,�ٍ���W�-��^��p7�吻�Y����*��"C�)�8ҽCyl׮]��?��g�y�_x&�2b�"?��}��v~��`֬Y���͎qc�X�w�=C���Xz���oh�/Ly��s��c��;e�w���#&bծ�3$�Np'�c�3ϏXkSFS��p��@�
��M-�k�B�;xU9	Rv	Z������;���)��O����ߐ�o��n>w��C��u��uĭ�����_{ܺ7����/�/F�߼�Ϳy�z+���{(n�׈�{����o~��Y�����1{��4/����(�z�E�l�I�#�|�F��ɠ�I���he% ���D�R�d�B�D�}�~�BZ&Ta�بx�wB!�x������� �wW`_O�m��R�c��C���0�s�k�Y���C�Y�M}C���^�{q�h���~�����?����ɭ� ���M�߆����ߞ��!����n޿���w��s��r1���.^o�,gr�o^~�+h*#�o���v���R���K/�%�\�����>�c�Z/ďtr_'<C�|��Mg�2���*����Ý��`���Uː;!6;!�̹�ڶ��@����&P��N-��Yim/o�ʫb�v],"���?�	{��Um�
��"�(�틍���p7\:���.~�n�]��w'�n���Y�y��@��ߝ�_�p�k������n����_ĺu�p����+�,X��[�r2_Q�l[�x���&!b�CFm�z(�7�
V�F ��X4�A���! =~B������JL�ƬQQ�3�J?�(%�B�"���}~���t(��a�f\$�+����gd���b�Bʦ��r,#�0[1VF�]tOl�¸K���-�ϫ^�޺��r�-ضm��.�������pص��߭��Þ�Hn������^�(rӻs빋�b����^��x�q+���߼��+�d�#�o>��x\����SO�G?����/J��}f�pb�EY����5�2�|=�Kم�պ���y�;�p��V�EĽ�B�
�	�g�"�ј��	����f�
Zi`�/ 2��S��g��xY�r;�n����؈[o�����kafB!�"�%K��oHm�����Ri^Ю"p�)J�G�-1&72H[��]ĺ��KL9�mf��(e.,)�W�c��'r_|�,���	!*D���? -ۀi5��UŌ�AT���Bq�����A��	aO8��!^�BJ�P���z���+C����À{��Xf�v�w�Y��_)�ם�<�;�C
�U�B!�x���z)�~����.?���B��X)x�V�U���>����%�Վ���X�T�(�n)�	� ��	"d1�n��@��,O-�g���*;�b�O��ŷ}�-[�;���� �B�5�lق뮻N����ZL�<�s��u����d�*-ɂUb�4�`r�Rm3�פ�!��Q61Jo�\X7��ݙf��}��/u"X'��3�rSj�0�:��5����wB!�z���ā� ��F�j'��"�~�lno-0ܮ�j��j1����澡y!V�ޡS^9z���z�����_����fB!��G�X�B*����q�EI�>�������d >�3To��Z�3�B��̛�=r�&������X����R��2'DeW������A�)e!J��M+������/RNPv���書�����B!�#�V�=U43,X�@%�h�y�\������ے{@V���É��m��h��`%o7�ޏ����m/9˷��AI�W�����l�@e �)ՃR�}R� �V��B!��	�����d�]�BH���p�~��[S!�\���`��+�#,c����7t+�N�P=������o�믿B!�X�������W^yE���c�)(�.�y�#�z�Av�mj�0� K`���8��+T��S�d�m_V]4g�7U1�NH0�N���:;�����p{�Ԃ*aJ)Z��T���X�B)Rv�O������׿�U
�`!�B
c�����o~#�V?��1{�lǛr]��(e�o>���<�_B�J�++�E��`�Ijj�*X�#"����Z�\0oVՃB,30��Ξ��*�1L�a��R=�	�C�c �BF:�+`~���P{k���ka���@���EnoI�bn���cۭ��Fޡ/��;���z���p8���_Z���@!���X�n�}�]\z���w�����C�'<A�z!�3�nt;<Ch�ܕ����7L\������ʽ�6�h��9S���C1ݽ!Y`����Ҭ �5"h$PY
��/�n7�Z�����N^�
Y���o��w�!�B�e͚5ذa���*\q��u�SM��{5�^�6��2������lj�$X�MTc�w�e?X�x�Ѷ�8�l<ɐ;!$O"�>��V,25��Tc\��WI-�����8!���oȏ�:#tE�#b�?�b�Bʏt��9=�M��Pr�g3��,��=BS�P�g�`��v1�����:��~�z�t�Mhll!�B
�����s�4#�(�:餓��|���1;����b{�v��9y�����=&�A��3�e���a��=���h�T��>��3��	q�/�aTw�$*�M�zU����������1]a�R���������tHK�,�c�=B!�8�h;3����O�Su�Q7-�^jM�nK��=��_�`���`��~�k4hדc�Vr?O�3xJ���A_|	�@o 5&��C1��Q�/��z�vM�g�?���B����P"����3�O-�h�gԇ�0�_B��@�R.�BO�A�7�z��<��!�h��a���S��a�]�z+�^�av�zgg��c.[��3>B!�m�6)�~����Ø1c<S��]/f��u��3@a��*u�(�Q���h­�pѼi���Rd>7=������4�R��n�ҋ�4ܮ]��)Sz�}�X���X^z�%�r�-ػw/!��<������·��m�����/Gee��"�v�Q��<�l3���	r���Ա|ꛚ�1��PmQ�i݁����S�4	!�0����V[#��*@����z�c�m��g����U�B
g0��4�4k#C�1Ѹ>0_��?�K��uB��I��C��K��k�Ê��!��7�l7���0ܮ��Y`�y�,5�P�ꫯ��#g|&�BF|���G�|���G�җ���KY���^/V��}�0a��y��� m�y��g��:���/�7˶@���OOab_#�`fk�B�2�����J?�S������R�������m�݆g�}�4XE!�gm���_�6w!Z͟?_��	�)ۺ�T�籲My��`S��a&V��V��i~F�v�̹s�\�!��}���sB!�B��n���&�a�����XJѺo�_�%p��+��S�b�g��Z�
�B)MMM��O~��~�����1~���ci��#���~�P��{�1��sG��!//���Z�bѼX^�iW	�
��OLaZt�xMR�@��n0�H�K�=-V��� UB�v/
TN�SbY�z5n��V477�B!�"Z�����K/�D���*GE'���b�RV�ɂUz�A�
�6���,d�~a����۱�F�2���!�B!�B��º�nW5�+�C�ٞs�g܍��f�a"�.}�������_|�E�;ܳg!�R|D��#�<��k��?�!�8�U�*0�z1��J�3�b|Xnp�x�>��Ɏ/�Vk瑯��G*�Be9V�n\0���g�)!V`���"P7>����Č(���)u��3E�@���Xe%ܞ
�g��<��	*ۺhmS
�Y�&34E!������=�܃w�}?���t��ˡ�!����n�Jy_Z�Y�J��vYf(X�o�����s�~C�B!�B�H��y��q��Vh�B�vP^�%ܮ_���!ʺ���v��@��׳����`�ҥx���B!`�޽��/���>�_=&N��I��ʹJ�3��"��T=�P���5���ؖ��=fҊe��,�_�uέ;O7𚎐l0�N��L�ǿU��`t8����^�H�R�ۃ9���1��v�He%��T���*;�|����?��o����B��ٴi���.�/��r隭�����l�[��1����u��^�)��{$�	}M���s���(!�B!�229k���M�R,=�Ь +�p��;4���v��(o(�C��� �~��ޡ@���b��B!�A�W�^���~����NS]#y�#�;��x�����ɞa�i]�"�3����s,��=�0N�}'N;b.^��b,B�`���P�ǉc�1��)����@f�=hw��0����/Rv�Y�zGG��<��� �B�������ߎ�����?�9���<��`��U��N+���1�s?1�O�Q`���O��[(XB!�B!#�/���ѐlOy���(�L۝	��c	2�C��K!�n����)y����B!�E���p����O~�1c�x�#�zl����l�v?�v�3��Vy�:!w��1�M��Ġ�3�~t6��Yuxu=CB�`���]�ǩ���ۯj`40�/�-��@rQ�18n�n�G_~�v��ٍ�mذ����� B!������ޒ�ܯ��:,^�X�heE�Ү{A�2ڷ�m�VYZ��*kX���%�J!ZE"�߅����N��B!�B)|nz�5"Taɞa��K��S�	?0�G1V��v��(�ǯs��J���!!�R���U�V������~�3�x�Ҹ��v���� ��y���@zfA��+����ZL��tn��%�.���i�N��{9�3!z0�N�T���Ξډ��1�`R�2�V0cIݝ�'�ţ�n�C\*'�*�c��0��n�w�}!�BJѦ��?�7n�~�L�:�VQ��w�ڭ��H�R��c�[�@yU�j��R?����H�W������w�!wB!�B!��9~J����t��v�0q;��ݩp�<^.�v/{�����^�u�]x��08H݈B)5�����W^y%��?�555յ�������m�z4�&<�t�=f0�]!w5�׃�XƸt�Dpxd�;�l9Ȑ;!Zp'�fB������쒚��۳TF!��U�p�|�PH��\*;)���-[����MB!���<�6oތ믿��~��*�I�^��U� {�����{��V=25����t��t���M�} k�&�%<B!�B!��'GO
b��.�|~�`���=�GLy�����z�a>�v�~��v�ns�X�uz��BHy �����c�����/~��;.o�P�^�л�����Tz�Z�Pr���Y�f׊�q�pnl�&�BC+C�(a��	��=/�ۏp{k�(�jo׈U����L�=d/�p{�)+��YѺ�d�����B!�������_�_|1����a��ўlb�����ؔ��!X�"���K�,��|n����-����)ڱz�0���#�B!�BHi2�� >�߃��Xf)����u}À�?�y��k~���a4�#�<�;�}}} �BHy�u�V\{�������/�\��s�#�;֋���6������ܕ�+0��2Wl>à{bc�0r?.�c�cOg�!D�wBl�º(z�&��m�!��v�@�h�t�=!J��KZ��/ܮ�Z��p{1D'�)��޽{�����úu�L�O�B)m�P�裏J�K7�p�=�Xך���`W ފ`U�ԃZ�.ٲ�2ȏ5��1����c�=�8oj+��B�z!�B!�R6L�ǿW��`tȴ��7�C�e��_��v'|�R���;w�č7ވ��z�B)?z{{q��cӦM�����ӧ�j���sٷ�<C�}M�r�=���	�+=@Ց
�0�3Ln�D�8a�r�gBdp'�&.��(iۋPEe�H���Su�=�6��?��n��+gE��"Pɷ_y��z�hjj!�BF|����i��ˤk;7��s�׭m^�r")\	V�XJ�J$Ī���CX8;�e�U�K�B!�B!��W�ǉcZ0�Q5��b�����@@�˟Q�e9ܮ�GZ���av��^xA*���� !�B�����k�a۶m�����|Eu���G�]�gh�g����)� 2������}5������	�x��?"��;!6��#��5!2hn�,�&��ͦT�T��S��m_�m̥K����CUU!�2��
�/�}�ᇒhu��{��!��d�Vʂ���k:�} e+��`e(Z%�*e+CO�A\0o�o�1|O!�B!���S��+S:��ݗ�+4�Xf��z,�����b,˾�N�]��nw��#�n���Ӄ;��V�B8!�BFį~�+�������kQ[[k�G�]��gh��U�0>(y�6c�/��_,�1L?~��D�g�����X�{4g&#�	)��N��P#�������4��$R�X��kU>b�����V���!�BF.����G}$M?x�I'���`��U�UM��wu�ݬCA��p{j9�����ƹus�t�$�B!�BJ��χf�!�ѥjnW.b��7(�c��n/�?0�p�֭Rk���Q��!�2�~Ճ>�M�6�n��������J��ݾ��g����
�����[1�2,e�=�����pW'Q��*��>2Ra����?9����T�Qs��􂁌����`6�`��ۋ-P9-H)o�RѺ�?�	��� �B�ڵ?��q�%������4��ӢT.�C�2z�vVv��3�\���к�p%?GE�=��mo��Ś�!B!�B!��X8o=�͉p�N)������>���J��K�`1��B�z�'p�M7���B!җޮ��\w�u��׿��t���	�d7�f��v��)=CO��r7�˖��9�y���ә��� ����z��ȅwB�dƸ ���Ɛ�o:���(�����go`�;ܮ�(�v�����-�c�����?�O>�$!�B����'�����_��f�rE�2ڷ�m�llp"�n$,%��n%��J�2���E)^�~��*�Ww�������}QB!�B!�48�}�{PQQ�[�U�e�g��{�4����#�nw𽥥��z+�z�)B!�����J_~۲e~�ӟb	���v�Av��x�3T�+�%���B��f��,�/Ly������8�nVs�g2Ba���<8�ڏ��6c``H��]!PemoO�SE��U�����^�r�WL'����~�!!�B�X�n���j)�~�i��E�b��!w-�s
����6�~���T��ah^t�i�*D"�݁����e�B!�B�6_��P[#B�
��v�G����,��r�;���+��o��&n��F�޽�B!z<��3���ǯ~�+|�S�*�g脟�g�\�#�n��kו	��jhm�]{\�_��1��g���]��ȃwBr�*�Ws�����%�t*K��z!����Y��R����*�"C4��oVvww�B!�
��Iܿ��o��k���/K!Ȟ�6χ��q�t�=��{RtҊU�N�5�rQ����#���š�S�����B!�B�W��� �:��bU�x��Y�����Y1VΥX�۶�ʱCCCx�Gp�m�a`` �B!f������}|����e�]��{��f�uz���,���u3`��]}ݧ�eQ�<"������!�~��}\�	�O����r'#�	Ɂ�/����<��FPO��k`HTV���{6���v
T��zzz��=�P�vBH�"^c���v�z-> CA����GͨZi���ae~�AFq�x�H���h���G�]��{/�mۆn�ӧO/�(et�B��-X�r����Ě�n�ߖjE+�k<�K?�X3=�B�����{Éc[���$t��B!�B!���	AL�	_0`\���;�bɋ�g����c����ۋ����oGG�T��z�jB!�X����ӟ��Ѐ���7n\^�v�˞��s�_^!�gV��L���tP=��R�d�5~��F�YC��3~�r'#�	Ɂ����ڒnW�܍��u�uE*���I{�R�A��bTV���Ԅ���wظq#!��xݭ��AeUe|��^�+*+��V�ە����4���� B����_�gE�D�����'9,��M۶c��G*5�+_W����2�����M4I��F㷓�`��il@�9�9Ab���!��o���}�{R���'��(��y��=�b����ۭ�U�ǣZ��R������l�F�����W���=��^E!�B!�x���8�b/�P{���vc�PY�����e�0�R�R�;��3��e������ZX	!凔�P̰!f���X��t��\�3���@3jg�w0*�@�L��4kphC��%~[�
�c���I�9b�eBʋU�V��?����㎳��e_;<C��s�wt:�nt�1��b����)g���U>�|��qi�Qc�[�~����0���ȀwB,r�<?z[vJ�G�p{����:��n��2��:�
�C���^x�������B�7a��j��֢�v������&L�~VƷUUWI�fdF��r��xL`��	����"�p{�>~K�S�:�Gs�����c�QuR轿��}}菠��}�۽�=���	K?	!�k�.\����kp�WH׊^�̶�-X���+䞥�A{=�K݂�҂�,N��*�sd܇R�J��ub��*<�!�B!�B��j?Nӌ���~1��K�g�W���٬ˬ�����l��W,˗/��7�,��B��xm�Q��,Œ���vQ��L���m��6_vlo�G��nD�]�`� ��s0����0+"|¾~�,K�?E"�m�	�6"����@�,X�q�V
��ٶR�[E}�S�?R�v3�0t��(^�O�Њg����8)p'�'�b��!-P�U�Z���T�`ZA����z�
&�%��X%�eQ�����s�=X�t���hBH����ѣ1f�Ԍ!�T�֢������ޝmm��ݎ�8�8s.�����:���`�O��=c��q�`{F>�����3��}��Ĩ�@uu��(w�)���8F_o���{z��FO8�t���>��L�Z3:-��%[�lI�|sB�$�����'Ɇc @��l`CH�$˙d�KHv��`ccl�C�-[�uߧ�?�=�]]]=�#�)�ߏ��S]]]����zߧ��BgG�QM�ID|`A�Gy�\17������ډ�@=Ҳd�b�kZ��*־��0��f��^�?1Xe	�u����
7��{�⼅���n�AAAD*��Θ݉ޮ>�Q����)V�)t�,nW��r1_8�����Ʋ���?�0�{�9�z�h�M����'`x`Eӧcڌ�F��B ������Y�	�75cn�<�lp���^�Q��'�E�9ϴA����Nlذ�!���P��Q�0�<��^���]���E���w�%��g�0��Ӄs�s�B]Fu�:� &$p'�(,-���Y*���W)pe���
FPq�1 %���a�^&��
J%3� USS�q���o� ����/S�OCaQah*��:u�1��v�gYu�'ڳ��܉Y���򱺶k�B����]�D��O*W�Tu�n��v�Ƶ�jY(*��T:{�n�8�í�9�ww���ۘ�ԝm��n_�}�+�����z�_�˖-�{�IU7��7&��OGu��=����Y�*�# �@��Víu8���5�� � � � ��������{��#Mf�0�0�
:\�#���<��+���s����&2��k�.�u�]غu+�H�z:E�#M-
�M1{�����MF�q"���s�g�TL������=l����'�:2L�j�H4�~���Ǟ={p�m����*�B�X��Ĝ��>Rΐ����!�tqgm�?C,�0���?{�y��|!��;Z���xi	܉�	�	"�Xlݔgy�<��r�*�pmz8/d�w� �,nw�08���hq{�T~�W[�l�w��]�߿SB��L%��>�N�j�3#�1��m����x��|�#�'��������y���yv]E�#���hi5&��J�� ����'�vĀ���v�~���툡}�q.u�e�mس�Cu��]�]����YZ�M�fL��0�-6�!sy�7��P���)�"��y��˶/���Lض��+U��T�֤�z��}oll�5�\cA�v�ZG�$��D,K�z��܍��A����Z���;X%׳�S�IX��b��jlmAAAA����-�F,��a�#?�qo�M��s{,�X���&`)��1V����)?�'w��?��0�jkkA�]ۘ}���(�65,d��E"9�� v�٤b���0�b�wf���م���Щ�S�DeӦM���G�|��8�Ӓ*d�2��X�%K�I�B�џչ�pNWN�/�G�m�����?���^����-1q!�;Ax��v�Z܆���q/�Reyܹ�=zpJ��Bv98E���.c�o�[�������x�G�����|�L�ʾC��w��f�&�M�Z��=UwC웛���3�iƌ�z���Q�k
Zp�]$�vsŎ�6#xR\Z�lג�;�o��ڝ�P�d��<�v�cWu��B����5��]��"a#v��,s���\vp���cdt��������n��H��R��g�<������d�lh�T>\����[F"���y��nP_��׌{��:1�gY&�"����J�����>��k;28�9�U�9Ȧ�!��>����n
XAAAD���� F[����>�"v����y�9COs,1o����Oq{"���<��>��Sx��ǍXR&c��S*H�)X*Mr�w��G�� '���5�4�2��S,�Qn�#&�#̭�Ә�
s"���0ͶR@g{�v�Iɶٵ���C��	�Fax��9�s�X����=n��L`fY��YOf3��Il�8��,�|�wફ�W^i�W��3�3��,�����I�.�
�����v{9��y���G���k�a�7�^��ʫ�N#��ALLH�N
؏��UC�m�����s�-r�;��r�N��385���P1�࣏>�'�|2%hD���U�%31-,dg���mX�x����%]|c^�t������vE�B�csm�.�R}�I�\�v��_0�7 �ӽ���>y��]��ڎ��Z����o {���t�4��Gttvt������>l������x�	c$�o�%%%)sb�� >�+"wi���o�%|�F�'4����r=�r�����������L��ȝ � � � ��� ��j�)?�0�r�y�0`Or�19�;F|����D�c]��Յ�������;L�Y;������"��`�4��G�K)=���PR63fcFq1��^�%�=t�	�S�PP��3�W-�Iɶ���q��s+�d��u(�7���bn��mm�H�̬�e%�+��y~O0�̙2a��z��� uuu���PTT4n����D���5-��?[b��D��ײ�z,�Y�ݭ�3�#�DAw�PpA�������؜��Ђ^�Fs`�<�S���� U��R��Ǻ�СC���	�P���o�Kf�����Be��{��'���jk��bjM]�ol��k�[d��k�bM/q{�]�5��:�-/�^�i���E�\��ܖ] ��2�G�T��*{�^跌��W�T[�����r��-�hi>�CM�)u '�t��#��ۇ���cٲe	��uY:����͠�5����D�r�E����wk>��n��9��So�������]�AAAAĉ�),6bd8�!f��7t;��e����۳�|����#��eR�L��`�e������;�i�&�`v3f�4�졉�
��P�{o�D�D�a�SS�O3���F��vwv�����	ߓ1"4Ad2����iܛ���(g8�u8E��?�W.r��Et��F��2K�6��4���!��9Mh/���>2�"&$p'��0�R�����:�G^P�`��󲸝�s2Yܞ��۷cÆ���A�	�3��Y������9��Zᠹ��{�\۝�jaA����Ĺ�;�����]۝�v�k�)$�kٕ����+�O܎���k���hn�r.��hj�1-XXc������͇��Ԍ��0�Bg�H'���7���r�-8�3"o�rT��,�V��y��~��Z�^�#�<��W�JX�2+��T!z�����C�=��tM>^�Mw� � � �HyAങm���4ƒ��y(�۝BvQ��-j��S,����[�kN/��n����o��;���� �MaQ��C���3Jf:�������UF�3���C�����H"R���lٲ_��׌�ᩧ����a�e)g���M�s-	����,��T��l�9C!�444�O���o�O�=DL H�Nk��۱���w2�T�۽��5����I�nϧ>�����xTlH�{��b� &3�:�Q%����M�"�`܀K�񤺶Q�]��{��r���%nWu�[^���M�i���������暳̽��ޫ�]&���u<�]-++Ms�b�Y���M��`�7���ALV:::�`ss���+�{�x�=`e<X�kµ���Q$G��y���]8f�pq�Ԧ#���C�`��-�pFu5^�K�^AAAD<a���W����!nF��b�@��m��@0�1V &S,�9�w���3!?mi�������}� 3�X\Z��ٳ03�ʜڳs�A�B�s����a�nAkhb�A�W� �C������W_�/|����3��,�y�t���푞�Q�a��W��K��ς9/׭bĜ!o�O���:qAe>��C���ā��bZ �G��H�%��]5A������r�eׅ�C
�Yܞ� ��?��{��"&%,�T:{6J�f[�(M!�v~�Q�Rܮ��we�jܵ��\ۙ[w�I��n5/��p�R��C�c�O�vCt.��vy;^�|Yܮ��Q9����\�y��]�pIhZ�ب��ى��8x� �����L��9~�a4���k�����IX1����K��]��DsdP�sF
XY'ɕ������X���ű�5�{#Y2AAAD����im�tn�:�s�����3�&pW�b�yC�cw�p"���������������1�	f���-S�ٳȝ�H:�ww��9��`����:�d8�3�;��d���=���ߏo�����O��a�6Ɠ[L���|�ոG<F8�Μ!ˢM�����y+��� �		�	"DaN�+:���Q��#�T�<H%����/A*y�A!h%��?n��v��.n����<�_��W ���f�a��}��2)�)�زf;�k�umR�,h�צ񺶻���������e�T@�ڮ��?��:s�8�ݧ�Eum��O�v�k�k���'vV�<�N���ӧc��%FQOw7��1�{K�!�d�����׿���q��c�ܹ�@��%ӱ!=D�Z���{l��]���|����M;`�Kx����01w6��ˇ��2����&AAAA��ӫ�l݃��W�З�]toL����Y�ܡ������a��!q{�m455a���x��A�v�*-��Yef�pz�G� ����r�lZS����f�55�dlHL6�}�Y�fݺu(--�؜��z�[_���u�6	���f����eR��Fݱ��i���X���"�!�;1�aOX���Co[�Z�*FR�������T��ݿ��ʅ��w7�4e��
DeJ𪹹w�y'��׿� &:�S�P~��tV)��k�
YܮKK�VU�v�[!G�\���Q��a��mJ�E�ф�*!���<�i7��.��Usbvmw��%<�[�ԩXĦeK��{[��1��Cc�~]�u��J���z�~��[oŲe���m�o�x�#��ݸJ�j��*X���z7wY�΍�y�	�@U��d,���!�ݖ�����AAAA��e�A�u�"̎*n�ruX�vٹ=K�ǖ7�l�%���q��"n�G��߱c�!���AL�u���g�)S�bDf��Y6J9���\n9��߈�����C�BbR��k����ظq#�,Y��9C���>{k��%�U|�g�?�3��(n��C3����6��ۆ�-?Ӵ޽X4sv����DfCwb�s~����C��풘ݽ,,l8�ݢ�,O�����\��LM$q{�쑖�ڵ���W�����C��T/Y�9��hjQ�ڈ�k��[X�,�v��.��Hb�q��]�V��M���8\�M!�%׷�E=�]�8��;�������bgE�sAگpG�,s��1��N<h>xuu�ݽ�� ��FCC�����[n��g�9�U�e�,r���D�R��92DO��nl�2^��Bw��*���M���8g^>���3G� � � ����)YX܏=�S�)���{�3��g�6�r	�yC���63!q{�˘(lÆhooALd
�LAY�C�ΦS,��TD�����tک8�Ԅ�����1Qٽ{7���:�p����>��9C��'r�Ж[����q�Q���P��l-�r����:�{c�X�} �eh�;��TH�NLjN��P�oq{80)Pe��;�����p_P�0�^��@9P�Qd���,{��׍�)@EL4rrs1{n���bny��TzE͂��Esmw
�!�U����xK��Z;�k;�`��O�./����-�wtS�,�v�~�H�k�(&W�_���ݵ]�ɵ�т���x���4E_���<TU/M�8��G[�a4�գv�^���� &
�����{��e�]f�c2��#QcY'^"w�9�M��V�ۓ�ً9��)n��y�*<���ۋ4��ƹ5��nAAA١?�O�Չ��G�0E�.`��Àe�������b���y���2"��)'���`�z,���s��_��_08H)�ă��O�6'-[b�~	b2�����U������4��lj=�QgC�HGG�!r��w��K.�ĥ1�w��O��K���s�G6���{k��?ԅ�!,)�����l��3fwㅺ��1�������,�D�@=4/a{�@U �`��K���[�.�g�F�Jp\��VV�څ!Q���(n� 1Q�RT�y��7>���R��[M�\�5$͵])$��!nK�����'�N��brm���
��p8�z���>j�5��?��]ؚR����cum�����\:{�1{��ho���z��p7�6� 2���a<�����;Z���%T��Ht i,������k���<�U���)Xe��%G�p�<������j��G����h�A� � � ��˧�G���a�ۃ1��Y~P�Ypo�k�%���ڕ�X^#?G��SN0��,_��� �<�b"���U6s�S~A>�v�!q;A��:}�1-Y������C���݇��A�3������~|�[�2�s���F����c��?{߿"l�%�c����?u�0�н����)�Kd�Ed($p'&%E�YX3�	Cp�ڃ�80X�����`���^�A��9V�omtq��d�G�ǞN{����SO� 2�¢B#5��ųJ�r[��丶C!n]��]˔}�uy��?V���b|
ۍ?_����G ���~Im� �0.�v�X�k��,�k���横�u�;����j��>i�:�eF�cZu����`_]v�܅�#��D���kmm5ݧO����X���^�ږ-r_����=9X���,h���#ݟ�e�m=h��EΡc�JP9���$r'� � � �h|rA�-���*a{4q{0 ��v>Q�3s�ޣ?˂v�(K�b��+n��l�v?����ꫯ� &y�y�;�a�U2{�k�I� �0w����tdt���ذ����& �_KKn��1�#-�$���XE��,nמ7���/�e�%���=gȄ��������QD�Awb����]ރގ�1�����T�H���,�}AZ��ۅ!ҏo�瓵~2����O&����Ad*�)r�bC�M��Xf
xn�.|����н��pmR��.��ua�HZ.w��!��ro'v�P�]}<��L�k���p=ͪ���Q������%�:ˋta=sU�Q��Wy�uW?U뱾O)���+W����kOcC�|��{k1:J��ǟ��'477���FEEEF�)r�X%���Э�2V��TA+�����n���&v�PY�����S|�e���c�4���]���AAAAx��,�����|a���XcS,o����yC��a���bv�}��.ng# �[�۶mAd2��3o�a�5{���8�
�V�ߧ��ߊ�v�������� �L��:�6`����3�:�j�6������϶���t��v|��ãAv�aiI5v��DfAwb�q�B=--�����Ә���<wY�)@�r_�DA�Ӆ��8���Bܞ� �I[�~=6m���4���	�+��[��Z�'��v��]%��E��>�;�h��p��.�)�s;��Ph\��*�v���X�ǵݽY��{?uE���mW�4Kq�I����5��4g=(]��m��fwGjk��ݵ_�J��>��jj�v?}���E͢E�480���Z|�m���N�K�]s�5��}ɒ%��g�Q~�%#x�G�.���e汓]ܳ�C�����*��'/�Z�T��}���*�ŋ�S0��]'� � � ����� *�F	�an�	�CY��*W��f��M��X��!뵙/t����D2A�>��`�z,fv��"w��D�b^U���>��A��;sV�1�>��nAc�>��v���� 2�͛7�;����.,]�4�9C?m���]Ŀ�=��0���ʣ?k�|a�џ�W�9V�������j#�����X�݈�eh�;��H�NL*>Z���ûMq{����)@�}A��n�?�p�h�vU��{��;w�4>{����-���A)��la�7��ڮ�%nwmZ�����M�D��C!�v���%$W���Mu���]d�]�U����bn�wm/ѥ2�E���͸����4���|]��b��T��#�]l+7?K�/3���>���aǖmhnjAd�~���&6n܈�N:)��u���-r�
j�E��u����B���)�ٞW��ay�J��6|M�UO{έ)�ov� � � � �� pjq�z�=s�^��\��;4��bsn��s��2u�0��t��*����q�w���ĉDf��UL�^Y����<�onI�{Ǧ�����6c�}���QAd
,gx��Wǜ3d��`},��K�.�����o�?[�>k�Gfx��l9�C0Â�<!�
���ϟ�Յ
1Bw"C �;1iX83�i�{�%�������C@p_���GT���C2b	R�%($����X�mݺ��r�m�HxP�9�3���h�)��\�3�\ە��Q��x��C�'[�m�K�k�K��,�v�$��C�����n.-(���+VS{{;�|�;�mGWg'"�imm���_o��]�6�n~�e��ݹ=y��!9�_u��U��������v+`�R�S*j�AAAar~�0zۺ��v��ݕG�	�R�P=�stc�,���*�x�c%#�7���/����Z��ߏ��<D�îs����s�8rA��3���9�nj6���cxx���^�o���K|�l��d�/����{�g���U��6ms,����'�ź�\!�z��p~u>^� Ad$p'&�9Y8*�4Y J�<ە�(�Ђf`�����Q�`U�;0�zn�%m�{���-(�����Ђ �t�}�K�f��f�+*��L4��]����#\��+;�ʞ�v��
1��>;���>(���z���+8廉��&�jA�?�v�v�;��G껣�(_v>�y<� ����}0�������u.������]'Jߥ���˻z7��ǟt"�;��:���w`�@�Joo/֯_o<�q�e�������XJ�<{�;.s^E���M��W�";���(#@e;h��G�{�f�աrz%�;FAAAA���k���r 9��Qs�*��@8wP���X~M�����C4c�v��)��&Q9��l#��D���4�x�	<��#�<A�3�PV>�q{ @"4�HW�o�9e�4r��ۏ��z45��J��=������6r��A��3�I��ݙ/4J�yD�8������N��r����=���tD5���[������������Ĥ`mE?z��L���k�A1Xe/p/�Z0�
Hy��;�ܮ����|JEP��:�c��K/�� E�)�S���T��j��
F3�º�D��b]�Brg�\��^[%�p
�]�AW
�=��Z�v]�w�k;��O/q��OBr��v�L�hS)܆[����.��E��s�\���v}�V�&���/������2���vg����?q%��Q��z�a�Y����}����� ҍ���>�������m��fZ�*m�E�Z��Sts���5� "���*�"i�xpJ
PAz/���"`548����g&(^EAAALbV��{]#=��Jq��;:r������vA����ܡ��$k>�ǫ���z�!<�� �tf괩���6��|a� 2vO0A�1���������Bb�HGX���DSS���jCW��9����D�>g��X*���Q���P��jΛ���rS�.��8	&YY]�XZ� ;SҐHoH�NLx��d���	���� �/q{@b09@ɅAv\��VV����L�.�t	>����z~�ӟ��G��(�S����WV`��j̜Uj��S����n\�a�9�k���n��K�n����#�g�;wS��/C)��ݵ].��)���x���tm� ̏�w��;�k���¾)>����?_׹��O���Oe�5�����v�ל����U6�KJp��?�Ύ��`;>غ�== �t�g�A__n��c8�LX�m�$B�n��o��!W�JzPu�|u�2��O�X���Ἢix~7�� � � ��Ɍ�,,�:��`��J"�H�v{�g��=�1V$�v��nq��SHD�/Q��T��\I��>���7"������
TV/��Ad>��X�t	�Ο�C���{j���"�x����ڊu��aʔ)�y2F2\�Ǜ'�wn�k��̈́EJc,�G���q_�#?��23g�p�a�;/NG#=[�B���h̝��A݈H_(�MLhV�Ά־���AQ�.�\�)G�J�#/�e�|�����@�xF"��J�:��B6� ^� ҉¢B�*+��WA*�x�]��f<*q���) �����ׇ�k�R��
���߮F#��K�g���)X���FT��p	�!��"�ve]��]*�$lw��r��U�N!���x\�UsN%�Uյ¹#tTފ�37��ӵ]:?<��l_��A�i�g��SN��9	���a��7��;�V��W�BOOn��6et�*��r��YƯQ�u����C���#92�a��`�����Lv��.��ҝ�v����gTW�ս�0(AAA1���N?��=]C�e�>+r���k{0<�37�
�D�\��K%h]�Ŝ�#�0���d��Zv��a�_����@�Ƭ9eX�����!�۳1!�RX����}՚��߰u���pS3"����~gc�{�3f�4�7�u��E+r7s�,_h��f=��?��k!	ݝ�A�K*��/�?����}xn7�C�/$p'&,��C#��vPJ�<��f���v��rap
�Š<�qo�ma�q�_�1���u�S�������/� ����[1Ջ�pjz��q�?��nV�!��k�Y7��Nնk]U�L�_��J�,���r�NY�C®�vH墛�&W��ס�U]�{;Ϊ�|Wg����!��?wW=�a����sQ�����z�黠]�� <���Gw�qm�ͅ�	�+�0��2t=�m`��� A��W_}�8�����dt�*��,�m󺠇����<J�`��t�2��w���b��U,XfMB���w�bYi5�Ӱ�AAA�$��ݭ��	c}��d���s�����?�"l�h�%�Y��i2�����x�8p 7�|3�n�
�HX,oμr̫����� br�tGl�61�@��=�ݵC�� �t��^õ�^�{�eee���1���*�mE���l,���������򽬘/G~�-�r�QF���\���zkk���rq'��ÁaN7���� �jxA��/�T��])l�>��%hU� ��r�e�It�*Ձ�X�a����/��2"�L)*D��E���Fn^�Q���k��7����}�����Xׯ���:����06�vsYl���Ϳ�-�>��t�]�U�Nq�s\�U�w�p���q�k8ޮ��j�YO�w|����[y|�z��X쥭U=� ձ�%���*��w�S���vT}�M���?�{҉�W[���mAݞ� �T��o��o�ƍ1w�ܔ��E�!x��d���,|��$w-�������]�y��+8�%rwM�;��l6��,t��	� � � b�qlyC-{|�U9�@ `���GV��,c�5Ų̱��!���D��D2-��ZV[[��n�	�v�A�3fc������Bwg�i�AĤ���:�h�X�
�5b��8t�	�j6o�l��+++Ǖ��[/Y"w�D���2�u0�^.�zޝ3�.��{��{�-��<�V��s���A2�"�����#90��T�/$q{�����~�t���v��=U"�T�bY����peOD*)+��E˖a��2�rݧ`]7+������;છ@�vQ ,���b��sA��(�D�b}I��Aֱ
k�>~���T`k�������w;~��ȵ=r߅�9�>G��R�n�9�]�-U5ա�---x��M���mA��M�6��3VUUU)�'*x5^�
���(q.�.�n���Y�tqĠ�3@��9t��+)X580�O�����|+�FAAA��)����E��=j�P4�
�"vU�p���Ǳ���.��t��ر��744� RI0;��U�Y��fLA�����ü�
cjomÞ������#$4%R����q�5���{�ŢE�&��=тw�����}=wq�yC������_{�gu�P��a�)�/�G��`AZ��ɝH/H�NL8�/��P�n����y��tl��UkR�kxA�{����u�ReZ *��>�[o�o��6"�?6���\�b9�N���c� B��}��Q]�b��B��|sQ�Z���[��^sl��j�����;�:ŅΉsmw���G�;����]W�K�k�]�9��^:��}u�߬6V�vm�}�W��Jq����wն�����8�3p��>�w����|=�� �d��,`�D�K�.��"���'�6:��.�7w��IRq�����΃V^�`P=� u=~��ނ��U�ov� �� L����n�<����t����-|�����=����Q:����!���>�ͻ� � ��?�O+mG_���;������v���+�)�h�%������#1Qr��e���[nAss3"UL),D��X��u� �/l���N>��;�{���m;���	"ٰqX�����ի'��=��]d<"ws���P��,c�M�<F~�9Ax�ew1_(
އ��p��.�X7�d�E�$p'&s��3T?f�q!���C��CR�:��;h�z�Y�-tO|`i,��td�߿�֭�֭[A�&� Ջ�f�"���zֳn`�����f��7�����}���n������rmג��W�5�~&ҵ�YW5����;�ێ�0_�^O�c�x��;���� ��d|7�Bv�>z�]�^�w���ꃺ���C���T�q<��煮/��9��>
{w��;}�(C$���:#`u��wc͚5i%rIa���?��wV�ְ@zP����yQ�.��T~�Vb���nۋ5sb;HAd8L����_�I�+��\{ɩ�^��[~�rҷ=uJ^h�y�Ȱ�{��/���¦]� � &7��9������*�r�jq����1�����ͱ��He~1����o��a��F&�T����-���J��AD�d�dc��%�M��k�N:��H6���V��Nr��&�V�8E�F�s���;߮<�2Ĳs��s��\�"g��=m8�����HH�NL�C��S����sdLjq�-f��T.1{�v�z�=V��OA{�Y�w���7ߌ={�� �Iq�Lí}���)Sh�f�����)6�E��b��B��|���qvm7���S�\ەhH�k���ǎ��졦,soGCl��
��b.~��vU�s��~s��zv5]:���y�]^/��[�v�O"uq��.�=Q��Q��o,\��B���Flz�]�ڹ�,���p�u�)V���K K-r���]l���vq�2DzP��u�I�r�<��+�F4̡a	Lx9<2�ށ!&��9����	A������'.Kq;����C=����"�L-�ų���"��` sgNE:��݇��A�!/'�iS��G��>AaN�������A)o��/��@x�g��=�O�9Cٽ��ˇ{�ʵ����a���Y��#֯_���>D2a���h�R�,-AD<a�s�SG[�!t�W[o��	"Y��������ߎ3�<�̰b�h�e�+󅬢`����s��M�n��,�'��z�4!��o�����0�W}�����r���vu�*�s�g���i��L��S2��~�!n��444� �EɬR,]�e�ч8�Dn>�9����]ۥz��Vs�e��D�������$�b�Lخ��T~u�^<\�]
k��Bl� �%����>v��x���oG�?�vu=W��ǵ]� ƶ7�����8A��r�7�r�q��8?T�tn�rm׌o�e�,a���}��3�s>�WŻ＃�����QD����7��N�+C"E�"�Xi�F���ӭd���]re�T�,��;�;�+X���*.v���a���"����|����՟Ƽ�i����v��?���^~ã�/q������p�E�`IE�Q�x��<�[����{�������5�t����o|uM� �xS������4��휛��	��߂��u;��3QE�9�<~��q�q��4�t�[��k|�	di��O��`���������{� �T��x���9�s{0,j��oc�H��	�`����^��Tc%#/q�K/����CC�02�<؃35K��y�{�$� ҃���8���`嚣�k���ڍ�!�ɡ�����s�!3,�nc,Y�6�
���ݾ���<�w>Qe�e9��^K0�hv�&�H=$p'&ǖ�߲'������#�b^0"v�tj���ܹ���۷�h�w�	ڗ��pn��8n�=�����˵=\S^ٱ~b\���IqmWvJø]��n��v�f	��#���\۝N����w<��=|�|����vݟ�|.H;��|U�u���\�}w(�.�Aq��e��d��������q~���יQ<��uN<�d���&��λ��!X�[�w�qǸ]�p�I]��(�u���T�\ /���W/w��O��U�+COG+�V����{���|�/W:���@��=w}�l\u�q��~���܏�E�����Ū�2Gyy�4<}�e�����g^݄tᴣk��-�ή����<�t�U���'Q{�/����۾��WT"a����ع�0v�o&��=����x�p�'�������G��g���*���ጣq��V��_���W5��	�0a�>�PԊ�^&Bu;�g�$n
�v/��(�l���!�R��X�t�G�;�����^0��### �d���ՋaѲ%���AD��/��QǮ1t�{�b������h�a����/L+��H����m��Y2S$c���.���o�g�Y'��<� �2�/�a�����~/����)���Ǒ��}�����=z���|��k����#���T���|�o������"��]�����������:�ͩ�����y�+�ӥ:�C,+�U�g%��/�Z��k�����v�R}��^�vYoK�Ocpm����x	Wv�[���?q;�z�sm��bu>פ��E��y���4i�]�����:b7���pHW�]�V��H:�cqm�z@zo��E9&��w-�]),,�)�~Ǟp�mق���-z�H(�����l䀳�>;�E���r������ŝ��_m'w�#C@�Ƞ[.�^w�ɝ;2�ߏ��a����L�/�����ϒ�]dѼ�������x���b�s�'��_?��x���q�v�6����kj��͗b�te�̩�9t��?Ǉ�� �.�b��8n�<d2��9x캋q΍���~��D������D�/�u%>s�hh� ?J�O�S�.�ы�#K2��mW���W��w�A��_=���N��Q�}:�[�C������"ve���m��HA{<s����Ƴ�>�x�F�$��.\�Ջ"+�FM#br��k.]b<t���;�lCwW"�0��~��ƽ�E]��o�C�0Q�_���Bwݺ�����W1O��G�/�&p�Ŝax����[3���H)��"0��i����9�vo��� �ۃ.q{��r�da�+P�)l7zQ�H���x�O"�dmٲ��777� s`�Y�KV,Gn^���L���^���ZU"�����z*Q�؀ ��pmw����4Kծ�
'x=�X^(W�5��:��a������[E�K
!�s��um��w�&��u>w�s}򹠉���k?� �U-Z�P����wm��>o]�����q4���+y�k�q'��k�`�����EoO"���l�ڵ%r�$xO,���H.�r���ێ����`���Sl��t�.�la� �rg�{���Ŋ���!��0Q���L
���Y�)n��/֦Z�~�1�>���vά�xq㕸�'I�N�&X����ql���9˫f�o���=�"�Đ�"�t�s�'���*�Ǒs���m_@���u�:~�iB�� &='��F_K��7
yC��}�v�˯{��/�G}�̱&^�/��_��x衇H�N$���%X�r9��+OQ�� "2잣�z*Ta}v��m4�"�8��9L��\�/��Ҵ�{�:��QK���Z
��x<ͱc�F�{��BW[^��7�hID�H��AD��� zZ[� U�����]N�R��L^0��X�ڼy3n��&���8~��
?�=Y��=RE*�Ͽ+�D��l~uj/6��b����PԶb�ctd4J��TXnQ��ha���O"X�����кYf�˷���@ +����/�Gپ:W����*��έ;֮r&?�qe�dl�튦��pe�3ʎ����!5��.��-�V�s��c�}��������h�Q/�_M<��ύ=�=:��uٵ�ѧ�����st��}�L�;~�v���xpB�3��GFGB��/������y|�4i�'�Q�d�R,Z��v~����d&�o�����u�>�,`u�w��\W��H*K����%����Uve��T�1�e^n�^.�V�:��;�n�= ��!�	"��1���s�-�_|����@"w"v�P�?��,.�D�SW�/���?�"1d��=��&r����=�}�H�>�_:O�r	��� ��Q�g�S���ͱ���ͱ<��nc�(�����)z�I�p݋t�/2X<�'��~��1�A��	ۗ�Za�	� 2v/1��Ҙl����C[K+"�{�|��^q����$:��Dn�)r7J�eJwV?��{��a�w1�(�ٲy��7���d�E����~��������Xbv9@���G�J=���s���r�2cx����z��w�~�z��� //񀋾R%|c�3U�r�l���g7@�ھ����;sV)f�)CNnz���)���#�L�<���)L�PiKU4��H˭m۳�ѹ���$J��zh��t*�u]]nm�7�Gt���׹f�?�v������sn0�p�[��k��
:mvN57���w��6]�Q=M1�t��@cc�}�v��Z�>���j��v�w���]�]��<4ڊ7��ѫ�췣��A���<T>x��$�ϡ��Qt�����Σ���a�w���C~~��7ԇ�o>`�\R�[�ީr�a��{����=�������k�g>�q�"zR-N�׼����o�f~sٱc�Qte�B���:U�3�틎b Jpl�
XqW��ĂV�-qzU�TG��Μq�"<~��2J�αD��;� �2mJ���
�h.&"�|�ll�sИ�Đi"�L�s�1'��I�>>}�r<���d�o<A��@�o��fu��+�Q��	V�%n�#B���Ja�%^�"w��-ng�g+Ѣ�L�/2X��?�)~��g<`��M*He<����~:�RU�/�6���a�̙�����?����m���a��;K�~e���;;12<��޾�l?��>22����m�����[�J�N�}������$� �������v�kH�'���s]P�̩ؾ���T��c����x��=]��ݾh�%�ew)o��_�y����/s�f.P�e�%����!�1����;��,(:Fd$�9YX<��р��EG�H��*W��3@�v`H�z<D�j����2��;:��7��8�Ͽ�/50�z�����qO�O�;��=�D͒�X�b�!d��o�8�۰�݀�|Y�`֜2��)zSiX�:�RD��jn�����d]^5_����&D/S�I՟��A̫�p�Ŷ\}���y}���6��n�Kf�:��ɵݵ?R���0*j�؎�x��[��b��ja]�ٵ�%@W}nBف}�Q8m*�M�f�I����Z�Spc�ك%�,Q�Gҹ��y�Br=j������e�<�7��QM�H!l�I.3��֑����ĩ�lۆ���/F�<Y��]��}�@
�����;φd���.��D�>E�&�`2�ijw�`-oG|��#��:�+_�V<@%�1�)�]��P�F"w�HG�Б	��1S)�6/l�"��	�0q��q���3�����g^���A$�L�g����D�υ��>�����{t"���Oĝ_:�tj#"&�� =�m֨��>G}���b�0(�����\�?�v�������;LF~��rK?�����c�!��8H�rWl?S��#�d�w�}�:˙^\l�SJf�J��y�:'/5F1욗�m�z����ܜIy�#,қ��g��HY)2"Sw��H�hJ�_:�,t�Eu�"��p7:B�J�f����բ$j��o]�`#�����+_���l��э�4��Frq�m�r��]����`0���.	�{�[pւ*�~/��ɇ�DF�v� z��M����0����AZ�.� l�����ʅ����XĽ�؞���7�4�흝� �xR�x!��^���|K������̑���w?2�K�m���y�=����-�b��^� ؽ&�r����B�+mǫ��-nW�ý⮺J���7��ۅG�C$��ˌ}�e�U�ե��9=J=��!��~)>_�9C ��z=�}W
୾kR���P�� ��)nW}w�A���!���p}�=X��#��C�m�yM�X�6���^�+W`������ X@��{�5~�>���&$�$���x��}����bpc��/��]X��Eq��R�1����#8v�a��,��h��A���v����c{=��	o&�s�HU�<�������8����;�»���=���s���ƫp�m$r�C0��{��W�},���Us�1ں�l;o��Aר�YR�0�-lW�`��v3�ǅ�$n��>�C���?��?�x�>����	�X��m?�s6U�O�3X��[Lоb�*���Nڶ����x s�O���l۩�>s�RX���))�~*�}xh}��O����;P8�����T{3ޯ��;?��Ҙ���m5���E*���>k��ֱ�'C��x��G��x��ER��׼h�e;����^Bw�C���rѻ�kR:���A{ ���K��acɅ�D�qFuݭ��ӝ�ク�A�1808VQ�����)��+���T{,A�M�6��[o%q;7�w��r>��gb��eVY,�	�u�"x��J[���:8���C+�ϕ���m�I ,�����*�/oRզB��*��+��
�=l�s�@\W��Z�c��OA#�藏�x�]�k����R��q~hb�z����s�}���Ƈ��k������Ֆ.���<���v���n<5i���Sף�	o����x��;�#�(�R t���c�r�Jl۲y���O��91�`����ϸ7fN�vU�Iu *�~���G�"�����1�n�VG�E7w/76��t��ixiWj��$��yY�G��ف��4E�W��۞$�;�dza��}T͜����p��y�F�+V��*�YT>�6�?y9�|�����z���`^�Z�Lႏ�0��~au��r|����y��A�Ω�k�ܙ�{S�ܽ����Ǯ�g���9A����jЈ�@�!l��ޮ���g�F}��da�Cܮ�ٌ�̱�C����x�b�D�ۉ�Mn^.V�Y�yU ��,̞;ǘlw6���/����_�*���K�n��R��~A6�b.�����B�aV �0�\6�R�#����+s��/�����N$�E� r;k�%
�E�����2H���m�AU��^��j�/�x��A�͛7�n@kk+"̚S����iӧ���ݖ�ݿ���e�zItm�b;
�xF��{��XW�)���U�-��]MK�
vَ��\��\m��ޡ�������.w>w-�����j�N9��z����U���p=���-]%Z�<�����{��%$w�]�ﰲ�C��(?��8?T�)
��ڮE�>z���òU+���w���H�S��ą��ٽ�\�T1z$R#`����i���iJ��j�A���ܙ��� �{�H��E71`�xN���_�zA��	^x�EJ�Ι9���3'��A�EL��E��.������������0~ے�>}�e�Ȋ�q�s�?���w�ǖ=�*���u��[d
O����������9�.N�I��1D�w]��n}�D�
ʊ��ԭ��t�#��Y���>h8T}��l��W�7��\�y�P%l�m�gL(q�L<�eq���G$n'�ʔ�)X�r�#q;A�����yg��~�nڌ��D<`"wvo��/9a"w�T��3��3�}��������n��ϑ��9�5�`�5�߇s*���n�Ƀ�6"c�]��+:��^�rk�
R�V��=R� ��u�[�.��T6*��4�2���֭[q��ד������kV��d�U6�]�òXw7#	��6����>"
����Cخ�OO�v�G�J�v(��k���[�n���{�]S�E��.���<����d����Ӫ�j�1���Oa]���＼|�t��X�z�z��x��M����������kצ��B2�=X��r�5�};��,8$�2�`���۴E�b��^�D���2x
�E'!`5s`f����"U|�����5!��#*0��Kw]e�L7�N'e"uL/�3ܵc}��+�?�?����w`����Zw)>zԂ1�ÄΏ]w1θ�1����{�s럊Y�Μ���+R.r���vN�ܙ����uO�����e����m_@y�T16Ψ���	9�Q�-�`��=�s{Б+�D.q�۽G|�f�%��+��I�_2�*q�O~����?Aă��,;j%�V�׺]{@1�a�%�A���P�{/�oي��~�x���7��ϯ�⊄��3I��c,9_��K��9Ckh#ox�a�%�]9C�,<�۲�V-�kud�E$�ù�:�Z�� UPREpa0�� U�%n����rb��0q)n߾};n��F��h�T�X}��q�}�ĸ�×^�*d���&صݵ}�(W)�7�
!���{
x�y��S���S,��K,=�vc[.���?�O���յ=�~T�v�s
1��<R�����������wK���h��~�.���}1�)��Q�x�ßk;;��_O��y�MZO���0�h*�\�)w�	x��~�1V���p�=���g�yfZ���u���M¿��¯Ztw.xw��Eѻ������� Λ�-w�jpp���๽ "�\���x�;"��!w��ڌT����:��پ��f���~m��K1s���X^5��:�]}�|�/�iW�]���q�ݿ��}��b�t���'��L�����-�ണkb^��W6%���[2߼�C��&r>����'�ߨ��Ǐ�ƿ��9��=� �FŴ r;�Q�-a�Os,y�g�e��˿{;�	q�r��H��=��S�����1^�)�ңVb�E�
��w!��,�{���QQ]��;vb���1<D�ネ���/��҄���
ʓ+Z��͈�X�\�c,ކ���'s��˞Wb9\�]Y9��S��S�p��D�D�!�;��.b�ew��\u�*�C��
#�ۣ;0h^����C:Γ|�&ng��MM��&�{�s�ꕡ?�9n�3���) ���%���WJ��rgOm�K+���Gj4�vQ�X�tnõu.V�g�]��s���vR�ڮ��q�\�5Y �X�5�k��ϱ����{�:���Q�X�� ���8]��:�Ee͋�����3�q����	���?���Ac�9��_���-��'?I"��+�$�j1`�_�C�^�*�2_�XY*���!j�WG���8����`A$�>���gb��t�"���J~���xrݥ�W:��:3�����3'�]��>an�/l��p6�˾C�t���ݘ>�	L�~�]����\jY��U�:���8����&r����йq��"��͝x���0kF��u�/�w^i���o�d�g����v��� M �w�	���ߣY�X�ܵ=�)�רϼ�;wY�M�nbF��=��X� ��E�xꩧ���?��ILl�w����8z5r��2� �h�{��+W�z�B�ܶ�>�a�.�X`���c$[�az$�3�6�r	�a�y;�+���e�.c�.�G�xb������씙�x���8� 	܉�gJ���&�cR��vS�΅�{�,n���1��Q0� JO��]�ߵkn��8@	kbl����eK�?��sW@���S�ڮ��U��.�c���(���mE�;��u�rY.��\H�k�����>j�e�rx;Q]�5�W��<����|���õ]�S�Br���N�{��יl�r_�k�k۪��~���z:7�v�mM<n�`hB�xϘ;>.�WaǶ�x�OBwW7"Vp������~�� R���ɞ���Ќ%cv���@�s�A;h�P^NUx
t֢r�Է�ȝ ��g>���Ӆ1�ߘ`���R/ngl�kƙ�����9|dE����M�ó����p�&��X��-]���'�{�104�+����8��cj�9d_}�)����A�'SD����������_�-e�v�{�c|�M��앳g�^oIE)~u�U���P{&_=�Dl�ҧ|�l�͹5:z[;g�l��=�)V�Q�M1��Q���+_(�Ϳ�U�X��K�y����'q;1n��+����)E��#� Lrrs�꘣����mނ�u ����J>��q�|�%�P�з1��8���ce)^���9� r���]vr�r�R���gWO��{�A"����H{ήF[��
z�Da�������gx�D;0D#�L����L�~�uס���D��"k���/(p-�/lO�k�R���{�`����v�8�7�\�\7�MC�?V�*�v�=�������r]���vm7�";��c��O]Ѧ����'�ZW��D�*�v�8[��v�1V��5���_
�����rm�r����޸��������L�]ۭ�T��{Ͷ���X���,��o��7��W�� b����pr�����'��cB��H񜏴��ί��;�DvPR�6mA���Õ!�ҝ.�`�J���<�㧵a�4�R�� ʅ[�G�sᘜ��E��i��3����y���վ�3D���L����Sgg&~�KS[7.�����s��G�����Oo�<>y��1�qř��__x[�!�XHw�{�:��44w��c\3w����+1db"w�;1`���^y�y�� b|,+b�u����5�s�����]��QG}vc��Y��yD�����yղ^x��?��c��d&V����?0KA�)�:'��QZԄ-߄��vD�����z��^p����t��z�)rg�Ǉ������ +�1�S�.�ܭџ�������a�5�V��3`w�("Q���HkN(�FoK�ہAZ���a�{�R��^0]b!��6��ۇ�n��x%�X�1�kN8ť%�S���<�/���F��õ��u�z�׵�-���k�������k�S�<v�sޖ�<�-��}S|��z��{��K�%ӵ�%�������1�]U�e~��:�P�v�?��%lZ)���j��3�r�ǰ�c����M�����X�n���pL�<�(<��X�k�5�"m�[W��T���=R����]܍���+6�vv`m�4�v�H_8�h<���M�HGq;�	|�������&����|�[�����Q2m�����w`�o���?�:84�������ŧNX������;�$l��+ b#]E���.�x������������^����B�{��?��"w�����v.?s��A�r�0�;W�gyC/S,[�p�����G}VO���W��I�y*��/����^���8����)S��أ1��AD|�5��<�l4���w��@?"���q�=����sN���W4�:Y���smAX�ȷ�����2��]��|��34���B�Φ�ZP�>��*� H�N�-�Y(i�/a�5p�/���'�C�HT?>�;���� �X`�,?zj�,v����k����*��"Xq���W)P�M�.�]��1����f���
a���K�.W��EBre]���SW��)�v�I�Tۚ���~�Ӑ�Õby(����{i����.���������/��5g�z��q�qlT}ڒ���Y�ӵ=�-���En�:nN!��������?sHe�}
����_��)����g��+�Z�W^��6� ���ى�o��pfX�bE܂=�h��v��|�}ݓ��<`��BW���̕!,xծ�a��Y�j��KKj���Fx �x3��"?��7����^w�!��^��i�}�~�Y3
���+Gg��ߥ|�E�_�9���#�����ǿ��9�u��׿�S���Ͽ��J$�J��ܙ���?�3�[�Lܾ��@�q���8ƿ����_�W�6n���'��=1�m�y��p�G�� ��sN��[��������b���AK䞌Q���1�<_:��㙻����+$n'���.\��V�]H�B�(ؽLeM5�++���رu��B��oܸ�����'>�+?���x���c3Ɗ$t7G~s��P�=����B�nc�t����nDB��|"m���>�����T��]���],a{��)nD��ہ!�H��g"�[o�;v� A��}�Vc�Ն����ο�o&�z��,zU���F=����\݀-Z�k��O��X-�w�G!(�ۊ�w��ڽ;TN�\~����vI�5+� 
�ݮ����v�}7߹�Ϣ�PO~����ӵ��٫�ݿk����D�&��#�Q��r��9]�=�7�nWQ��nh�����k����O�;m��ֶ�����:��D��r\��/aۖ-��W�����)< �{��[n1��.\�Dw����@�S����,(v�nP�vrgx�ۙ+���]��� U�`��5�<� j���wFDt���_?o�9|w7ο����KQ1۟ӯ!2]�!r�D��o]tJL�v�??�g��·�4�h_��9������ĥ1�[���sNZ�g^�"v�������W�~�������˱���ҏ�� ���19�?��i��.S{����^�������xn����>���������y���A��5s���9��]�����}��>K�X<W��!�W .�.y����7�����o��"��+���Ea����� ����^���*����qp��_�~�z��OW>0]���cTc,�w��	Bw�����\����N��������qpp���KQD��X���Ob��~&��t{A�[�%ƈhc,1�رDA�F�*R�(W����3�3󴙝�{��7��vg�y�;�3�;��g>��/r��Y4����Gk�z��3�m���D�!�;��;(��[}<����]������#M�x��܌+��o��&���AA����&O@�JU��k{x� m�iT�vYt*��U�f��W�;"DU�tEq�{��vS�S'��t`����)��6<��3Ko���.t�6�v(�T��\��퐘k�鬔�&��YyU��ۿL[�m�m�.l]�\_�x�]�FHȵ��ݳ��,��b���l7�!]�w���~�v����E:~ŵ����د�|��P��CǍÐa���/��7���ƍq��c��0`@�N�����䞏7[�҉�M˝Nuq����w��}o�����c�@D�3{<n��r^�n����;-'�ic���S�%�<��Ex��u r� ��~��^@G�9��w�#��_�btt��$�N"��j����{yp��������^<��ۗ����v6��7�y��l��������xnX�+N�Օ���l��H�.%��p R,�ꆶ9�W�woq��	����#���d�۳I �����ۖ1ց@A�\Qa	����� "3�s�c�ƖM�-�{cC#"���V�����=Ǝ�qy*E��ZNl"w��S7���\���C�k���y'w�џ���&�|��>-��V݁H.$p'��>!�7m l1{�����=| ��*���&���T�td�(=Y��]xW_}5�.]
�BiY�0jj��>����G.�X��ڮ�s�k;08m�fS�ڮ��%��,'k]��-�C̵]��H�Y����/���W���_D�����Z�ݐ&)��!L3M��w\���"��W{l�!�w���&����1y����\��,��]����	����sg���I;n��Ǔ���VD4V�Ze%���{uuu���{'��dw��g�����*���IX	.�19qr߻c#����ɑ� �����<��0��W܏�ߙ�o�41�<�J��𒯑�=�a_u���/l�]h�M�?؆�-X����|���<H�DaN�]~�"�Da��{~s:��0,�y�����<��;?����)������'�=+��gcH�*�f�߇杭�{{W?�����v�{{&F}�T�.Y$3��?����џ��;���>#ǎvrbADfa�i����?���>짛ֈ����㷿�-n��&6,�&S�ɾ�����!�]Ï���|��~"w��.�
�ڠ�fȮ�t��}��avM+]Mrd"��Ed̩pz�.47�(..R����RT�;KL����{�	�ˁ���N�"V��9s]�����3π �0pH�%n/.QݱbumG\�k��?v���ѩ��K+ί���?T���	�u����$mw)�e�q"7]��<�S�rrf)T}[��W����M�>��m�D���
R<�45v�g�sm���ziں�+�,~�v�_��4B�X\�����ƦG��͵]Z��S��Ը�ێ�rLr?�^��.�e�sl�~}���V��.���������zp����ҥK�D��{=���C�+a%'��iz��;�`4w/�;��P�M���7�Z:�А 2Eiq!n��]��l�Մ�\z>ٸ��p៟Ƨ[�qŷf#�ɛ��o��1�����?>޸�W����L�~�����O�>:j�U�v���,�8L�~�s��G_>2m�<�������ث¹]fQ����������4s;g7=����Q>������� �Ì�B4�Xg��\$�ci̱��aaH5�*�ܨ�:�������֭�DM[�nM���}�����Љn� ��:�o�cF������[�|sn�m�Բe�\t�E����z�gb��t5�w}�������K�n��lJuC{���X���1u����nv!�	܉�b����$�Nܮs`p���v�J+n�=Q�i�hdCRJ�}y�z�X�d	"]�Ub��I���y���T���n��b,z��]�Mh����µ]GZ]�q{j]�݆Fd�I.ں�Z��<-�B1��kE��Ivmw7��Ov?_e_T�3|lhb����n��˓��������'v�Q���4h��cCwA��k; �d"n7S�F]�׺�?w�˖�uΝ��C�7��sO?�O>��ǲeˬ�����Z˝+Ӊ�L�ٽ��"ww���Vr������%r�Vm\�JrP��p0򷵥'؏���@q��\�\�����c��:��_A��Ҩ�+;��Oִ�'�����̺���3�x�۸mθr!��4�Hmi �<2�<�*�v@q����q�϶�����K���]:� ��P]^��{�[�>y���3�r��B���:�F}֑5�T=߼y3~��`��� �h���4� A�ݰ��w4�lڌ�����͔� �Y�f�%r_�`z��l�fK]�����sK���!<j��߰ȝ5���S74#uC}������l݈ne��s/�DI$�@YC��!�v�C�-h�PEA;�����ݝN>y��u��с!R���Һ뮻�׿��}G�א���e*	*��bHص�PE���zi��S+a�BaE�nǭt���.	���Ʈn]Pn�h��3K�$��݀# ��CX�n9nGB;S�N�{?K����Z�ݐfW��~��V��]�u���c�������.�3"q�X5��u��<������e���Ƶ]]W�7� �y<��د-l�	�v�S�<�?Ye	ݛ��@^�����?L�Ά�tB)�DO�c���c�qc�V�����}���7��NN�D�V��'����L!A%'�t���1��P��e?�H-�(n���۫��܃�.:��v�m��L#��+��B��D�?��c��z�r��Žۿ���p��`1��l�?�����n�%�qh-��t.+A�cf�&4�jci��^�f(�a�<j�Y7곎l�'򼮮���Z�
�;������nn!� :lԍ�_����a�G�� �X�r%.��b�p��֭��N�-uE_c,��uJ[�S��k�����;����Z�%n���k���[[Zp\�}xd�G��@w"+`����w�y��$��^�Ђ��U�A������ rǁ!�.�'���w�	��W�>?e�u7�������hFo��k{�m�|������kgֈ[���Z/���N�̉����e�:���Vl�퐦vm��k���ѵ5�.�C�/	���.W�|���D/L�vm�֋�������F�0v��7+��!��)��=f�� �D+$�C��u�)qm�n#gk:�(�+�p/���uس{7�\�:'�|UUU��l�^��QM�.�;Ye�ݳð���_YܮzP'r;3r	���#����Α�~�&|R�����@�䞧��Iq�ͪM;p���]�>�
zq�So��O�u��v���g7?�K�z=������Z`ۮF�m���v��Ȝq�a�tH�8�~�1��O��BHO��F�ƈ�jD>s��B4�oEqI��v�qo����υ��]��T#�,�9�"b�z��ЀK/�+V� A�Qٽ�5�s�U � :&E��7�R�寿E�X�/o��6���J\s�5�ԩSƅ���S�[ߠ1�Bd����o�g޵ݒOp"w����ꆼ�ݳfx���3L�7�6 A$
	܉����B4�ׅ$���h��"r���u�Ar`�|�ҥ�+���/-���.hƎ��Çjߏյ=�`=�ފ!a�vM:[����sm��wm��Iڎ=Ů��[�tN�,u��v~}LCޞ��r�յ]��1qmwo�5�6е��%��$vg�ܿFH���Ǖ���<�=V���|��Cjd W]��e[7���eC>�	s�X���%ر=wExDb��~*++q��
��Չ��.?G%a��5�]��I,�����E�vM�ud��T�ߖ�V̮iţ�)�@Db�j܋3�\��ߙ�o�4Qy��'�Ꮛ_���l�����Z���|i�(��Ó��b��:q���IY_v�˵���<�
���; �|�{�tٻm�EQG|V!�9V<�CY؞ͣ>G#�u���V̟?˖-AxQXT�1��Ð�Җ$� RKe��8d0���������_�~/�"�N0�<�%��X�)���s����t5C[����n	�պ����]/��lDeY��K�=�Ty&2N�J6 ��]#nW\�ei�A9)�� /�����_Q�9�2�-�� ��{�=\}��طoBG��}-煲N�a�c�#�L���M��ڮ���յҙ�S��.'~�vY��N���r[9N?�v���k���q�֬G������ns>����s����1Y��F�����`�ُ�8��v�����NM�6����k���o��$M3�s
��	m<�ùI!�k;߯rc���v�y��E�~���e������Ժ�%�[n����8餓2��ʤ���ا��KXy9�&�9�s�FU��{[�폃���;6��>C��r�%"1lÅ~m؆k�;���������%���_v7�� ���S��?��u��~~�Q��YG'����p������@pl�f4�<6Ɗ�����{{dZH�%�#=�C/�v�G8�ٱF}�F����7�|3�~�i�=z�Ąi�ѹ�ADn�~#}�����^{�?�
���F�����?�AJF��l�%�"�0�{���0Tc,�����}�5B� ˴����B���]7Z3�---8�_�1� �gFu�w�(..SE>	*G�n'�
݄��P��+Bw;	%%�\�d�w�JG���?��S\xᅨ��AȰc�9/5B��-l,n�,��hPvM��kD�B;,��mՋ��0Uq�:gx��Fl��.x� %v�}��#t��CS
\��vnx40M��Fb���JqM�(���>_Av��fx��vS�8�x"�;���k�C��]=���}�8�Lӣ���M����ekjL���4�6P�p+����\+��ҝ'����,"W�>m���ۇ��L�y��'}۶RҊan��Ȯ]�bڴi�gR��{&7_���M���9NL��ΰ�m��=t��C2�����G�������������>߉�f7�;�F� ��'����jވ�u�L����V�قo��;6m�� �i5�h���%���vχ�s{AD��ݣ>g�Η,���~.A�(*.��q�bȈ�q��� ����i������x�o��~*"*��s�U3��׿��H]&�ꊉcI���b�e�4�3�3_#�k���=,n?�u�(.�RݐՀ�vlƤ~C��f���Cw"�[BC�������$�Tn�AA���������ޮKT%!I�#WE�۶m��_��>�!ӧ?��D�>������ 8?�����+K�P�v��FT�Jm�\�����R��.^=��r����hp����'͵]3��$��.Ϋ���.']���x��έ���F��ڵ���p��#5N�硉=�k��=L�6�����!hc4u}k>s6�����n�/�{]R��n��r>]����������?�^y���	6���_�?��=ztƓK��MhɎ�C:r���eX�����$�=�nPv��������=�`�_;iղ�'֚xl��v#������A0��H��J�9|��˯�(O���}~vڌ�����m�Z�� �M�ʲ�Z6����1��=���uuC}�0�{{�G}Nv�|��O��nA�`B�#�MF��rA����Cѫoo���ױ���	l�g��>g�dS�0�uE[���ٵ��Y�/,������eq�m�řbEj�Q]ܹ��=�_�&���FSK�o�%����<����F�����'�d��B;!%&��\<U��v��&��T*�E�HU�����%}��G ���b��2	����M���GK���DU&��O\N$BUt*�����{��.�vy]ൎ^�=��J�N��Ĕ"�vqY�g�r$ߵ���MH����'���ihb������n�c��#i?T���i��I����*�V�i�Mb���~m�ѵ]����E��~f�6��5�.�6��q�/,,�Ga���x�n����ĒV5559�tJ�o_G�?�IX�N�^Cڂv1iŹ4pN�m'�X]��n_��zÊ�ɑ� �H.e�E "��9n0�z�(.
!�a?��~{�;yr�}����w>��Ͻ� \f�ۋ���(f�X��~�v�n��e�{ �v��%��k��T�ԓ�_:����K���,�F��)*.�������A�Iy��8*���������TK \��0w�\TVVb����f^�.��cYF��g���Y�U+��c��p}P�D����h϶)�麵{���hiiŜ�xtU�獈�@w"cݫM������so�%���۩]NT���;���v_��Ƽ�G:D2*���~X̛7���:����O�6e�ʴ�̵]'�T��d����ku~3�O��P�nq+�gXCTl���4�^+���k��rL�޵=��Aq`�v�ێ�ą��ŋ��vIvm��|�l����x�ͮ����R_[ǆ܆#p���"�,��(�caߐ��X\�}���F2�����~��{Ӛ���ǋ�΅�;s�}[l��4ͱf۽D��gajڨ󙦦/ݱyC���F�z��y?�>^^�b���ͦM���n��&TUU�=�ēM	-�|˝[��uN�;2D��#��B�;a�qqg�!�-���-�!� �e� "{�2������~���־��_��g�O���;q�5b�*� x�(D��uV�Ppo�e)�nX����������9�5�l��������+�w�^O��}0��)V�pݪ5 � 򛰛{���kؾu¦���]v�5��ȑ#�R�Γ�Z��1�S7����j��z!���L��Q���(Ϧ�1�3_/�\ܛ�o���C��gt3;��u$����P��%�Jr�(��]v`pU�DU���˽��a���D#��)�J@�}	����ǳ�>��a����b��C�?��ƵP��V�4��k�j��rm�Ϥ�[��Z�fZ,��i��fDTۢpZ�'��q����������a;�z��Wi�Z��1��%ϵ��A�凧��ڮo#n� Br;ص]8^4}����d�m���9 �p�2�e;�aM�_ &�v��-lcbE�cf�!Æb�#��k�.c�ʕ�ꪫ,����ҬL4Ų�d������pn�Vq;2���&����U�ZN���܌jM,Y� �H�:�� ��`�!��eg�Si*0����7.�>X���{���A.%��z!g�U$	��q�[���fXќ۽��M�k��HG�q�����K����&Z� ��_�;�c�YX���x��w��A0�o�nc1�{���3*f��Z"_���	9c,�nh8}�źaA�^X�&:����{,.�������Z����i�[Y�6�G[a�ց�NJ��0�!7Y�sm��W~�����;0���]~�h�"<��� ��=�0q�TTt�}���sj+
���?�y�6� ���z�`��5��b�J� X�����{	x�������v�^��˵J�����!��4Vד�Hk����"i�]p�v1�3/�sh�Eqm���nv��&����>֔��v�җ�3�/��؅�H'n�쳺����Wq�VH.k^Bri_�ɵ�	)E�����������&��u�X9S��h]
Є;��j��~�C���g�Λo� l�o����o������V�]A�����'w;a���OVX�GΕA�����5����Q=o? � �HU];� ��3aD,��l�����
L�~ӏO����p_�y{5��`1�[@���-�[ߊ�bo�vOq��n�������Y;��4��&�͑���T/��ڙ�}Æ �h�C� �`9={��/��]�;A�O?�W\q�U7���["����YK���	axG����>�uP�O�fh/�]/�k��������Q3tD�]7liه��U �X �;�v���;�P\\�80��0J�цԹ0x����줔����7a�QPA�?�������`��gب�=�P빌�&?Ln�v��+z��"r�5��e`!�03�mլc�iU\�*�U�OMԵ]I{��)n�c������ ^v�T���P����sC3���څ��<vg�;���S>y_0����Wi�{6���p޹��cP���\��(m��b�v�uyz�}�\�q�ǲ�󰦍�/���.��v����h���y��&��)'c�C��Ë-�g�X�x���p��M������X�s���WF�I����	���'��_7Q�2�ޮ��<����Xmt����	� �Օ "���/=��r_�^*��~�U|q�!	�u�o಻�����9�_!�v����ݯf�<��a�X;�cy���bzs,F*�:�%z�g�---�7o�5:A0��	� B�KeW{�|��J|���q�f!r���~�_=.��2���h�'�j�:c,�t56��{�uW3�E=|%��,
�M� �K��y���5�o��
	܉�rx�"4֭��9�ǽ�ׅ� ��B!���/�&�d�v'Q��b'���T6ٔ�Je���>��JR��O_8й��fi90�H�k{���sr3Sjc��T���V�_����R�v�vN��S{
۵Bx9&/�vS�3m��ܼ��y�rm7�MWT�l�\�5면K�k;?_$��������M���=���.�^��|e��ej�U�6
�Fخ�l/Z]���Q/�ר�Muy~}��L)�aÇ�����=�֭Y"�a���7ߌ�}�b֬Y9%fO�?��gw�92�U���a�����JT����M{vcVmw<���AD��Mw��$cj{㑫���Υ�u�
C��W_ŉ�G&�ρ�m��g�i�2��Q\��h	���~#?�$Q{ac,�v���˵C��fMܞ��]2�H���a�X�� ]�`⴩��C� ����6u�X���o��M�� ���z
}���~�m�,���d�Zy�K�1_?T�^�B�z�-~o3�a����m��R3�����Ë�⣂�8��	܉�Q2P[���v9)�9� �P����ON9mb*�$��l����[���+���$��kpđ�QTT��g���#�Dm��H��R#Ƅ���sm�*��
���ڮVUQ�:�-4��5XO������{��n��bqmW�����׳���@\�<�}AZ/����^��8_���}Í]�A�	�vV����;!%۵]����Rn^�z#��<��~�w��q��Z��i#�Y��&���� �'&n�WL�qη��7^}�~�_օ.���$��W_���jv�aJ̞���_L�#wHE�����:���î�+����c�As����-AA�0��'��Bh�O�)�nF���!�a登~u*�L�P?���;�?����A�9a���%%%��ݯ~�{�"w�+�׫n�-j��Q��G2�?���X�h�1pH-�<�:^	� "^z��Y_<��&6|�q��Z�?�r�)Y#f��|-�U!��0v;�n�U3O+����|�P#l����u�����mj���xj� �`�U�6N�5�I��(��B�D�΁�����5�톒��$l�Da���6�}Ē�
����f̝;�V��߰cm��0t���c�ۃ���E �-�Ř�����R[�4l����g��=��i|���W��!l�
�5b{h�Ŗ��(�e����Js��d��r;թ\��@r]��J� ������몾��5�h�Ь��.�ؕ�Hڷ�Ⱦ-�$��G��c53�5r��Ҿ�k; ��S�=�,+�k�܋�Y��6r<��uOӹ���s5'l��n��B폩ӧa���X��Cصs��eϞ=���Kq뭷b��Y�tJv�A�K�#������D�)
܅�F�~P����bz�f<�P� �H��]:�'L����:�H̹��W��n�/n�TZ��.:3�M��u���׮Z����QAxQ۽��ִ_O)5�"��aa�S�7�
�J�0�l0_Cd$Cl�|�&z_�t)~��߁ ���0~�D�� �H�eҌ#ѫ_K�~`��3ƚ?�e�u�Gvx1{���ͧ7�r�u4Y\ݐ��}��H�P7��j�e���Ba�g��}�z��Z�M��&�Cw"-��Tk�����E�CH���%�x'�{Ȃ7�t%���G���KP�X����H���bd
��0t��� �랬嗔�b`� ���a�⛖�Q�?�ٽ-��	��HZO�v��TC��=�h��k*57�D����ؿ�}�[���գ����O���ʳE&�޵׮c�cj�=kk@umwE�{ڗ�a���K����߷�ِe�564�M�W��5=����F��~'>]�Z]��צּ0M���D�s��0;����U���U�3|P�T���X�u�YW�ҲNڮ��ZYe���M\���G+?�ϧ���M��YF����8p� �����J�~���?A�,u�l�|+��mFqQ�FA�?ނ�cžt��[���wV�E�(�;���G��Wb�σE��ߊ� ���%���v�܉y���n@EEE\	�lJh�ۇ�}��;~���]N\y&�"�v{�A�V�����$�l�;{�P�S�k�� � �g�%/��F�ICTD:8lH<tE����vљ����}���p�Ջ�}W��îa'tى憐֭������a�h�ŋ����џ�ڡ"|w��:q{���td����?�F�ۿ�����=�,b�
AD�8����y��W�4�������+��m�݆!C�䬘=�X|�P���B�w�f�ꃦ��]�ٮ!��aj�n<�;1�!����H��D�@�
*���d�ށA�k��n��?I���ʄV�E���]w݅%K� ��d�޽���*SɶL�{2�_;|(ƌ;���'�k;;�*�wCIiI�"4�N�e��rϙ��_� �S����.�T�B;/�mX6��}�7�ك�޽�]ۃ��v���J�]�d�oݏ>5���((�՘���]9������_d���	/L�Ɔ~}tbg��4�bIl__Wg���^]-��S�)��/�bl��#ܚ9��(�����͐c��ئ��������C���؎���L�|�p���6nBE������n�m�{N�nY�2������6Kx����X\��I��`wӰ���}Vs\��KwR4\�;�n5��PVV�����0�e)��04��x��3q��ч8}��*����I�o3v�axoŻx�ɧ�^?����gɍL�ѿ���vg�e�~c���[�+�W\Uȟ.��L�!��;2��aDqd�v�MV(�*�mD���=E������"�:��Ž���[� "�`�֘�Wv.��~x�%%"�L:d ��,Tt���x������Ƅ����k��G��V�ͱ��а�><�s��X�C4�rM�x�,YԮ�*Y�ꅆv�]L��U��m߾���<\"�Xl�|^��Z��,w�	2iX���LpسOo��|����n�d�]u�X��e�k�km��;�2��Lo�L.����2�*̐^&ם��1Xk��'̌���5�F ��ٹ;c۞��z}Scfn�ϥc~��a��V���~߰ߏ�]�`��ڙ�ms�)�477c�ܹ�1ssOTp��Qk�"FDN�j-���Y茱���a�F��,cYm۬�a[[�qs���ȝ���7������xe������H9�*t�T��B,I*>A�&�D����������O&D���O~��SOY�d���2��n�Z~&�=�峡���:��(�E��X����c5TH��G�*����l_n����qS6��N����[�.����X�P!��k�5Br� V'�5�y�27��{Q��l��]#�Ո��mUq���`78�Ķ�J
�#M�־1EVH�*h��l�i�_�|�Y�)��~������w�I2~?Ҭ����\w�v�s3���`��=�]��=���~h����y��^�$���qG�Q�8Ӵ7}�/��|S\\�OT�e���i����#�%;��ISnc���k^�	� ��,��ذ�l�N���-Y9�h�=J;gy�1���w���.&��]���lʄI1�v��B�ؾ^��I��=oǐ	���駟F���q���	�t��y��G��ud��
?
\A;����+g�A3�����ĥƑ��ef״����HA��{{u�OO�x��'�w�0w��M�����/�:�e� ������W��qC�&�σ�]�_��8���B��v*KЩiL�s{s,�^�덱B��]�:���t|�TW;�IW/}$k9LTĜ3W�\�Daۖ�ۛ�23�Eii�e��X#�dj�������f�u*���G�g�^q��Ď��A�X����򙸞�w�v����3��3��m�}��]*Щsfn���3���Ϸ�oMb7t��w��R�<}dr�3S��=����2Qr�g��[6m�[�,�jxe�J���"S���]���X��2�K���u��u�]g-+��l�%��X��#����s~���ڡ�o�Ż�[�Y[{h�nئwp�k�e�{��z�&���AScސ��H),IUޜH��@IX�C�n�!u�*Q�0�'�d���|�Nt���{��L&v��R٭�=];�`Pq{�GS��&� ��풟��<���j�Zi�-�V����}Z�US�S'浻�������eA��>�~==]�u�$6��#�0e���i�5qX�N��%�E������� ��ɭ���&����:�t�{C�F������['nw�<r�r��M �k��e�x�����k|,��&����3&C�a�۵]\VP�vmD�[�ӝF$�ۛѶ��t6��Yj����]�������K��� ���I'���	(��R*�QX������k?x7w�}~�A'iIJ��q:'w>QŦ�ݱ#������@A�\s�QZ\��}iJ�y�����v+^�p�H.G���/9她/n�TZ��.>3aq�_��~{�S��A����;Z	�)Vpq�X7�넺�ew�ڡ�9#���#֚#��_�`^}�U�K�^=1y�4K�NA�O�~�u�X��˨�1�"r��^z	7�|3~�_8f���w�Z��1�>bu;c,�f���G�cq5C�^h_��uB^��F�=� [����	܉�2���cKR�%��$����5Ġ���/Dsqg$C(K�Tӓ���m�p�UW���D~2pH-�O���Im	���v��@�v�8TO0�vA���,G#�׵ݐ���SbJе�#vOq�S�]��ͥ��JJ�cS�·�Sd�$�t��5�a����(Z��h��R��NX]/����@[������~�ˎ�9���.���m"��uN�Y7eWn���gB��M�bM�;8��X>�F�,���pmW�1�x�y���Csޓ��n'�>������d�x��+�"<�ȗO?�C��ǞH�]�D���_=jjj0f̘�K@%�_,��m��g�5��p���>䄕��Ҹ��!A�nZ����'��e;��膃$�!� 8���s��R�S��}Q� w��8��w㳺= "9?a8���i(.JNq�݄2��d#e%EXx��0eTb���ث���� ���[�ƺu(..�4�ҏ�vjwj��zc,�v(�<j��kH�v���&���x�KWmQ~�p�B<��� 򗡇���G��� "�uꄙsfa��w�����O-Z�A���NK��=�����u�.���P�������=�wq���ᑞE���!r�[Bw� k�s(Vn��?���D�8�O!wĞ���U�%IŻ1�ɩ���DU���:�)1��7ʇ9��Y�D�Q�~�>ij5C��,�  ��IDATE�c%���t���m��M�!�k�( ���%����Jۣ��C����DD�o�s�ļv�IrmW���5b{@���ĵ]#:�����.��u>��.�vx�3�?ޟ����	�qe>֥�!]����ݞ�)���daz� ���y�S�lϛ>4�A�gbqm�۸=z�$�1#;�|�̵]�����i��j��1I�t�y	���|�Ï8�z��C�?�];w��/��ك+����z+z��v1{2Z�����ב���V�k'�����i'�L+Q��3��� 9�7�ٍY�Uxv-�EA����q��p��ӧ�^~6N��/�ݴA$���q���'n_�����g����"�`�F��[}"���+����� ���2��%�EL��b�Y������ uCK���b@���^�d��1_�k�̵���n��0�	GNA�� � �l���;~��{��W�ak+��㦛n�D�'NLj�'���xbvtK�1V�=�1_;�k�|��wqgӬ�ad�g�-d�#uD�^��a�uÑ���Q���������H	�@m�s'I��P�T�D����$��\��R`�DO:����J�KP=��� ���z�t��߰��������h-��#ҏ�o�u/�{S��TH�)��2=�k�6��N챴���J(�vm��]�j�H�k��/�����{�csmOf쎰�;f��� �C�I�.�9�gݔ�]+$��3��O�/̔��v��)����;�%'������,S�G�G���q��/�v�D]������v~"yq����o�~��O~�G��0>��#��ڵk��1���Z����U̞H߱����s�{�g{��9	+{>Y�n�������`��d���ɨ��)$�G)Qe%��l@U��knAA�l�~��M��[�2L?�6�<#j�-��s�=��-�AD|�2}4n���(%���~Z��pÃ/��0���f1�����g��v����@D0Nl?���5���4\���7�*�������ꆱ�cE7��MKU=1��R�ߺu�Q��A�Tv�)3��sEgAD��w@w����K�M�Xy�޽{q��W�[n���B�k���1�^bu;�n�W3�녎������a{�������=�=�
O���!�Bw"%̮-@s]�%6qSEE1&�ć����tI*��#r�%���ǻ�T;0����~�G���0i���;F�۳յ]�Ih�*}�u@�>��6&�=L9v����R���O������f=3��.
�����c2ܵݾ���2��ɢ�d���䷕�@�]��]����b���rkn���n�����7ͨm"W���M�umW��T��G�GD�R<�,?�k���L.ve���K��w��ƞVVV��}�,���X�or��7�.]��o�?��O�"`O��=�>�ik��&��s¯���k �C�V^.�,Y��c"{������d��� 	�YA��-X��A���z�����s0�`�L��貳p��Eh�Gn]+_�9��)I��c�'7/��/�D6RԾ�w��T?aXB�0�>��	"8}��@����D�VX�c��n(
��ڡW�PW+t_�)7[�^��$ې*��%Rglhh���۶m�1�M<�:�� "[�ܥǜ8o/{֮�_lܸ���x�(//�j1{�5����uR�>��Y����.����P�V����C]���Yvrg��ףW�A��H�?"$p'�NuyƮ�(��'�
�$�޽]��RD��4p�����3������˗[_�A��D�0b�(�9�0�QX�\��sn���1j��]����b�T��+1�ѵ��	����n@j�^�ve�힀�n��`
�A�������]���]d#���PHn�o��_sG�rw��o~�!�)��y��/����y�@\�1�VL\�@2]ەs�&�hm����g�a���?������~��1t�P|�_L��=}�2�_[_G�KZE^��ܽ\�CQ�U���;KV��mڱcz��[� � x��9W/£W��1���3u�@,��k$r'���	G`��N�����mg�u�X��H���-?�2�L�P?�=�<��δ�=h�m��B�l�%��5D^���������=�\�H�ks��MV-0���u���_o����?�LĠ�C@A��:�����xD~��o�w��.����@&�&Y��CG,�X&���y��puC��F�Kg���j��Ԋ۵uC� kF��x���Cw"����;�@�v�Ђ�I*�{�_�� @�J&UB�t͗H[�l�W\���&�CaQ!&9���h�	.l�V�v�V�_/m�Jb�B1E��d*�r+Ź��@�J�ib7����{�[�>���z+�k���pcu�[:�]��5�۩�kYo��ڕxwve��m�
kyvu�|��z��@����Sb�F;חt�"ޭ+ƙ�k�!F�x2=����$$�nK�k��I4�����I�C9~#��H���y8�<߯���=� ��TU��S��%�h���x#�܆��G2g�s�|�	�۷D~����Ϸ�<�0�F�t;+��G��qd�q�Ǣ������n���.�z������<�$��d������莃ts
A!��iκ�,�曨��=�<L��׋����=h��	���'L���Iж��-��Z�1��f#L�~�_���1:�~n_����9�I����~�8�s s,�Q����'n��V�0�9#�fX:�A�~�����'�����S����� � �����Cѥ��zeZ[�!�x���1r�H�~��I�󤻖�nc,��ϲ1�+n?��!m�PW;�	����>C����.$p'���>E�'�u(.�$�4.�k{t����T����&��xS�p``B�y��aÆ ���8��е[%75",n��3����Z y���\�j"���b��^��ٱ{�'ku�5�ve�FDx�!n׶�b�tm��'2As^���B;S�W���-�� ��Ϲv�]�֟(qn����Y�(U����	���τ���t��qr��#��}�����T߯f�����g��O2�c͞��x�����ԉ���J�y"�h��K�Qo�ќg4Ǯ��nu%�@|��7D�������97��m�sy��U8��YX��;��Ï@���͸��p�M7�gϞ)K@%Ý!��b�Y���ܰ��-p����{$��u����&�tɪ�s/q{$YU(��76����z�Oi�A� Be��F�v���ǵ�B���@��8�O���5��ذu���N��_?.)}����;�!�j܋l�����/��3�$��#K�#q;A�HQ�@?s���B�ݰ@��۽=h��5ȂS/�oO�x=u�D�x�p�w��/��}��(�T� ��0��'Oć+�Î�;@��^XSS�)S��]̞�ZbPc,C��o�E[�S7�����.���1ƒj�^�?����E��Q�����B�$p'�F��$7�x;���Cz%���T���T�k�_�*�O�%��ξ n��v��� �^}�`�Q�PT�������\��`RC������Q��$�?�صB�@m��99��V�]ۡ�k������	��i��p4��r����	��i=M[�-�Q�m���@
\۹�=ۄ?y�Fÿ_g����.�F���}�����u#��?��ǀ�������G��ˊ�՗�[�����#�"�>F�;�#��3�6����N���E8���ťK��g�"?ظq#���j,X��r���w�lrd0�O®u��Wwq�'��d�=Y%	��뢦��,�]{I�NA�lܶ�]�7<q�7ѽK�@��Wn�!^X�6+�ܯ��9l޾�	���_�1�<sfR�{j�G����b_�d#l}�K�9��'�Ͽ��?�y�.%I�s��=��������O�.�]���b����k�D�X�f��k9p ;��Dj8�GL����� � ::�7�I���O�n�Z�3x������?����O�=��X�K��SJ�5/����NB����v[�λ��5C/w������{0���]K5C"	܉�q\�����J�*T��IHRQ�T��y&���Ɠ�>�{�9,\�D�0b�!3~w�D��������3#?���L�k�����ʵ]��K,�YN���t[��mL����k��[�,�6�yU�z,�G�r�:�k��;�>V����.��z�/.��D�y9�K�����	��!��)��=�k�sN	Я���C�ε]�&�6�va>�yB#���qΝ�r�c4��ؿt�H�k�f�	ʹx]����ie�6<��cQUU��=L��<��_�=�܃��??�T2�b�#�mE�3���a�C��*9a庸�n,q�0�bHVqw��jmi�1�Z��j*�v�C��\�\��� Ad�6������^�������0�HyY1κ�D�	��y�bo�;�|���,ڲT��~������&$�ϊ5[�����e�H�����ϳ�`"[�.o��ܵ^[+�3��?D���� 2ژ���U7v:Oo��#��Yɘ/H̍��֨�uuu �v̌w(F�� ��%��τiSн����U� r��۷c�ܹ��{YYYRM��YK�Jc,�uC�Ktq�G��j���{[�������,6�{��o�� �;�$����a#��!}�TZ����$�d'1I$+I�7�d$��90\w�u�#.O`���'`Ȉ�´����\ۃ��|��ѩ��C+��,��*a�BaE�nǭ�+N��[Irm��h�S'׋r����ůlcu��}�79������v뮄�>'ӵ]�A\w�h|h�C��R��4B򤹶s���G��͵=2��i��9�v�db��=�~ma�N //[�ڮ�[6h�����c�?ǻ74yl5T�6�,ʷ����N>��c����j����D���rfΜ�Qz�	� ���VLV�� �uU�+����?a�9-Y���Ѓ{wlĈ��x;ݐ��̙4��kA������>�/?��;�}����ҴQx�@���q�_��G&.\c�+���߸����o��|ab��6�V�s��Ջ~��ϕ�݂�?���[����8@�w"C��݌杦�)�}��m�%��l���!{΋/x�,��Ea��CetD3�x��{��?�˗/���`��3Pݫ'� "W<|(:�����^���V�ϛo��;�?��O��'��*���ۖSRn�Pg�Ů��i�U ���5��\�Cj�PW/���5Ö�ݷ����9`"9�^@$涷�����Ib�un�=I�ﾐ�$��lIhu``��ܹD�S�~|������``q;|���l�c��ipm���Ԭc:]�MgN�?Y쫛�����"�u����Q�61�vW�.+�r"+��k�</�|���wm�9bhe_��=r#���P�Ӻ�b7�IB�n�����|�������;����y�Br�1e��k�t\�; �ṮBnmL�^�Nx�yB#"��qΝJ?�\�u���H�]�����D�^�+�@�6V?���>j>#Sl��{�޷__����o���Dn���ٰ�������I��=�>2�6�#��h��{;����N�#������j�U���Nu�����|EA��\�s�y�_�5K�ۑ��'��k��q"�t�T��.>SGL�������Ó�}�l�s���O��|���3~x?�a��e?�[��u�|���x�h޷�j�S�ƺu(..I�n(��,��Z��������uD/�-t��|��O<�ŋ��JJK0y�tTt�� ��uz��cN8���456��}��~�9'�pBZ����RUK��'��8���n�g�e�Y�Ю��hk�|�P~��6�؄��C�c�=$p'fXUa�IELR�
cb�@��������^I��lpcHgb�~�7bŊ r���v�L�m�n�f�Gpa{Gvm�I�âO5LU(���N=\�#B_^�_G5vu��r;�E���Y�&��z�4���c)��v��]L��:��*���<յܾ�h+m�f	��K�{�إ�#(q����׎ݧ����c^�8�-��\�+�k���^q"i��J�\o^�����˶��:�������
�})�qͶ6ܘ���cW����� �����m���.�ML�*++q����<��>�n�8[�l�n�dnc�a��ΐ�dT��+���$�,�v.i�'r�'�dG���<g���wafM���dA�����Gx���+�����r�����H?x߉���r,��l��;�v5��7�y�>؀l��g১N��a�!��&��a���xqŧ�M6��A�~%��&�lCKH?�s0a{��@�!�G|���YvJ���mRe�K�d�����`�� ��=�0t�p�AyE�ʮ8�s��җ�c�6��G]w�u<x0���:`�}�2_<m�5ƒ�^5C�5o��j�^5� �X��{�ctY>&c����D�VQ�����+A%&�
<W�JR�Ȕ�=]��K�,�D�SճG}���`܃����c�mg
��ԋEe!�!�e�Ipm�W���ڠb{��Ib_i��Wa��ۃ����x�����5�����*�1y�E,�qm��	sN�´d�����MSE�q���}��G��h����cwmO�G+$��3�M����ř�N�v#|�����;u���(ˇv�|um����v~ZiI)���x��g���/��m�z�-�~������c�T$���B�j_;B�J��b�k|�*,x��ŝOVَ]�mFyqo4��ʆ ��f��+-��?��� ����Y�[��/}D�QS��۷}>Pӫ]~��p_���Ys��M;����� ��
0q� ��3����t���;A$����\׀��OS,�;W;�j���=H�PW/t��<�l�K����k�.̛7MMM r�AC�`����]O�|A�Gq��ԣ�?�{�u�_�)��f��ݘ;w.n��6TTT$\��Uc,G[y�����B�Цs��ŝ��"�B�fشg���zD�Bw"!f,D��z�����ޮ^09I*��,&���Lґmn~mW�\i909�ACc��I�1�����"xF�sm��k{X�)k,U��{`�v�O,��ж�d�m�M֌j�4؞�1�z�v��sU�,�vA�m5zP�D�]�kcw&��sq\L�إ�Ҏݯ���L�6�vs��p0²�}�Ǫ{�����x#��<Q$��C�GX#m��<��ˀ��s�o|NL]��`�s���]��/����~0<�H�F_�憄X]ەx4�M��>��P٭;�||�u�L�.<� F��9s�dm2*�|��̑��~}�����b�����l'��]�-[���hii���6,Y�� ���W��K'��#s��'a���:�h87�/�v��VQ�\gdMO<x���SU�p_l=��Eؾ�c��t*�/N==+;�+�G�>��ӽS
wo t�X����X!�~�=��\3,p����X�xj���'c>�9�Fgu�?���Q���-{�� � ���q�������� �T��trl��/�8��_�k����c�]�����ۣ>����vq�j��QҼ	�%}��B�h�Bw"n����ʖ�8XTNJEN81����e��D�Tn�JLR���$U,m�:0̟?��� r�cFa��q�s���AT�\���M�� �����������K�mg>E������{	x�NW�����sm7x�4�^P���	���_�.��\N\ۅU7����J;e�s�`�Q�cMn�Y�Թ��q�?M�q���n��\wAc���wԘ<��A]�M�4�<�]��bqΝ�r�xLu���2���2�ڮóo�h�O�.ە�#�N��O�|�T�����އ��� r����a����R��e�#��*<�;wY�F���)9y�VV�#sa���n9��~#�T�bK92A����k�Z^���6���b���3p�/����	yo���CYIr���⾋�L��{��5��u�qoǸvb�oQaDp&2 ���8㊅ �D9�o+��ڒ�ޮ�٫n}�g�:��mfX��M�|�93	xꩧ@�6�x�|�4���AA�a���Ν��˯�1V��裏bԨQ��W����'��bi�1����n�����cuq���1����8c�-$p'�f�@���PR�{{d[Ĺ=SI�l��:���p�7bݺu r��>y"����!�p=���E�:���*:�y�`5�{���0Uq�:gx���k�(�Uc��ĺ��9�v}[�@V�Ƒ�$ͨ�@���c9�LM�d���q�N��0��Iqmw���&�ؕ��?v^!�Ǥ����ʉݧ���L�6��Ո����r_�]�ݾMi���p+���h['��E�@�GHν���~m��k�]�x�`��"q��(���nM ��k��:-���r;!��wذ��q����{；n��a���q�UW�O�����J*ś�J�X=X[�#�;��ǫ}�A9ae_˙N�J������{6��r�$� �s���-A���4�!}�,��7�}���"
��\p������|r�3{�p���SQZ�x�g���W�=��;N���I2&� �H�!�Ѵc�����¨�vYܮ�ٮ'1�E�{�t�a�fX~m�����{�����`ڱ3QU�AA��T�N���_�ĴD��4sÇǘ1c:DM0������ȝ�Y4�j��"w�nh=صc�vȋ�[�7�o���l��	܉�`C��7��h�qo�ەU|��+I�̾���4���F{��'-q������=��)@;�]��E-f�\ە4m�����3��*����rm��DZ���]����.�uն�A@����ۅv^�튃:\��?�2-ݮ�B�L��+�Y�)e����CP�!6�v7$�����ӵ�_(Ǐ�qmW:P���9�t}A;�r�34���t��!�h�+v������<�6	��kcҋ��i��~��sǝ������a��\p�1%�:��Bl}q�+ұ�;�	�D���n��udЋ�cuqo�ۂ1������AAѸ�/�BE�R�5k:*s&��OO���~	D��ѵ��W0��Z�_;n�����?إ�����ぃmh޷�Jsߩ� ��û�F���+Ƚ]��5�PLuC�A��{�,��a:��|uuu��k�?]{�2�+:c�qǠs�
A��{u̜3/�g)���@�&��l�ܹVݰ��2�z]�u�\3���a,���urg5Ķ6�����l="�X�V�cM�n��{�+!�;G�mž��R	纠�{&�
d7uhA]b�Oܞ�$U2O:2����Op뭷��]���t�г�����҈��֎\��刂u����]�)\۹?�4u9�ؕv��]�]ۍ��U�����d��]�7M�b��f�1Į�7�b��BL������N�4�X�n#n�,pm��,M�.Hm?���~���yا��� ��v;a���>1Y���<b�&��B��34�|�F,�������h�u�]x�j;uuPU���ɏ�{�ņ��A�&l��C=�f��ɨxWA������
7�we�sc'�l7ޑ���῜�]��PIRr	+[�>���� "�{�W�?�n�8q�HtT~s��X��3<���s����NEuebfL,�8��ɘ��9��Y������#/���ʶ]�Ի���i��H�#���~;JJJ���Q놼9�ƹ=S,�fh8�<��\7-�a*L���]w�����~J�X9L�U�s{Ii)� ��KeWs�l��ߥ�U�Dn�j�*K?w�EE��udc��my����� �ˮ�uDo'w��\��b4wf�5��P��F.��	܉���^���Q\\�8�j�vI����E�^I*х!�I*�rcH$���@�7ov��"7��f��.]���;���Nx����.���R[�PU��5�q���tI1�5�A��^^�/%v>6a�V�/�����9�05����>4m��x#�rx
���������z�,C#�v7��s��K}mr>�����)L3���v��?)&k����X5�۸�MwS ۽ɑ,�vML��¾i��ڮ�kjڨ󙦦/�k؇�ԗ��F��Epo���U!9��qo
Pۤµ=�	�$};nZ���������Ea�W�Ax�#,��#0`���AAخCtd��p���=���]k���>"w�I�vd�\��߂��]'n�]t"��]�8r@^��1DeA��O�N���%�y�c��v�� sm��Ÿ��3p�������Eq�g���[/�2���l�k ����4��;+)N�?��	d3l���۳�ݓ''�מ�|{���һ��#��?�q��ǀ�ܿq�C �x	���lG����ۣ�c��v�K?�3/n��{���H�Y9u��a<}i�H=�G�F}&r�^}�`���(*�QM� "(e��p����ŗ���- r�ŋ[�X'�|rR��T?�֒!����.�b�i���Bc,q�g��]qr�pqY�]ú"o �;3*�XC�B�0��ɩ/q����O�ŉ!LbI�lvc�4I��<{�=k�*�}�-X\R\����qڙ��sm���k�4]])��$�ڮk��̵ݔ��b�Ȋ����z�����nM�m���,�k;�Ů�7��r���K�C�3���ʾ�d�vg9�}��� b{�BM~P n_�Y�ޯ_ �\�=�o��R�����(�SW���a쬯���Y��^D�m�6̟?7�t�u��L6�,��69�-�dM��΍3�ލ��^��$��aC���wqw�T�=�yz܂����� ����NDM�J��~�FlmmDG�u�A�u��a�оxಳPեS\��n��Wp�e�D�Dl����?�N�6*��%�%w=�%�|�l���7���2}t�}}^߀��.���~���O,�Y��a`/rq��֝�8����n�sLm��{���$t�Ź��ꌱb�z�cu�a��~�!n���ˠ��1~�$�!� "6
�
q�13��+˰��u rV/5j����<����1���\�ЮF7�r놊1V�=�sHk�常kF~nڳ�kz��ۨ���11�O��m��U^"��M�Jp`��r\ $;I����1<���x�!r_�U�{�Ĵc��~`ǂ�ID��'SigJm�����'nk$�pm��r�vL����r})��ӽ\�S���_�I]OS�N�=bvm�׷�=�ߵn;G n�G~���^�k�kh"��E����+}i��z���k;�:�k��wy�����q��7����웩umc�m#)#�vq�Yv4��i��\Ѻ�	�vZ�yd(�bWVO�����6�4Sm��k{����ݿ4�Li�M�rک(++�KK_ �{���k�����|�C$�R���U�9�~����v9i����&�Z�)��]qq�$���}{�0��'�^C?� �c�|�g8�����o�sY|N�SGįΜ�k>"8��;u*���p_��⻞���|�J������gb��~	����8���sf䀽-����G��:B��{����_�g;�� ⥴(o�����#>s�>茱���b� ��l��������d ��Dnrȡc0zܡ � "~�o�I3�DIi)V}���c�Ν��k�?Ym8��]��e�1�Xӷk�|��K���������q;g�U�j����]?�j�Ņ=�J����D`���
������U�ƿ������r�C
&H#��@�QP��S���g�)>�PCB�"�  �#%��!���{��gvg洙��;{�?���3�9����s��N\��	K��T�4���O�>�k#U>�1lٲ^x�u 
��	㭡���pEO�"5bL�[����նjj����\u��<�N�wm7 ��U!E�����VS͚�#��7v�>vfitm��)�Gl{9Z[����J���]ە�ںK��R��:h��@�|��qb�?��n'�w_�{�;Iǵ�-��R�_I���vn�X�	⡖e���;�dM��o�d��|>Mݵ�;FW�x�|��q˷R%q{�\ۅE=�M�/n��}�|�XT��#�D�z�jx��X�paV���J�q�<�g�ȧ~#�����%r�l������g?G����.��Ka6m�ЊIh��� "��q'�q�_p�/NFiqr�����R<�n#�[�1���z�|��
e�wy�G�c~��A�����W��ǭ�8���r^�7�~y��QH<��&�ꆇ�/��Rٟ���Ӎ��ޅW�ߊ��݊�ތ�#�%�H�L��U����^���]3곟1Vq{��]g��Hg`����'[����/�Q����þ��AA����棢�o��D���k�����g��e�O0�r�C��}��X?`d~?'p��u�w��P5�bn�:q�`�I�ܻ:;q��"<@�X��Y>���!K$1��0�E1���qJn����O��7R�ȶН���Ӄ?��ؽ{7��c��)Xx��@C:7#�5M��dE�š�S�1De��!���O�k{̍ٔ���G˺yj��J�FخYO���Nщre��k�!����
�5�Ǘ��y��+��垟���Υ���޿��^�w�ܪ��q^���p���I���k��e���Η�
��:*/�8�m��d\��� [*K[?a��fjˆ��͖&�v+I*�y!��������ǉq�L5&����ǎ�ˁ��hH?ڑG��AU��]w�(,���q���[V#G�L��(Wb��920��}N���b�un�s?��he=���)���Hr�ˑA�Gһ�{q��^ܳ���&� ���>����}�8��x�:�.����{�X�T���A�(/-AMU��`>a���!����DZ�`��﮼w?��¿�>1k�e��r^�e���f����f�}/ZSX��W�����,��zz����]X��v�۰�Y������� �DUU����US,Nܮ�7���dq�W��W��o�YB����0_�}��Gq�]w�(<�>>�"L�1AA��}��FIi	ֽ�J\�>����kٲe���D+��X�'I����7����ɽ�3Ų�ͦ-V9$r���Dei�5�`�ƹ�n��f�Ht_�i��+nGLX�����ah�ґ.�믿�>�,��c�'f�����"��q��J��T]ۙ�Zjߢ ҍՉzUQ��d�fK�Sa��	_[�-��&�ij9�
�ڮI�|J�k;��)N�}=�=i��Rݳ�ڎ811Et�]�U1���-�w�B�Vl��|�����]�{�趑��̵�Y+}y\������8/���}�G�.��umO:.�^�{	�z�k�o����tt饗ZB�d��<�l�JG��|7]�n �sC��m�*�9��#ߣC��V��{d�س����Mt,�w>ޝע�t��bƄ� �H�;{�ƍ����4��x�7_??��>�y3��3?�r>�e�(+G ��*��xmJ��PUY�|/���Ŗ-Q�3AWw/���w����|��%�q��?�W��?܁u3[;@�}�]xw�nl�Q�rg'��a�]訇�oȞ�>�?��5��v{�g~����3��)S�fX^u`m!��F}.<��h�L�<	AAd�i��DYY���t?U`�������=�O����ڤ����?�,���K�3�r�<��#{�*�&w�g�~C��	ݻ���||���D�Cw"GN�GO]��+D������SQ���f�~��H�x,Be͚5��`����ܸq�`)@��V(c�Ce1���t�vU���k��)��G�:!�*浳L�k�$�t�5b{x�����
��ɔ����Z,K���x	��q�:j?�~w9-Y�v�����=CSW�u������J^����oۿ��{�u7�^���h�m��҇,w��B����u\rmw�SW��fj��c�8M^ʺG�Rum緛Z-7ͫ�Z!x�'�Tc���n�?z4L���$�>r��s��o��5���F�!
�x |0�=�ج6Fe��)����J���ЃZa��9�H�5�`�5Ԡ5G��92�D�asS�����������2���'��� ����[ǾG�S���'9�?�:^|g3��>�[�@���_�Ýxr�F�+�{���C:��/����+�P`���ۺfY����*A�M(+/�>��vI�^�هX��E��8�3�W(��E3,�Q���X6��G�L^Ab�ϬM�.��={@�;d�2�W� � 2�ĩSPRZ��|���
��;w��/����#S�X���1�"a��B�o�1��:�s�>�t�Œ)��Y�oh����L��Y���M��� 
�qVY4n��0J�^������UR㔟����@��F�t��ә�Wlkk+.��tuQ�D��\�g̊�L��ߜċLݵ��_�ӶjjSqmg�+u
�k;':W��b5�t[�-��&�i����Tѷ>��ԕ�Y�v؛Q��z�{\��X\��G��!�����z����b��}��H�rm��;���ә���f7���;�^M�\VԵ]��d̵=�(�J2<c��Ja��]z����k;԰��l���g̰D�ׯZM"��������2eJR�B��ؔ��h�t/c����]��.�C�UE�Zq��Ƚe�N�=o�� ���3�t����0{ʘ��g���9e9���Z�aOcN��-xs�N�#���w�_�Ԃ����ۛ��oEkG7� �e������v��]/rWG}���F{֚bA�Fd��͇~�t�h�-�܂�Da�\d=r9F����	� "[�N��G��=��WQH<��c���q�'��'���X��%�1�)�3<��Ϫ1��/F.r��t��Z�;3�ڊ����!�;��zѹ��奊���E��B�V��%r�5Xɓ����'�	�����A���꫱~�z�żE1�3}c�փ�����kD����WY:��r��sm��q4���J���R��V���]ۅ4�'#&&���|B�!��7ky	ĥ���4ݮ톽w{�]ُ�};]�u�y)�ȶk�������SW��fj��-=���f��F�������>X��]x#n��f�1�um��(w*��7�;�������6��Ι��ի���	�0hhh�^e��S��)G�l6\%3_����� ��&7T�C�V�C_�5�`��Ƞ9Ȇ�7h7Zͩj�ۨAA�	����߁G.>C�+^����`Ѭ���6�^6l݋��>�Հ|���מ{�Z0#-�=��&���ۭ}� "Y�Ֆ��a�5�,n/��s�X¨�na�ϰ8��]~6�3��"�}����������w}�pQ^Q��>y$�
� � �˨1������z�d>ZP\y�8������R؞l��L`c,��19c,n��1�_�!��yc����3f:��E.�	�	_�.FW�f�Qʧ�J7Ġ+t/�:0�6P�'���5���T#T����?��S���;A��}f�wb%"Xg�M�k;4b{��7k�������ea�.�Cܮ���-Ŧ�ڮ]ayC���)�Bq]۽�n8�
���.&�:�r)��[q���u{�uϪk���),gW]�������1Et�\ۥ��s��v���͗o�?��o��:!9����Z��Z���o�dEw��ȼk��y�u�J���#l��튰]:���(����RX�eh��q'M��g~��ttt�(�}�Y�q�8��Ss��Hl���3�}XkD|��� �2XS1/lw��9E��~��ū;�� ��w5��K���?;�j�L��?{0	��̿�݂�~w�ۑ��Q�[~qrR��:}�|�w���:��H�ie{��]�����>�"{�g�ɝ��B������C8����ܹ�:?yy��گ.�����絎H��
��$n'� �2l�p�z��#���D�CKK�e��r�JTT�����?�Krp����XŜ1V��+�_ا1��c�X��ϳ5�-T�(\H�N�r�.t���T��*a��"w�Aѱ��ӵݯ�J��S��r����'���*�V�v���,����Ҝ��Ⱥ���oTdaӆ�R~SCc��T�4�����zl[Kkdj��J�bB��8}��nR��O}�"��G��PY������V���ݝ]hkmX
Ww�j�~$C^>Jc]=�wMAЯ[V-�õ]�َlV��:������TѺ�v�W� 'ώX�}�޽H�7�����{��o��]󒅫]��8`���ڍ�ֽ�U��_�3L_��6\^M�MVC{EE�Z��e�x�H�y���k�N���J�'xd���ղ�q��C��=��9���ȿ���_����D���&�M�����m߲/<�^����,�!l���:��ް�"1�d~	��D8d�x��/[�1O����MUUn���}?���p��c͚5�?>fϞ�5a{>96��U≺(�o��*�F+~�Ag�A���;�Aލ�5^M-݋W1A6yy���s��	�&��g��VaOc��">w>�ι�>���!�5y.8�3?�&-�=F�v� �Ē��hil����>Ø�@��Ήܭ��?��9�~C�Y��/�Q}�:��e��o�������
X��]n�����\�h٬�}��Q=x0�R����a��~��}9�3s��l�9\��o���?��{ֶ���ތ���9��t�����6��|fϷ�kj��#���OjG��=_�\��{,��_~7�|3��o���	c�`��r���3����X�Q�Ց�������7dϗ�џ���b���xe�y*$p'<�:�m{7���<�Hk��5R	UE���/r�7X�7R�+v���F*�h�b�/��R����J[[n;�rU�-~����0�A֝��]���L��1M�R�:3q��ӼJE&]�wnݎa�FX�Ysm�����L�9]y�.�Zw� �v�BN>L���Ԍ1��i�Q�u��tm�Ҹ����6�������L��~�����nHu�%n���'�f�StVVHR��OV~_&0g7��ǎլS�������ob��k�w��vLS�Ѭ�]'�uҭ�[��Ü�x����K1ޮ�R}4y��G:lHdqE=��bt����}�_um��c�AĲ�󄜏��?wj���I�N�����7���s�㜼}�ĥ9�}�����x�"���A���� ?�Z�M}����>g	��$}�����ƆF�ܱ����, mRbq�.�5�_���Va~.��}t��g�v�����o�/�W_}5��N�l�,�3�D��tVJ��*^����M3����1�9��e7���,�8�m!w� "|\p������5ytB˕D�����_|D������͏��>�|�	�%�i��_�l����=�)�'"<G�����BW�?��3���F|v��ɣ��K��=ڳj��?+�Z����^z	w�}7*++֮$.S�|V6ۿX�D����ee�g�t�6�XS��������}�Y�֦f�ز��%�sU~G{������rA��}.�omi����93���[�}.޵)S474�쏶�\�ߤ��=9�?��|�η��o66���b���{,v��{,v�+c�T��ڵk-c�y��eM��Hl����}�����~C3j�U�:�������џYڔ�x��Y	�	OkE{��@%��{5R�SBcU�!}��O���*H^?�0��~�;-[�	�'i�7��2��}dq�)��R9^"Xi��|QZ�r+���uub���Ԋy�,�dK�*��v�zz�(�׏��\S�=b�)�X]OS����-�*G#X�t�B�(*��d@�|nx���3�P��M�ۻ�iĄ˦�&T�KS��q����)���M�:Hߝ���8��4���
W��ԗq�}YF.O�y'G�:I1^ǵ!�7����+��'l�XE ���+����F~�+u��XIܞ���;Ǝ�
�uy�j7��po��`��֝8����G���}C��(���z%o��c��[g���/���"��o��n�g�yfʍQ�uIHn~b�UjC���{.c������n���F+ޑ!�|�r�o����{)ƚ�Pl�@_�:d� "Yz����5���_}%�e�T��H���|���亍�w�%ng��_��/$n'"->��-(//wG{��Y4ǒ��,����Xq���Z��T��G��н��]t��7l[��FC�6�o���)�E]��O�m?��
���rnO]�h����	���~�����,���lD��!Æ�����wo߉��T���Ps��=�=سs�M������n�qֽC.��g/U�5�`T혜��K�۬�oǌ�'~�a���{,���=��ٔұ������^k���������J�h����u��^����ϱ���س��6�*��-c�g7��{!BwB˾�Jвw��HU�i�����8��C�'<�[>�	4�F�x�ݰ�μ�oߎK.�$go����-=�G�ߛ7N/rԔ�����cz�y��{���8�|U���������q�,���1q�R''v�����^r���bE�v��'N���5�)��[w�:��py�N���ݽ\�Mn�h�*І�{b��鬻#l�S+���� .�� v�:u�����A��&��þN+y�/����ߒw�1�'�;�,#u�v]4�=ͱk�I�~��Sm���q�D�^yi�K/����M(i�tm�.�[sm�>N��P���ر�cq�����/�\qr'�ɚ5k�`�|���llJ�|�gc�ΫїO��^�̱�k��>G�ss���!��*{�A�(�ڂe�F㉏��� �����51o���Dr�ߴ���;�yW#
L��_�]�t�DD�C�w������r�a�=�Ї���L�t��'p���+��>�Db�%�_�r%>���A��jv���ȝ � ����<��������BG[�D�D�x�w�j�*�s�9NZ>�zŦk~��X�6Ag�e����X��B�h�c{�r�X�1֘~f�5���
�Z��nBG3�@�5�7�`�ƅ�gx���Sh�JW#V��3%tg'o&n߳g��c��'NQ�^uo��To��5�v�d�_���2O['VS^RS'KY���g(�|>�P7*:��IYK��5+��n/�U�d %�v�X>&�Ӳ����CF�Ʀ-�6��r�tm�rU��vx-�y)@�}�-(�sI��7�2V�Cm�tǪF�ĵ�9Wh��������rXk���<U!�['�:qQ�!��Ju�
G�.��smwʉ�D���v��.Mү{<�v'�K=z�ɜ�W^"�0'	v}�uס��:m�M�#\6_==��bG��|f�~����8�n��F,ٽ���F����QZ4=�I� ��y�J�㮜/�m�i���n~��N��cC��������GGW
$n'"�9�u(��pD�}����E��%n��;��o(bpSz��tdZȞ��֣�>����� 
�ʪAX��$n'� �P5�ˏ>
O<�:�;@���n��2�:��CD���|Ay�|R��bi��B���1Vt�g�K�7dZV�+j�Պ�'��c��-�� �;�0��-��Q^^�
�97uhAۅ!��λ�;�ũ	�E�g���5�/���;{�1���ŋ0i�%=�`�9�͞k�Nڞ]�v��Jz"���>'v$��k�'nc+��k�!�%�|�Õ���\ۡIc�ޯ���eε]ZQ����+ʏe��kҴBr�r�K|��P��-(����ė�r�r��6�|����`<��N(��A^w���O�qm�뮋ќQ���~�E�I؍���]q��e�e��0�]���V[[�3�s6nX�D�ٰaV�^���NZ�\r�0�W?1Fj��~�~�jCUl�Aٍ��_�;Ϟ�#Cql�����)�xhcn�'b���D����<���`F�e�*�@�=^]|Ǔ�(2�iv-(H�ND��*3Pּ��!����Ms�
�~� �vm�!���Lp&�\��e��P7�޽�{;QT�Ï>U�� � "0�����'������.��"̞=Æ+���Ԍ�T݁�o��1z�2�*�:��L��џ9c����(-�EO� j ���P�V^���R��ʫ�J��^$4V��z9/$�ޮ�a#U�n[�nŕW^	�0�w�BL�!K튋�/T�ȝk{t�ZMS�������㺶�����i��XE�K׊�ݥ�*j]��b���zF�ޮ�J��8G-ĩ�kY|*q�:�{�J�a��Y\Z/��=�I�ߚP��먩;�]ݹ�$�[�K�\��U���+˽N�|��a'���.�\۵Ǌ�w����Wٯ5��]���ï�]v<����
)����IQH��ɣ�@�y���������4�������gƵ]9���89�HԵ]�&���ƍÂ���g�AgG'�ps뭷Zn�-�HcP���.���CN#,�]��*�y.d���	�9n�#�0�"iF�VT��GٸA!�/O��������F�$-�]8�ҿᡗ��@���Ad�����n��X�7��;,Ҍ���%�<ڳ�g�?���k`����^q�زe��SQY��>�Ճ� � �p��߇}$^x����?����;�<'-�����w�E�O<c,]ߡ�o���
��Xa�g�!?��-t���Ċ��H�B������hi��1k�
4̠�&M��P���4�ܔX#�.-�������@�&n���L!-�`�9Ƌ��,UѦc�C����f��V=]�!���\Oq�R��>A��'o��]+nW�6�sm���n3��{`�vy=bqZ!�	�0޳�r mw������|1�:De����]KC�����v׋�uu��@��v��܏!�4�i�u҈˕�b���դi��r���\ە��p�7u9��I�lJbwnI��ג�r�r9��S*G�Cp�vC>W��v���k|<AzPѺ��K����v^���4���n�Yumא	�vS7�f0N��Xu�U���^Xc�e�]�U�Va��#1�� ��l�O���{�Fvc���rC�W�#Ck�*
�P�>wu��*�� � B�3olJ(���xw�n|�wb��z$H�ND&Z��4}y.����"w��]5���;��GQZ��ӥ�k�������?����O��Cj@AD8\S�IS�ཷ�AwW�ps�wbɒ%X�tiF�s-l�W?Nu�!p���}�|��)c1��~[�����)�bYi%(i�F�X	�	�q؍{�A{� �E���=��X����v&8O2B�x��ٍ�����#�<"��p� nw�D�*�g�ε=&DU��
��yJ��zK�&���IF5�d>]��<�SsrfY(�m�vE��H��89M��f[���k��fH�خ���%j�����u��i�>�Vwa;p�r���A���>ism�21M�y�A96L��Rum׊����~KS�����c���C����+�,���.�7>�9�xM�8'&���n7ϼM5&��Jݳ��nh��0#}��n���S&��3���W^�����w���7ވ��:K� ��Ʀ�6f	gc'F���=ܠ鸷��EG���{�v�A;�Dh��6V�i��'������ � ��6���vf/-)�s�?���s`݋�������A�d��^t�����\�3�?�+l/*�o���H�_ȋ�S�ӑo}���֋�D�)�(���k�AA�ƺ��O=�(c��G�r�Jx���1V���ҙWN���?�zO��P�7����r�����E���Xv��m�%cu��������
��0���&TT$6Ġ3��5���D]2�H��F�d��*k��ݸ����E�?��= 3f��T���k���#�e�]�����Uŭ\���b{���x� W/KzF؊f�L2���+�Պ���W���o�m�vC�#�eҵ][^��k�sw�<�����vO��'������:�i���C�ε]�&����u򪳝&���Q���~����2�_���/Ɗ��>�c�P�Ѽ��)e�v�r�1푷t�s�RqmOPoh..��	�,4?�u��ƥ۵]7u�}��3Nǟ�����fn��&ˑa޼yy#<ϖ�]l�RNx�=�t�����z�8�����E�؝�t��1w���n�:bp�� � �P��/�:�1���ƿ�݂���ćD���i�)��٘g_�7���h<��C|������ ��3�����3,��P�Ct�	��7ƲӴ}�|?!�=��ܤ�/}���O�~��p˖- �MYY;�H:AAC��ң����z=��e�B�>��իq�9�8i���:?k�XV�~�g���;T�M����+�+�����mS,���Mh�F�X	�	�q�t��C�Z�R�Hh�*�3uapO��T�\��ǫS���a;w�n�k���X�]�P�傊���v^�TH.�n+}ե�� ѻf�.�N��m��(N�N��m�_G~�N�˭��zʢ]N�,e���x�m�nw?a����k�����B������lx1-{��B�|�߶u��A�EN]���Hu���3���$]ۅ�\�XT�|�
��.}�v>��])KSv"������Y�sm��A�;/4yl��b���!��m���k��@0��',mǩ�]��m�;0�/i��3��"��3f�?��_�a��A��q�%�XV����,���wi�V�Fl�5ܠ����1D�)�#ϓ�1W��"}C/r���d4oCu��vӐ�AD������j�߹�^|��>+e�ۍ��v����`B�E�&8����6⫿�]��b-A����}�CB���1���@ߡ�)����?/�}�٘��3���{�n�$��8���AQ�9K�<O=���+��v�mX�l:� ��0��X��D�o��w�>�s/B��X�����w�s�������� �;aq���65&��n-�5R�\	ۡ;щT�6Rś�o�P��?��x��@��I�L��E��A��1^d\�a�;5ǜ-����<E�nih���=Ĳ|^��;�IU���vN�n��B��M��qZ�v)����&�|�����ٹu�_e_T�3zlh�$-���\']�)I�����>�����)c���;���%��b����/�xݺ�ǉz�Y���9E��[�����Qʇv�@��bz��O��UwUH�َ��-��ڮM�^�
˵]'��s��8�?���o�DxY�~=֮]�o~��ƞ\7,%���26q��F-��
���*Sh����|�L�Rc��p�ݥƪ�'��!	� ����G���^������-8���h���_�Z������^�@��7��ݎN���V����%c��"Y�n����N7�����4�J&�\�oii���^j�N���/Y�#F�AA�ɈQ#���C��O[}D8a��]t���zTW����?�=c,Q�K֐��X�)V��H/p�0�b�@���
�㍽����:18�TE\#U�\���xRmJf�\ͯ�����p3�f0.Y�|�aTo�׵�O��!���&�Kл��BaE�n�[�4��J��L�T��@�rrf)}�^ +ocu��	�!��+ǀ��Ų��-�v�U2�P����h+1N�޵]\�%��y	U���F �"J=eq���,\2�ڮ�G�� t�'���S'S�K��������u��Bs������=���8q�N���M���_�v�N	���'4%�OqmWҌl������ �������DxY�f�.]�ٳgn�����D���rc��A�������"O��wc�VT��G[��p� � ���RQV��"�Z;�?��⢤���׏A]s{�;����f|��w��� ���|���h���T�c��j��=kj'p��<�����L���W^y%6n�"��}x��%3�AA6��cᡋ��g���&��lذ���;�����Z��	c,y~\c,��t�c1�����y���w�
Y���7�r��&������X<�-���8.n#U��*��ʷqJn���8��H��<�=��������A���c�`��I�}�(���9Ƌ��n�j='6S��U��q�A��:�3'���5\OjEܞ�k;�tS#Xw�)�]%q}]YA��pc��Nŵ�]uw���^H˵k�U��.ޏ�u�^s��G+l���따k;�oͱar_��BSGSS~����o���I�g�U�kFr���cM�;�E��=�d�e��<�h�9�+ŉ)���#o��ν���]�+yk��� "xum���C�8.ۮ�"�[qԑ�����>"�tvv��/�5�\���2+-^�O&�g�1K�?O��nP�ˍUѡ�}�u.��'��� �PAw�;Mm]��G'��,��v;򧳎���Mx��(D�z��[���� �L���{>v���
}�v?bQ���еܔ���L��|9��^��w�"܌?�LAA�IS�������2��r��7cٲe�;wn���0c���ÐF~��2�*v�
���c,��=f�U,c�l#c����ס3Q�v������C�Bwم���J<A�T�\;+d"� �T�=���^�e��X�|��%���7<�]�%ѩ��*��h����D\�U��	5S/����S�����j���[2��.�O�n��(˺	��,�k��jƅ��Hٵ]~K�g�:vE�}���Y��R�ĵ]WwC��Oݝd9��\+nW�+��>1�F2=b���v��5�����oH�k;���q��
�w���_�#l���C��h�Τk�����\U��W�ȼk�P3vĩ�]�R�Zk��D�Еk���m"�殯��L�m'���c>�)tv��ǟN֭[���'�|r���1K��3��*HW���+w^�n���5V�V9HA����bTU����׷�^z'�����I<�<����J"�~���ذu/
�����6����A�������k���X�;���n��eO�����퉎��3���u_����с�+WZ��Dx����}K�{A� � 
�i��DWg�~��G�+dzzz,c�իW����JK�+���cI��ee#Ic����ݚ�ѕ�����
�pO(AkSC ��"n�x]#�ށ�cx��❴��%�L��Lv��Hu�WP#U��<K�8�q��#������]���Sqm���=���!=�j9�n�b��vmc^#-���++h9�|��2G���z���(���R�'�ڮ�]#����ѻ*u��S�{h~7M=u�U��Ǹ��NH�@�c&]����Y��Ԥ%�ڮ�C�./h�Kε=&$�~�x�������R��si��)�A�������}�hlh��^>�����.]��'�B؞�2�Jb�i���<���L�o�*�L��+b�T��U:��&| � "d��c`��1����ڇ^)8q�́��%��;0����~�����R���C�+q[d�������ЊB�����_�B�v� 2JM����͊s{P������-&����/t�3�E���>B��7�x#�}�]�e���a��fa�R�A�@d���������p�~�z�y�8��R����|.�u��E��+��G~�`1a{��	ڣ�����hَ�����8�	�8��Б�{{�F�D\Dn�|�T2�dc�ڵk��*ĔW�c�'�@EeE�Xӄ�����ѩ��*�o[۪���T����TU����.
x�:z�]��b�?�sm�qL�+kF'\Y�OS�1���.�)u����k�f����[���-Kֵ=u��&�����;�V���1�Ƹ�t�!�/K��Z~|�v8y��v�Ÿ+���>�y�C��mq��[D�������ܥ����#l��+�j�s�\w��HU�_�Fx���]Y�D����.ot�?q�u,l��~q�l��]�ߓŴ�qn�j\T�{�i����|��Fᣱ��V���矯m�	[�S2��k�29�{"�U��]h�*r����|����^5o��*� �����|�q�A3����O�1���=�k���es��`���9�z���S1e찄��8z(n������n�(���{p������Ad�#&�讋���7�>���Xv����v��]���dK��}���n��&�e��i�oށ � b`3�������?N�1�a��)S��0]&W��ɩP,
7�3�|�?�}���Ϧ��9���XEE�M�lc�#&�1V�!�� f��R�46�<%�v��a�I�*?7��$t�����*İc���Q]]�g4�k�c"KU{(ƈ�T)6�k��CJ�햴j�ᬧ�W-'�k�R!hE��t[�.�BJO̵]���5qirm�Y����|����-FYAF�,ʽ>`h���d�j�f�������|�#���\ۍ� �?��j�Ǹ��NH�;���:i��/n�wm����(P�v'��Ƹu��]�#n����Sz��=��Jޚ8;6��rm7�8S�(����f�!V�k�5�V^^�o|�t���Oؽk7�����bŊ�TOk���^BwY�n7^ɍU	��G����:qsq'4� �PP\d��� ����������t����s��ĄM�=h|�������W_���D9`Z-V��E�����/�/�m�ی�Ͽ�� ��$̽��qK��Ŏ1V�3��ϾCO���gܽ]G����W]u�5�3Nj'����� � ��`��ֽ��;A����6\~��袋�}m�"l�d�d<c,Y���=S�c%���&2�
7$p�L*�k���s`���{;�He(U^0�*��r��#��T��r�J����l�?��e>r�o�i��&�dq�.9�Ft*���*Tw�̸���Yqm�V�R_)�]N�,����n7���c8�ʂ|�ZN��J����v�����0�:����'C���o�������'Pwq'��;�꤫���v�D��G�n]ۥ4�~X2�ڮ��-����������-L���@��v���$���/����	๪�/�CxT��	�v�\��k��K��:�v�hs��z�Ĕ��Y)	����TUU���9�^t1��@�v,���bȐ!����g�1˿��m��j����CT����{o/�^B�UD�2a�JK�-���&c��J�o��w<��{��Yh|������;��9h��Ə����]��r�g���,�eZ:�0��Њ/��F�����h�Ą�?r�t�����\q��o�/�}� rCԽ���	��q�X��X�s�"l<���M��ԇx���駟N�����-��}� � ��-z�G���"|<��x��q�1�d]�o~>c9#?'`���yW��)VPw���rq'c��B�ʂ�%hi�Gyy�{p�xQܞ�{���
j���X�T��Y&Wn��w�y��d�!�0v|�oLT�/����+�NI �um�3Ј[�<�Y	V//��Rw>�C�.�Vź��v!��v�صH�k��D]��
*�&��.�"Ĺ�u7��w��K���ڮ�ŭ;��h���Hڷqm�z	@�N��vy��5�cZSǴ���u
(���F���oajb��,�1���+uJµ]WwAH�QwUH��1�KjLJ��X/q{�8�е�[�ƙ)�A���k�s/96�:�L\v����	"\l޼k֬�w��]�F�|l�J�2�J���X���[�^�U�96��P�:#���I���XE�5O���>��
;��d6~z�
L�.�;b�4���[��f���?s���S��o�l���C��-3zX5���C^��m��76�v������ϗ,�z���'{A��;�B��Q׌�2&�����AD����{���X)����Q� v7%�ޞ���t�w�^�^�D8�\m��\RJ�� � DJ�J��#�����D�`��W\q-Zd��曉U�c%��n�)r�Xd�^�	j�2��%��0�:���*�{�,b��C/J��*_�t$�gCCV�Z"��7� L����|�"'#K<���p���Br>Nl�5�vM�Z�n�2�xq�R'U�kIU�FH�k�4/��d��٭WC%.��	q�&.ݮ�8�����O��ƚ��i��I�k����u���쥮ʊA�T�A�(��|��wf��?R�^vC�3"����n���F�����r�ܴ���a]/���"��RkYLyd~wOtxy�sd>�E�|K�����:��Յ����Չ�Ύ��N+N�}ma����7Y�vΑ\�7����k����|9v�&F�p\�5��@���k�V��#X�]�]ۣ��_�L��k~�X}D!�u:�
у
�����Ԏ�ӿ�-\u���y���z+V�X�9s�d�a)O�,��XŻ1��X%���t/�;���k�*nۆ��q���n#�0��+��y�w�����G!QY�c���N<�&���Ԏ�{~{��˛�~�.�AO��('9#�T��e��a�ܓGUEb�팦���bdGW��f~�Y��&���'-���͸��u 2Ϥ1CqǯN%w�	�O�\������"��=�v�з�Px�4�I%�����o�5�\�]��8����C�\���
1�`״ʊ����#�GG�g�[��/Bww7����Y�_�kA�GEe%�F���#��۶m�7܀s�9�IK�p*���d�e��ߓqq�ͱlc��'�$c��A�ȬQ%h��k5R�B ~�AU����ۓso�?a����=�XW_}5v��	"|L�1���㷟�"�Ћ���/:�c��G�v[L�&�bY7O��Z���]+��딄k�����Ă�����tû��]��J�ڵ=v\xם�QL%��++/ð�!�\��j+�4#7��0��g����hmnA��]hkk�&&�ʦM��أ�"U�5���
���<�G��¬�k���(vg"��Hݙ��n��o�p�&I�k;�����	ۥ�D\��"yE%m��q>�����B�8uW ��1N�Fx���n��d˵=V��T�q=���j���3�A���k�{��`�ҦϘ��N=���D�`��]v����:#�vdϖ^D�:ȍU@��*/w������ϭ����n;2tuva��"<�)��� �@iI1�;�8�ww��u���`�	��;�Ì	#����U?:KϾ
Da�?�L�ńQC|�>�p���i��ooC}s;�ʲ�Zn����:t����/��-8��	-�ne�x�g�������g�ԅl�g��5?>��� ����$�ִM�;}��bw/c,�_���h>C���X�\���ه�5��^����7���8�kj@D�(�\�BU� TE�V�~���43f?w�6����L�^QQ��.�0��?��\��B���	��2����c��e$���2tv1s��h��i����s�$3
imo��cvt��=���j���#�ӏ<F�X!���o����Ν�R�\������3��xc,��P��{�������cՂL��	� �մ���k��pq����f�wg�wo��d��6P%�Ho~>�5x���q�=��#ǌƼ�j��+�hĘ�5�1ѐ��\�*"��H�õ]�rBaW��;* ��cˈu��s�Z��<ëRV���p���u��f-�O�n���+��,ȧ��,8+$9����3���nW3���\���q�=���bjנ�(Byi9fΜi��Ʀ��>t��[C�n��c455��"�_KK�5���#F�@EI)fN��\���u�5p�76���YݟyA��ES��.��7{��=�@<Z��#�+Y���N�tm�
�u��g���+���=�v�pm��P�Ο������K�̵�>#��;�#M#n75q��=����>"\���+���{q�����)��v��J����� .�ȝwq�����]l�������B�1
}q��"l����Ɵ~_�Ƚ��?<�0�}��(�ܳ�9y�s��үn½��_qŰ�g����N��-ؼ�ac�Ա���'&��ۼ��n� ���ꆇ���??�Ȅ�-�l�?��%|�gk���p����G�ˑ}>�h� q��3��:��O2�]߃rf���z��}�Ŏ{{q���a�3��M*�b|��2�����^��'�S�`��������KDn`��Æ[��!CPlĞ�b�����1�x;Z�6`g�KH��9�����[H'���̱l���cƣzpuԔ��D`�^L�2v��5ԣ�'���D!2j�h,\�/=��p�^,Z�r%V�Ze����vI�a�&���X�wC2�R��l���X1s,f��tr1�(mlD�0&)Fk��ȉ�<���o��M�Нo������*z��n�bd�q)[�$2�=D0�D܁���=$�|���˘&<.�<�8Tc�1Q�~?��n������n�K������H��׈�=��Z!��E�(W��ӵ]���%.�k�X�O�\�_\��������u���/�_S��p�;�k;k|*��Q#��'�fo_�f�DC}=6���%`���F$���������%�c磡C�bܸq�6aJJ��@q$�Mm-���CgW�}�R���>+o�[�B�ߵ�s���]Zέ��c���iA��k���������v�sH���wu���r�6�+���83`�U�4��L�v7�[.�=���Ϣ�����e�5T-[��F�J�q�{~�]�SYƻn��"`c����m����,w�"K�9h5RIn����V,�P��P�QxT���柟���x7|�]����N���>3'�Jx���R�����8�o����Z]�;m���������>؎�0�v8n��)<�<�对�y"���Y��w������p���2��S����=M�w�
����8���ȝ�<���?�A��b�De�N���(#>{	�3���L�&�YT&_D�:�чx�-����>��;�&N A��]�ƌ�qc�b�0vl-F�n5�3{�޽عy+�m|+�:Vg�_��齵Cf����&��������"�Vl߹���"�L�g
Z"��;o���"�[��2�=���.\�7?��X:w^��cY.��X�n�1����=��E�ZD( �� �Q]託��i���\a{L�^\H�.7P�����T�¼��.r����p�޼[z�(/;(�x�Rum����
R�X�|;w�Z�-4VoNLmy~by.ݳ��v�Ny��.J�=ʉ�P�\�c[͐����T�e��C�>|E��+���*�[���j��N�H�غe�Y�&����������a���GCC�5�_��Ig���c�b�ĉ�0����7[�z�������h�
��O�.�=b�|c%�^B	����Y'.-��h���IU��q�ܒ��ӵ�TӴ���q�X/1�����vII^�C�-+%�z��vq�����I۝5 ���S�w�l��1��'��t�M8�s�������BjJ.�B�{���<��G��C:��In��%g��i(�)-)��sO�D��?�� ������g%$H�).Jn9"�a�'��V������~�V��~�5�{�����ב�Ԏ�;��Ը�^l�݈���NMk��2v7��s��F�
ۇ����4�v"Ӭ۰�=}I����Y��g쥦�,Q�1q�P����X�oj"���}���
� �ǲI��ljGyy�22���4�ﰘspWM�\q����k�����(�0�J��t�u�V�́S��}��A�ePe��P>nl-J"�(�oX��1�{o��?�[7o���L���^/MUF�]mm-�?E�%(++Eqi	v�ك�w���Ad����֖Vl�h�p�z�j~��3fL����3�e1ƲRݨ���(rf�Ż�k��Z��x�h<��D8 �� bTU��[R�  ���������;1�'!���
��*�|i�Je� y2��뮻���!��ߋ�/Cu�`!�4�{3���bL1������0X��U)+Kg˵�� �R����S{
۵Bx��g�@��m���-n�r�ܟѣ/a��g4ή�>�~wM1J��8Cg�7CSW�{P������1���Zמ��>455Zo*3q6�^؍>s|g�p�ԩ�>a2��ˬ����	{,������$�x��h�&/C���'^�r���浜WݵB�81N�FP���.	�}�؅��]�c��C�]�_#��=Z��\ot�ڄ�q�F�n��E�H {Y��o���~�A����G}4�̙S���t7V�.���i��<���,������Bf?����Á�#��j�"
&r���/��7?f��3̵������G��Os�;���چm8�w��_�W�̄�l�5y�_�/������A��}Ҙ�_���-��sw�y��wq�ooÍ?�rܗ#x�k"˰���<�����s�}X���~��y������Ww>ܞ?�&����c1��"�~��Q<��C�=F��Fgq��_�3�E�Zc��"!�˹�S��Y�yI:�~�N���l�&Sv:���k�J�p1r�h�_L#�D�6d(��2U���vv�hjl¶�[��Hw� �Pl�ƍ�dî�#G�Ĥ����}c�Z�[��Mhj�kAd������V���"<���c�ڵ8��s���8�g���3�3�]��>C&rgϙ�VaL�ޗ�1����Hmj@�� ������E��p�1��#���m��D�]i�R���L&����/�믿�r$���E1z��{V]�!��|k��Țk��'���=��)nW�ԉ]ˉΕ��X{%��1��!|��Tˉ�P\�v��ԕkz���q��C��������׵(--��1��)����ض�?��ըB䆶�6���[��`�x���iӬ�{J����Չ�;w����m��!n���1�.)�v���y�vM��(i9G�-	��k���ō���~��m��s���|S����jjj𭳾�?]xzzz@����^\q����+���vTHG#S���l������9��Sq���}V�V��s,���s�Qь�1𜙈�s4��iGb��1��GWw~��Q3��r�������ܖy�e"w<��&|�¿���91����-�A���3.�+6�ʯ�m�v&�N���ڄ��z�?ϼ�N��Z���S0�&�5���&��g\t���I���(-)��g���}Ƅ�x���y��ͱ�?{	��_;_��´�w�O��{�A�c��R�67����w�g/c,�+�|'��U�v�ȝ�?�bpS���&����^x>� �pQ=��,_f��A��oj�hL�0e�l��$����FKK����ߏݻw[����1y�d̛5Ǻ\���Y.�o�lj�����F{[�p��m�1�QG�y����a{`c,+I���Wߡ�gȄ{��X-��8p������� 	��ˋ���qtH�X�0a{��Jpp/vE���:��l����y!�e����۸뮻@��}���}fNw���x�ε]�_�!�+������8Y���S{
۵Bx�7���e�v7NW'���{�֥rM9ΐϴ��a�9��Hi�zj7CSW�# �kl���L7�G�B_o:�;��G���^!W�<�5f�رÚl�{��30a�8k��֎��pi�n|�@<��<m>�qK3�)O:��'N�nJi^������	�|�4��:�v�|I�Htn�I��M���N��EȞ	�v�t��c�&�פy��}�õ]}1�Ą��_����Dxx饗��C�3��LV��3�rRuq���ƪ�.{��#{��s\����ݘ1b:6��� :�z�����d��i�����X��ﭼ�7�B>p؁���~�F��媿=��y�����?��5JA<�;���[��<��L�����TL��s;��+�zDƺ�q�O����=�G?�w�ll�݈���/d�[�������}�r\}������uaoS�;����k�=s��MK~l�o{Ad��Euh�̰����,��H0ƒ'�(�C��-ˉ�4�ϣ�ϩ���2�gfzp��W�H0d���a�G���A�FyY9Ə�q��X�X����K���Kd���
�z�}�f��"�ע�Y#�E�%v����M��L�"%**+#����?AOw7�p�4�~����Bii�����v�vq���=�7S7ƚY�D�X!����'����q��*n�AQ@`;0�N
����J��bv��Jm��O�2����]Ԙ�#=���1�j1g�\�sb��O�l'��.d����ѵ=eq�R�]ۥ��]�iyC�fo61�D�\�c���乢h�Ȣk��um�����q�P=�
��ￏu/�L����w�^k�1bWѵ�4e2�뱧�N:5qCݿqm7�Ӈ�>8���Svm�-'��n9G�-	����n��g'm{�ܥMJ N���S�.��
��X_a;(nc�v�������?��c�{����,]�C�Q��KcU���2^�U�}��X�!r��w��y�b�^ϲΰ���}��6l��Nf"�����m�<�f�OK~��3�\�M��ȫ�XpOcn�}fM����G43�����Ǳ��W@>���>�q�]��/���D��E��y ��6#W0�/;�G�N)&�߲;�\��[��3�]�;��+�Ĥс�;�K�����	���ܻz���ǡ�8ywW����?=r�g��W�ӛ$+����,�+�Ғ��v� "��7�Mu�{��G�na�X^�v�y/]��:�Я�h���_�5�p���Ň/�F=%"q�14q�L�0��?lokǦ�>�3o�"�a�[�l�&���;̜���
�E�m�lh�T�M��!X��<��S��/���5"ӱ��p]���5Ʋ�⻸g�K�3l�ߍ�#��:z�8�!�� �,�+�l�K7R9U����w`��ۡi��5P�d۽=[Bwy�?��<�<9�����j�lIT��%��ϵ]C���r�JYYZ�Rng�>ub�1�%5�q��qm�S{
�5�
�vSZg'.K����)���Ҝ����Ԥi�G��Ѳ���j�?`��i۰����
���A.uuuسg�Ր���oc���<~J�ˬ�hˎ����Cs>���J�	%��D������g3n �<�+�N���qm�+��<h�z�ӥ��{�&TV]o݅@sΆk{B"�hj�8�4q��ݵ/
8�4qb�џ��oێ�^&_Xغu+n��f�y晁�����;'j�n��4X��Ѿ~ΑA�Pe5RI�ڍV-u;0a�4lm��*"�hh��q?�}��8�Ғgq��ӎY�/-? 7?�*n{t�۲���(���[��_��B,�*|NA	��o�'�>��I�Ł�C/�����]���D��>}����E\�����ډl�d����/[��T`�m��ч���-8��kq�/O����/���-{���3/����7��э�?:�e�w�����N�4���!���p���3����/�80my��Χ�[A�gVu3�{K���8}�n�a���^\�������ޮ#��0#�5k֐x)d�p>Fצgd�(0S���Lǐ��V���m���O�� ���A�{ ��a��sQSS���^��4����t���c������A���l�2:4+}��#l����z"]�aƍ��>C��ԥ����$p ,�T���nk(���TE������X��ޮ{�P����L�	���l�իW�%�%8��PZV�-��E�"���p]��r���)nWꔠk�RM�� ���[e)"xC��w��\��;+~�;�[w�K��}���DEy��3�e������o��Gz��(l��w�yǚ#G�Ĭٳ1�f0����������)�!��rm��Q�Ը|sm��\SVPq�sz��54�X?ز �I	�)�u�|�(n����15�X�%lW��ow3�v�D���W�c�v�ܾD8`�O}�S�g�}�.8�T#S���j�\ܹgC��J��VVC�Ƒ!޳�3���ЋEû����B�����߹�oX��6��kG�ƣ���{�51:#尉��Ճ��^'�	-m<sn�XSU���g�r���(�����Ҵ�[���߾�xr�F&6>��wc5sr�v̈́�?8q���!xw��k��G�𷮹�z��-��7�w�%2�E�wv����>��Ӄ"ϸL�<xP����1�>�R��a��J��ĄQCQ;���ʻ�w�'�>"y�y�?�7��D,�;-�2��U?<��l�m؎L�^���ooÚ�|9e7�Ic����)kjl���V4D�6F�����ȹ����{{���Սp����~��+�JQ��F��aՕ�>>"���Ze��n}�����>S����n��+<D����N_�6V�+�g��l_%�̪U���2��g�>S1���� 
v=_;�m�X��Ptuv������������Gcc#���K��Cuu5�O��A3�QVV�{va���8� ����~hjh��M�A���;w��o����='-_D���+�c�ֺ�W3ۛ{A�/ԫ[�������� �V�T\CbPq` <��*�l9&�;�D�a������0��=G��e�v��>�?.��>��Ғ��ݬ3��~Y��0R�z�<9�����}/!I=���ڮ[1�����-�.���cWX+l�f����Ų]]]�uo�"L�.)����::�#S��eu56Li�����푸��N456i�}ut���<�{��(U���*tF���Ǟ@kk�5��y�Ɖ\��;;ߖ���|&�@+����C���lڴ������g���Q��"`��=���҈�5�� ^ �9��ݳW���uo*)a�s��C\���aod}�[N��rP�4U�h؝v��:�w��W��kU��8I��mؽs�&;CyK�v�ruҍݡƱ���n�����P��f��u�׋���m�mعc��=M��Rj�m|����>r~�weu��=�ݩ���|�����.�����D�r_���*���K�.:2���~ˑ�s���o�'����n�VLEc'u���u��7^�`�%�7�&��W��X#"�l��{[q��wa{�zd|�]|뢻��G'�3�0��i���;{,A?{	�H�-O����_�q���;G���/���^�����o|��~��6�^�HC�+�)_�9"�,ށ���`~��;����8�vow>C��gR��t���O:�y�7p���C���C� =�2s�t�5��}���&lۼO<�8���+\�n����#L�<�Z���blߵ������%���Ԍ��F����oǧ?�i̜93�D��,vc,��3�Z<�m��Ld�8�+E{�����q���oq�F � @����l"�b�E�U�9�����ɓ<�嵝�Mlǉ�7��:�dK��%Q�����;)�"	6�$z�������������������������~�6dddH�SsaP��7��i�T���`soקUTT��w�U�m�Ѧ��7��|u�+`@�O�<	#G�BwWW��R��
ٰ���� `�b��=��x���4�V?�/>A��S}J��BX�ݝ�����ZZ)�[,Z�����L�m�p{�����޿9\�
=�g�G<����\�Mk���;��==��W�<��qIȘ�='���cİ������hn;وȮ��M|`e�]�]e�]>xv{��J�ng�,6b���Ŧ��kܩ��۞�F�b��{�{�Ɖ��یx)�bf���]�����{ݷ�C�
�Ƶ]H2VI���++�p�����F(_�@",�fnhi�����D�R����V߀"�HQ���c�
kwI�K�{�����X=.�\�v�l�`Sȭ�|��ʵ�|;�/e���G8t�V�^=�U<��U��*++�i��?���'�^�ąAKcϧ�E��2�ca�������?�<Z:C�}~�1��ŝ��<Al>|	��d�;B�{��?߄+����G��M���#K-mS������K��;�Ǜ�ת��_��7��5L.���������@�=��B뽛HMM�O!���)��1�"�/�:�C�7��#��D�Ň��ۣ���z&�c�>3��D���23��6�U>�K���@���i��1{&j+>�Kks3��o�X�3j�KDj�3�8Ю�;�:���@բ%��^���\�f�ύS�����!���TU��$�lև`�1v�u��Zo��7�`�6��	��:xP�������c�NKG���5wj�>O�`�5��,�N���v`�������v��Y���E��#v�c�FD}��u�~��������(d_�2Ɗ�1�1ݍκ
d�OBsW��">��}�S�ڈ. ��_��" M�.ua���}P�V�op�Hs�Н=��Q���v
.�,_�;0�d$��8K��|8k��� �=}��|����+n��r��,�0�Jd/�c���ra�I}t��i,U��)TT���1y���P6�ӡ����!��'�onh���_��s�ȏG8vE�&�I=��'o��n�l~aa M�/�&�_��%/nnΝ���5�Ǎ+�+%CV�~_����!5Սi�� {D�::p��yܺqӿ.�G������FӨQ�t�y�v��eÆ������?[�6�/¨�\�{�U��bbm� ����{ܭ���S����X"R7
�=a�h����{ow�:cŔ�ӂ����kZ&��pߵ�$Bt�;��\�'O��aÇ��	۵�Iru�i>��>}��qص]Q�G�Y>�[__�LfΞ�_����d��g6�>`~>k��e{"9�!��Z}g��^W������ݮw,vͳc��+V8���M)^RR���Na{<�U���U�"Xe%`�ڧ}.�C_�8 � |g�_}Ъ�
���	�`����~��h)�����b^��]����]A��4�E�/l=����[�c�_�|3�k���|��6����������)�q����������?�����ę��z�𱲰=u)��=Ԭ�����+�s�L���|��-b�S�9�ivo�s�N9r$&"�HaO��*�����Y�U��+V�%�J�7&/��1Ҙ���v�S�\��o�3:��m+����P�����f�x�{v-M_����p��p��ܺuK]�b�c�L�Z����Փ�]���<vv�c���gBܼ�<KF5M~M~~>�-Y���L�ܩ���e�pP���<+���卵���}�����x��H������fw�������~�����ٳ�ڵkcއ����c�}��5�ZSl�¡��}3%׍��{HOO�,P�.\�ʢs{�E�����x�����?u�v��"9����V��KD�$x�߾�,�N.�@'��ۥ��F��¥�yė	���/'���g"��'Bw@�:ydR?S!�XM����ן�r����̵�@\9j},�ݟO1�i�v~/�Ǹ�QܮK����׎�<�|���aʄI��6�Ο;�{�� �E[[~�sj�����%KT�{cK��b!� ]K�?�e�t���	��l_��<|5��>!]��b�(���ZYKE��mR������ }� ��R�:�|���˷�5��'{5���p���9y��p�6mڄ'�|�A�x�xB��߷D�.wrOᖠ��������
���V,��j���nBvÞ�m<�se����z
����I4�?��?��wPy�	!�������o�u�D"w&����D���w���������r�����o<���n$���|�����~�|���1�8r����p��A�G�n�2um9�f�e0ƒ��M�!͇�[|$ʽ=V��v�&��/�& bu���[��U>+W["aQ�2�u��zI��#$���~��.�ʷ����gW�Lp��x��<�S'MƤ�	�xO׮����#�uf.�j�69��so�Lv;�=��*_+;��X�����'�ϓ&M§�[�=�
�ߺ�[��b�y����z{]��[;�L�[�qE�1g�|��gh�;���cg�v�mV>��i�ʕ�0��6�pqW{%}�2c,S�{�����p)c��	/$	�1Kr;�Q�2��F��U����(^\�}�,X��`0�������_���)av]�X���=^�.��+d�v�ې-��D�.#�w��K%(l��[�����w�K2�ORw%�h�C����=$u�	���g��X<N�d����  27v�P�_�Ż�K�򐺶����4����V�o.�d��۝����dg�NMvl�F�."�0���W?��՜y��FyU��t�����=�h�!F�Ǘ'�hݲ >xK0䉗k�T�-y��򅯿���Y ��(�"��v�9QM����#����$Ͳ���|B|��}��O�j�-/E�W��uTWV�����a��^x=��:��l}"�L��Od�I�U�����?�`pq��|n���.�����_�-y$"8z��������Q|~�\V��������v����Dh��?���Ϟ�>���	���o���Q�P�W�����?���4�w�Z�[5xy�)$�^���o~�׫��g3��Z?xq'��	��7����1V3,��3�
�o(�;D�������m�x����a�\�~Dr0y�4L�91Ta��.�3i�Qv{w&f@(1�a3���+L�6�^���N��p� ���̹�hlh@��� ��ŋ�q�F<��S�	��K�/d�;;��jB*��1�!�� eTf
��k�#n��� �G̘�ۍ��@�&���c鼠O۱c�?��T�>��(AΨQ&k���˅����ɒ�z�]�}�v�>��Y*l7��Lx-�����˅�<֮����ȵ]��c�n���o�h�PE�������yy(�/ �B=}�::� ���b���ôIS�k���rQ��	>��	��[��\L��[1���<���ۏU�v-�����i�x���.�g�K��&�NH�,l����k;���w� ?���S�Φ��o�����`���&�K�����U|�*(r7��vj_�ߍ�O�
�����[��1o�h|\K�*"9hn��w~��N^ŏ��2��s������?{{O�<��u�����`"�dvr�����]TЬ	c���hn��s�K����g���'��6��k�jr���tu��/�{3��sA8���;�0�sHc,S�w�s;����Pt��xϭ�%��QWW��^{Dr02'�K�� �"ƍ��������chooA$�<�VvM]2331���\^U�+���>�	b�����u�hnj�l�����ǃ>��}K����l����ylJ���1�n�A�A�����y��v��/H�O/�2P�|�*�ta�qB�)�y����n��W����$aڬ�4m�����v�0�DH.1�5�]ShJdA��
�QP䬭��(_"0����v�A�:*�D]:'l��R���k�"pmαx�=�}��v]�>�6T���O��|*b�ظ�+���q�����=}���ܼv���{�X����`KAA,Z���lܮ�@k[�(v�a>{|y���a�(�H.O<]������D߶�1Z�vA�Ο-Ͳk;�|jJT�L�,����	�%?#�N�Y>+�v����B|�k_�+/�����7��g?�Y�?~H����b���`PJ�˝�mOc�*���

�-�����#��qm:"�xs�9��^�_���1k�v��?��P�L�D�|p������X�����a��2�e牫���_������7��BZ*�JI���q��m<�?�_��Ӹo�$7�����ĥ[w@�3XR�Fks�32C
�������f��r��;L1��}�@P�.�/.�i�!t�v?�楗^B}}=�ÌWV�_����P!;+��C�;W>��}��� �BGG�9�~�0q"�_�=}�8s�<ZZ[ACw��k�`����%C�SSS��_�>�lT}x���hc,���P�7�"�9�A��A�;p�Vy�#��]��)e*>0%����E�8/�$K��~�|�M\�v��ۓ���QX�l�dM���r���AA��7�k���}��� '�����k	um��G�W�O(���µ]���=��A\����K��z������)���҂㇏����L�F`Ͷ�sa鲥�5u:�5֋�6?X�D�)
�%e� ި��%̵]"��$�GV鶰,ngI����xq{��5b�<�|��Ua���*�KKp����!gÞ�/������>�6�]��*5Ű^�T�)X��S�ۺno����}�����Mk��Fa�4T�� Z,��6��)�5Y{/n�H�ؑ�Ă��s��o=�ov9RB\�N�9!��˻��&�C����/����O��>��z`<~��G	-���ǎ2OwOZm��%& ��^�o����礶�u���K���������z|���Iq��t����>H���`�N�uQN#�05��ݩ����b&x7�����'�'����vh1c��dro�~nܸ�6�H��Z���`�ݧgϘ�����؈c�F~�dn���Kzz:.^�ޯ+k�q��U2u#=#G�`��R=p��y��W�裏���hH���TQ���fc,���e�X�d��@H�>Y=х��.�[��s�\���b0E�/�k�!����8-��}3����_~�^�� &�\�~�:�'z�vN�n��X������]�k�v��vH*܁�8\����ܲ�]1�ת�=P'����!�G�O�D��mM>�յ]~q{aA�

��vl݆��~D2�\ݏ>�~�>cF���Ģ	�]Yaȗ�v��[�{ty�u��k;�ñt��pm���F1:�SX��)䋽�]�ϣ������k��n]�n�����O����(���|��x�'0o�<
V!x�V���ԃb�UZ�S���Yrd`"�^%�c{�^�Y��Ld���u�[4�4��C�wb(���oC��w���M�Z��l?	;�����=�o�;����()��d�����:�����@����ϣ������=�4"���:��O�E�c�����?|���ͦ������C��d����_���S
s��l@�W��5[��濼���^����O�pt��م�7��K1�-'0"3]�j��kUu��ߢ�N�R4�����:��D�.��ٞ�����`<Ÿ(��+O2��t?���/U�ٴ�4�f��b���<�.���|��6?��ΜA$]]]W��EEx`�Z4�����b03a�$ܭ���+4K��ь����!�F�X�c�rm����1��d��$H�>��C��< ҉A7͠��H�Sf�*��bD�-�>�c���o~�ܽ{��)�o���K�޵][��+� �tm�nle�vU�l&����	�?.�G�.
�9=#45�Dr'�v1ݪ�=&��|�$_�\۹�R_S0}�4�de���r�ܶ1)�z7o���#ǰd�Rd������T��C��M���=.��ϣ�)��x��C�fq[X�C�̊�k{0yyѹ/M<��	�}k�x4���{��v]u�y��R������_~���N΅M�����?��e�y������PdmH^�\R�a���`�*��B��j�F�{:i�NU<�������KX�`�asm��;�۽g��p������b�K���{�ǌ4�?r����7��i�t�Ld��߼�GJf�ϾxM��D�|t���>U�K����. #͍����w���k����u[�����g����ϞT���0����Vձ|(Q^ۨ�K����0oJA ���_�����8���o��?�����gJg�I\.��>7�_wƹ,�g����{N��G�Y,�UdX��<���l����p6%���'o'�֋���jz�i���M�o�m;}_a�vk"����ɓ'�k�.�'wL�.^���>�������p��1455� �꒕��qc�b��8y�4��i�#bp��d��Յp6�1����#�#c��c�u3?��?�(XQЇ�i��� �� c��T�46 #C��.�XCM3ȋ� �T�.� ,z�*j�e`���
o��&�3�x6
��Ңwm7���K��ǵ]"U���%K�Q��x~d�҂Չwm���XL���r�JrC>�$� ��1�k��p�`u<�܆Ӯ݃}�X�~��b�������xu5b(��mߺM\���"gTʫ*����� ���O�	�=b��\m���u�z���D�����DD��n.l7�v��HωGH�.�I�eq�\@�������/�$�uq����qEޘ<|�_���
��9p� �9��+W�&H�?Xe���`���tc�
)\�t�f"w5�D����������`��/��U|���X<�	�\�U�7v��E�����N^��k�{��xd�����������32b����j�$A���{����U�a� ��o��U�e�{�syy�)ܪm��|6#GY�=|��E�9u�m���E��\��
s���^��}�0f$��:�ܦc�r�Y�%u����}S�/�5N���/n;��^z��l������X�h�.����3Pq�I���(�<��+�j�T�Z5�2�ۃ}�b�a�i[NH�ԉtmV�dro��_�}��/~��>�w:���\w���&��F��ј;c6z��������AFZZZPq�G��E��3z�^��w� �}�t��޴�g�F8�x�����rc��˥cU!�=]�C��)	 �� c����Xwo7��SR$��������|K����N4YM�~^z�%��(PǓ�;
�hѹ����6�]���N�-����u���ks�vQ�������-���H�G�W�Z��0ߨ�ET���C�1�c�iV]ۇefbެb4����ӧ��:��B��v�ڥN�[��ESǣ�n-Ztׄx?���C�֍�v�N���˵]�BrѺUq;$�,�k���|J�]�%�: a�o��ඞOvB��E����a�iy.^�Uk����πp.����_�%%%��@KJ�*�o�d"r7wc3ݠ_�n�B(`ev�x������o��T�GwO^�}F]�Ρ�ԅ �2�_R"4�n���^�"��O/%���֣��1t`��{O_S�������GjF�Խ=lߡˬ�P��l�2/P�C�W�fǾw�ޭ:��g٪Rd�A&F��C��Gc}�ۏ��~�P���8zT}�3w�ŵ[7p��M�`aD����
� ��9x� >�U�V���7T��y9��[3ƚ���7h0�S �� b�pZ�j���jY��r��Tza��yAV�[ě��D��֡����>g�DF+֮Q��d$�k�o��k;?�D�{�]�a.��"�%q�dP�~[E��>M,'�$7��H�I]��O����q�u������?{�[۰w�nܼy'NAu��ȁ��#˖-��)�PU[���V㵪��nE�܊ܵ]E7Ї�[��ĵ]��>�F�4I.�̵���c|\�u}Zt�L�,���z�ָ��|��y�~�ш��|�I\�Z�� ��޻w/z�!�Jv��I\��X����*ƀ�&r�̑������T59�AA1xpy�Ri�����.��=Tߡ�oȷ����<�����;���/�v�~f�-f}&�d��o�͞������7�Į�4ؕ��g���/�˴�����5�t����&`ʌi�WC�8��������$�˴}��G�ͮ�� �	���}�S"
R�������W��漠wn������[|8!��H��鼜ϒ%���������ȥ��rm���B�(c����9ѵ"��SXBx� �Ӌ�����C����E�\^�0^�gb\�e�T���GH��ڞ���y3g�|�w�:�� ��>~�8N�8��K�B���*�wt��:�^)T����1�Qt1�E�0qm�vF!n��%sm%nx>���vs�QU^��[#6�����G!X7�g��r��`>�ݽ���^��^����տ#��x�;t����0�3M\����*N9�k��{۵��SY�Ϯ~�������a-8�AAA��w�������0�?��v��0�k;'n7.|�=H���E��-[���ŋ �ͨѹ��x!b00s�L�8	�=��'O���999 �VV�.��������nC>����D�d>ܾ���ΩS����I��`c,���ڌ�8[C�XN�����n��~����.h�(.� Y�
�EA$8A�m�>��c��A�����)��%!����/�Doѵ]-�#�{���n���ź+�W�*�	�e�p�w]��z��IZl]ە@5![ˉ�e�7�l<}-��RQ<s6��{���>BGG�{V�:y
gϜ����0{��WU���w)�\�RخO�u�zL\۹�,l�p���񣜴��]����g�fY�.�g"���w���[�G/��1|8��������\.]���[����=��}�i�! lS��I���c�����t������g6ژ�Sp���d&� � bp0!�m.�i��l0�6�8`��O���Y"n7������4M����/��2g�Nu��U�o� ����&cƔi�x�cl;�A�S]U�.�&M§�[����q��5D����'���}}} ��/�K�[�iii�w2Ʋn�%ӷFl�%���c�ц�Ha?$p$����܉�����9q�4��P������'	�����_��4Έ�l,)-7�W���3qQ���xѷB���e�vY�|Zl�b{M�m�k@$��ω��t��Z�;׵]�}b\�� w'T���O�wc��Ӯx_�\�3s�S�8|����AD�F��#Gq��	u
�YS��Bw�,�iq��h]�`-�?�"y��ۚ��%�)׻��uH�Y�vm�ϱ��{�v}]%k,�5y��XK\�z>��	Ο9¹0��~Xm�1�┐��oo�5��U27��x�_h���v�Q�J��µ�Y�mE��@AA��d���p��i>��C,�}�f��C���ͱ�&Q�Yy6l��7@8�ťˑ���HV�L���i3p���ؾe+��έ[��eʔ)����e�v���Dr�������� �KYY�j���㏇�_\}��1�2�il �X|���n5F���v2Ʋ�ƻ�aѵ]V�B	��`�4���=�/@�n�<NO�~�;�����p.�w�b�j��o�:Y�N{lUH���%����[��[�R��.VS�򺛊��:���a]Hn&n7�cE�����˄��r�JrC>�$_D��2��(Z��#�9��P��Aa���;�\ձ��#h�i�"&0���C���ѫV����B�WV��G���!^ky�|f��X����B�"�ܵ�w�t�k;�ٶ��'V��r�
�#�+}7auI����eܺq�M� �	����{�җ�dk��,-^��xQ�)>�_� sd���)��z��̉0l��.e,�<!/j� � � �S:��u)����Rhq�Q<R�-��3�Pt��d1��Eymmmx����E�2i�L�:��L�03&Oŭ7�e�f1p؀4�L�6�{ ��]Ey�mD�1m�L�Vՠ�v��y�2Ɗ�1�|�2�"i7�����6�d�C�A��l7Z�� =ݚ{�!H�2�1�"���휸ݸ���I�x��g��N8���`T��w��V�ߘ��Z�+~��k���~�:���V�����u@�/���ta�T/
�4q� WO���;�x��i�X'	sm��! nl8���S�"od:��&{����o�>�U:֭_��a����Њ@�.�!(n�%�H\�%w]i�"ӗF(n7�y��C^+�v���{����ػ���)j������Z"�2|�|�o�����p&�~U���琕�H�;X�� V����Bw�w1h%�nP��q��.��A�r�{WW'J�Rq�6��EAAD��N����:ҙ� m���L�Yt��`"�El3�8��*V�������\�g���� �d�pl��*��7�k�;�_��.�s�����ŏq��]D2�l�
��`3:�;@8���r�����l���<-^���1�g�1VjG���)�		�%��誋̹]&n7��%�Ԃ0�ۍ��z������}����	���Ɍ��Ys��u�:��ت�\�E/J���<f�v~[_�@\�%�A��ZZwSq;_��\���k}�`5ż��Q��,D�lh(�|>�x���|@��O�0����[P�����3q��y�<tAğ��.�ؾ�F�ªի��׃�u�L��V��rm�܈���vA`nL���o���G&l�t��@d�v���E���s����1pm�y0m��}`=>ܳ�3�s��z�-<��3�V�`���]��Tƴ�jS(`��x7��`� � � �����i�c��D����B���?T��!�W�XųOO��Z������p.췺|�
�SI>A$ÆÊ%��\߀��w�G.]��O.}���c���8x�:;A$l���W�Ý{@8���G%c�c����l�_��ڱt��*{@��В�TՅ�ֲ�B -���l��pn������ro�W��`�u�|�
��OO�]�%Jt��\gYl���ĵ��R"�6�K���(:M�nȫ*7��3{A�D��.w�W�k��>�O�������뵥���_\��������to!hhh��M�0s�,,^���5hmkU�yL�Ӳ����KH�k��B>�Ԕ��p�vm���Ks7vc�Y]��!B�ɵ=�5������K�����3aS��_@vv��ݩ������f"w��]�� �vPk��E�j��E���h�AAAD22Vi@��m�Kߎ��w(k�	�7�6|�a<S3�ЯhV/�oXWW¹̞7y�� �d��w�.X�w:�݇�]D"`��sgϩB�e%���=u��� ��_X��g��+ ��ݻw���o�w�w(*��XVL��n7&�5�2A�	ܓ�U��ֹ0D�&�/�J���T����*�o2�%�.Nvo߳gN�>¹L�9Y�Y�f�/4�q���\�e"k-�~[3q��]�C��T�.�I.���Wz> ��µ]Z��v1��'k��>���n���F2�����;s�eN�A�˕˗q�����b���v�8V���(<7�G#n�l+Л	֣qmW˒
�c��$�ĵ]��Do�	������=��<nw*���o�?�	X
��f��drq�E�^į'��4��V2'��������X�xi^*�@AA�tL�q���Խ�l௹1��H ��d��0��3��8�o0Z���ذa�=r$��A$3�M��	�q��a՜� ����ݍCDNN\�5U�t�DÄ�Y�t1��Ԣ��:@��믿�'�|R��0�+�1��g7c��ZfMCuc�	ܓ�|ԣ�saH1	T�#T\:q{�i��(���`Uh�����h�ÄC̅�p.�y�QP4� ����L\T%��������PBtױ:y�-e���g��.y[�K���=$�vUyi�k�c������Q$e��L]�����8���]۵X򔉓0nl�:�zru!G���G���ӧ�z�dd�����>��$6�C��s�`�_ [�=K�"��+FQ} �xێ�k;W� n��.�Lخ�9��c0�#�=A��f{��������#��,�n��)ʟz�!�
&�ި$"wM�n�������w��.���B������
�)��C�B� � �H2���A���{�m$�K�7��"w��1�P�k�����HD�T�oy��E��d���a�칸^V�m[�� �ill���;0i�$<��~��p��o�p0��d�J�ٲ���
sq�w�ˏUc,m�gK�X)�����,ۇZ@�	ܓ�i�n47�I]Rn���ǻ��+����]��!
�<g�b������̙3 �Izz:f�-&h�A3gT^T(|�BA_^��:�/kБщ۹􁺶+!�n*n��k;$�C��k����;/�O�k�$���0��Fdaa�\\�pg�� A΅ͪ�g�n���㾵kQ�Ԁ����z����v.ђh[����bw��&l����Bt�$-�7&�v]f��ٶ����ۍ�ʵ]�j1�髩ٻ���t�o<� .�?��@8�z��w�j��ؤ�׮}[3�+�̍��R���lf�~��u�>�#�q�3q�xWW'V��ay/� � � ��47��X%�q�L��3B�ۃ}����Pm2��ݸc�z��_���{��{��)�4#Ff� �Jff&�/\���&�ٹ+�ށ ��s��-���c��%X<w=�ήN�������sq��y΄���O��Xc�I]�����-���S
�K�Bl��I���Nt��S))a�U)~��@�ʕ�]����S��� ��;�`��?���Ԩt0KV� --��/�Z͊k��R����Pΰ^'l��[J�إ�v��Zs�5�K���=$�QW����!��M�����.�'=0���E�v��.��M~J`|>��9�̜�t�[u]�룩m"Y�s�6��6,X��g�V�mt�#�ik��"�<!���$ك@���|>����O�k{�"x��v��]ۣ�`]���]�r�M���vr���?�Ia�����\����[����??Do/	v�V=������V��`����Py�˰�RGp�^��9��J��>� � � �H�Lp���7`����,�Cti���>�C,I!�@�7��b.�X��D���|��7ɽ�����#���T�[���G��G���� �{�:qX�z���Å˟� ���VU���=΃c���{�ַ�R{��$W�`�4Q���1�oq���f�}!���~Cf�UZ��A2Ʋ�')�.ݍ��\D�vލA�j0d��T�P8I�� so?u�gR4y"�O�����������8�Y�v���,�Nt.�˫$<�<��O�ĵ]�ˏSVnT��]w�ssFaެb=rwjkADrr��9\�z>��:ۍ+-��KEےm�qm��Fat4�u�>�m�yC
�u����#I�ۍ�v~�yyc���㽷��<�`����o~s����Py�#MB�2�����.�v�>M�������i�i�!AAA����:t�ܦ3>��~�3>���Ӻ��j��a�C���q�0=�fXx뭷@8���T�ܷ���������ƪe%�p�<�ܦ�	"�������{0�����!:y�m� '��뗭^�]����Cy���Uw2Ɗ�K0�һ�{ۿ}C,��V�o�FaJ��>4���=IY]�BoS�%�k]���]?� ��`U�nħR��Ty<�4`�.�3IKO�⒒`�U* ���M\�Ec֠��߫�=�ϸ�����E��Z*����a�Bµݰ_]����qzd�$�#6��&�u�\π\�ŀW�+����s��m�n��G"b`ttt`�ƍ�2u*�F�Fzj:�{����8½]M�=Q�n*l�P��/D��<�1"�)n�۵=Z(�{�哽���!B�,X�@oR�uq���V�Y�sg��z�5΃�łUYY�����|N	8E�&��h�Sd�`pJ��td`���Y�J�^hlG��htn5� � � ��L�FksC���%�+��{x3,��v�;��%}����TN�ӋW����F���e���6|8	�	G���-FzJ*vl݆��~��TVT���
�J�ctv��8�pY�٘�p>Ο:�y�1V`MXc,��P6��K����#���f��-�P�5�-�~�hH����)��\t#HB�0�����]t`����k�!�����i��4zک,)]���t�Z���Ep����µݤ���U�D,:L^��\ص������j�H��:�H�ڎ`Q!��Qsc��Zrm���--�/���Sp`�~
p� ���U���by�r������ڿf��*Ҥ�	s�(���=��`ސ�v]Fö�|�\ۅ<�|\���!M��״�S:�N��t����em�/~�+�ɿ���4���`S���;�`U��ݭ��/��LD��E�� ��@�"���y<-5p)c����AAA$�Ey=�g>�W�w(k3�	d���c��oێ<ɘf����6l �L��b��� '1&w4�-\�ǎ�qB� �6H�ؑ�HOOǂ9s�����M8��s�QUQ��;��t"d���	o�e���h�H��3��O�n��?@|�~lj�`H���f�F�\$��.��L(`X�
�E�􁪡����1�vr_v&�E�1a�$�D�m��-lε:��a���Q����e4��Ʋ͎3>���9�����^ʱ���+͐&�� z�v.��v��d�"�VW���A^X�j��m�0aV�^��;5�û�ޮ&��۵�5|��\�u�yq����`����K�2�����p!%��>i^�X�\p?fL>���`��A8�z��1b���@�N���G�~!�o+�wi��_*�0����}yu3��׳�d�KŉJBAA�sq� }M5 ��@^i[�\��"�4��v�g	N��3K���o�[��׃p.�O����=�t�2�vucۖ��9 �AHCC*++�?���g��#���A�{o_��;7mE?�&��\ܿ�o$M_aB�� mT�K�Whj$�kO��ZZk�w��>��0H���,ۏ޺`'��T���2�v+.�`�4P5t\��:�cǎ�p�iiX��DP{��jɵ=�?�vA�.���9��*���@!\�����|V]�5q����$�XssFa鼅�p�>Q�JĠ���ۨz�m���~�����j�\��4�ʟf�G.X7������d�3��vq[�$-(n7B���=Ξ9�۷�A8�z����կ~5�A��m +�����q;�'
1|�b�Jtd���'N�h�	d� � � ©,����.ddd�S���?�c���!���5��,-N�k477��7��L�/Y�~L�����q(�>GFKف�`��+�>u���XW�
e�7Q^qa7Y#�Q�`.�>�y���+��;c!l�ahc,En��}���%���XT����= 	ܓw�x�iLSڈ�8�0���]�o�A#���e6,ӐpI�r~�*e��k�O�΋��ڮ+Ǫ�]�wK���vC�%�z�8]�����D&�W�k;L�)����^[<}�\���۶� ��saؽkƏ�5k�Cyu%����qmW��{9����&���u�d[k�v-_���H��d�3HO(�ľ�Ƶ�b^]��|L����~��Sg �k_|�_P�-e8�Q!�i�����~4���M9h\�-��R(k?Tz1��sk]-FeNAC]+AAA8�"w3��n���C����X��?�T��� ��&����<�DRg��ΜZ	�;&�f� A���.�3�2ұs�1t`���ڍ�`M�J:~��iۙ5�U��PG392�
|���g�e�m̷���i��pi 	ܓ�Ņ�hom�0H:��S��ȅA�Qsw��c�v��y|��G �G��BL�:9�]�K�r~tB�D��C���k�(����I^@�ڮ��k��H�ٍi�pmgI#G�`��blݲ�UU���AC6��;oo��~}#�q��^��dQܮ�	�O�����>�u+��y*l�ok͍�j��`4��������jM��ྠ� ��ضygQQQ�-�w�'�x���Ĥ��h�� �'D[5���2���I�*%��r��������~AAA�cTf
Z�� 5-U:����p����]Z�~@�﫾������+���6l �<�o�d�J�~�����\̘0�.\Tg$bhr��9dee�����3�[wa���ؽi�p l ��6�R��=c,��=�1���0\���;lk����h�r΀���1'lH{�K:B$N�\��`�n��M���qo'��������R�tWn�@2����9 ��ӄ�~Kq�_�pI|9F��_"l*�/W�2Z�v�X_f�8=jrt���O�|�E�R�����wmg�3�NG����y�F5�M������͛1w�<u�YQX��"O�˺G�g&l��k���$Ͳ�]k������Ͽ7�y��}0����{�~�>y�5� ��k����{,���@R����wQ�z1�PfV�vw׋܍�7��2גAAA8����z��Zǻ�)��1�����=�)����x�l����x�}���s��1g�|���A���������<r�H1tiii���[Q��S&NƱ�'@v12'�����s�p�o��V����<�۷g�1�L��c��f��z�;?���=V�K��} 	ܓ��i
�j�v>H%��i�1`&8�waЂUZ$J��ȅ!NRݸq����)������;UF��/W�{5������ⶮ�N���:���!h�f=�bf!U�s����y��+G�)���Z���e����._ՕI����ȮI�n�z�xKs�wi���2nb{}}����㧡�W/^
d�����K6f`B�����~q�:����W}�ioo��z���]S�655��͛����ݭ7���soױ3�<�������.v`米�\kk�z���k�NL�6]��o�D��5hjl�_T|X����D�ht޾U����o��ʵ} u��>盽Ϛ���ЋDD��[����}�;���7�:Uܾ�=�F���9s��Ҋha���h�5?��o�����~<��pjp)�4� ~Ќ�;��.f�
R����Li-��5&����	� � � � ��.�Y�!o�e���o��4��v�_����x��> row&#G�`Ɯ� �����}�+��s����+#bh��GAaa!Y� =����/����媶�p���:}�Q2Ɗ��0��d�g�Qf>����gZ��(H��D�,r��ރ�4y�{��z��=���sa��D��7��8L��a㋩ݎ��*?'w�.���M�\�����ѣ%��&��H\ۅ-}�n^)Ô�Ӎ�T�b�������#pm�'2q��Y3��HC'|}$N�fy�\�YBխ��?��c��L��zB�O�||�Z�¥���'_��9s��]���s�k{Ѹ��_�}{� 77W]L��Į�������rL�8v����'O�����F�ߜ{\W�<v�˿{�.�6��`���c���SũEEEa�vz�V�Z���
p��RM�ֵ���S�9{&��Ͻ��EwwF���L�~��uƆgĮ��Me�~Y��	�++*1�!_"\ۙ�}��حmm��;p���{�y��ڈ�����:~�(���۲����q`��߾�꫸���uלSI�[��K�78����N����b"��E�����Ơ�j�������t���AAA8���n��4###Cp�sE�w��l��uq{����B�	��X�m߾������v'ۇ]��4��Gf��0q"ʯݐ�okiEKSܩ��&��1�5[�fq����4��<�D�?zT.��x���͵��K�m644��4��|�g�4v�i��~����3�rV�]�;���ifx��Xݎ;�>��[[P����P������T�]���R~2��	�'��{S$��;����<�8��6�����
8p �ׯ����d�e����3���&�Ҳ�Қ�1-w4�Փ1V" �{1������;1��L��N����O��6m�,�osɊU�.<��d���L@&s{���ԯ3���	*�%�Ac<�t+��>5�Dh*$�i"n7��s� :���Mq���Vw�7a��?��瓈��`1�1��Iqa��E�}�&v��$��{�9t�*�_}�ܮ�R�\$�,EģO3�{�/���Wo1M,#�1��ݷƚ�=�|V�޺�<o��V�������{���p��y�f!�9sFh���:&�{�4�����KQ�>h%�vP��nɍA��94�4V#5e<z��AAA���Dg�[�p��
S�s��� �1�T������3;�Jc��z�~�8C�8��n��=^�O�5��3]_[Y������D�Dg�gL��l6�5����h�-��y�(��{W.]��ڻ�t�����3���ȑ�8es&�����V�ف������9ոq�l)����.��ܳ���3fL���w��K�b��I�{��*���~�3�d�!6��$�g3?�߸U��>�w���<���~��P��c����+�`ݺ�ɜ��
�j��ۧ����PhCs�� ���ݸVO�X���I¤Qn�6�#==���nű�X�F�D&n�[=��������r�3y�<Nx���)�=q�\�9�z��X�D`�龅]*�D���bLԥs�v��㔉����cހ�\vi��ۅ㑉�}*���2M�|�Q�"x��S�-��m.�8x@��G�K�9�,���{<�Au�����~m]hni�-���
u��N���h]ۥi����NQ}�U�j�/��v �jM�n�������ǟ~o����~+l�(&pק%C�i�if��N���v~@w�@�U7���N����AAA�M�KAwc�|��žC3w�8@�_���~5�L�-���E��δ������� �EFf&�-Y�H4cF�a���8��C�g�$"����eTUV����ȩhhjA$��%KQ[U��8B8�ӧO�ĉX�|�c��`�e6[Y8��@{��kzݾ�Z���y�?10H��$,݋�:]P*Dp�J��̉!.�$D�JcS'���{ �R�_��Dܮ`K~�qrm��A|-�[��Na-���]����]�%�Y^��H�k�pm�y�ߍ�vݱI��Ӯ��� �ǍǖM�b2z� ��s������j�j�E��Z�z���%I���桄�j�GL���2���ֈ�h���Cɵ=��k�(/]��G��ڕ� �Ç~��/bΜ9Ip�E�Q�΋��-fA*��g�C��f�AAA�ݬ.b3M��΀�����͍���ji�~B
d��x���~Cso'����K���
�H$�3faTV6�o��=� B�钶mي+W���W��� Ezz�:H���c ��f������������\�.���ٞ��nf��|\*�T�7K�P��IBJ�]�&��Q�n����T���
��B�mذ ����epkA*7s���#{ ��vA���Z�ih����vIݣum���`]�ײ�}���@�>_p���>\�(�7�$����\80q�@(�v�iάY�i�P�A������<y2V�Y�k�7}�$��u���|r�k����5�_�/_�I>������i�{?�;O�?~�o4h�Ah�����4������~��+�w��]����	�].�Ck}-r2������ � � �%/��n����)�����b}���/�HD�]�ģNgΜ��#G@8���0y"Q��a�e��s��AD����Çav�l�[�9Dg��1e�tܾqwjjA8��{��ҥK(..4"v�iF�����Bd�������R��f�I_H����FG{+�32MU�L5ȏH��Z1Tm���n��� �E^~>�&M�}�\�}zf�]�_�lTm��
�u�"qm7���#K�ב������-��k����r�:Q���������]۽N�%K���Ө��AD<�y�&������|w��3�.(n�!�4E�����O�f���{�m�H�v}M���g��ĵ=q{l�o-���Xǌ�Ǻ�Ǟ��@8�;v�;������ޗ�(�N?�����V)-����]?���G��B��� � � �6Fe����RS�B��[�7�������/�^�$ 2� ����/uz���Il�0�oq�rD��H���Ukp����׃ "�|r�����u`����>C��'�J�aצ�����4c�������#b��1���=E���$��@ߡ?�����&���ڃ��I���.t�����*E�2so���߅�N�����q��m΁����,��ٿpm�8���wm���q���Ţc�ڮ�3J�����9��#�Ӎ	�m���\�M>	'^	Vǣ�m8�
Ffgc��b�ٵ��� ��'l��o���yX�n���	��Y�^]#����,�ڵ=�zE ��k�l��z '�CsS3g��Յw�y���w#N�`L~�`A*�~��D�M?�;����r�6��`����ټ�@AAa%����+!�ۭ�bE��]��=\o^_����fR�\	g1k�1���Â�s�k�N��� "444`��]Xw�z\��	�6�sFb�외z�΁c=��(,,�z_N�So��~
c̱,c�wpWB��9w�Ѕ}�zA��;����m���B�a��~$�o��26��Ȳ�i��{��Y�(���#�ߴ���xKP]C&lק�E��nاt�M�k;/$GB]�E�;`��n̄�\ۃ�����w#C�+�<a�rr�y�&rc!"a��۶nò��1y�ܮ�����z�x�
��|��O�f��鶃׵]��t���f��|rzz}��x�A8����<���|�j'�dt��"bB�4q�<X�;1(�*]��d�\�Y9�n�AAA�d�5�C20W�X5��-���u}���ZbE�8��/Vi6l@o/��İ��1kn1",�7nO
�n�� �xÄ�l0Ͳeː7:�/] Aě9���-t�w�p���x��w�G�G��+LL��Q���3�c��!ۺ��o�+��{^
3�"~����,�Fwk���	"�
A��봗�D1���U��
�$`�C(�-�ĉ8s�琑��}����.�A�@[�݊�vٶ����������Q_m(�/DV)-��k�I^K��(]�ż&�<�|�pm�pi��d���}�i��-�� ��U�}|'� ����㨮����vu%����tc���$-J�vY��|�qm7����<a���&N���!�-X�G�Ƶ�2΀Mm�e�|�_t\*�ei�Q�7-`�}6����~]�"P�:1D�.,��AAA	�0+-�u� u���P�wy�v����B��=`��`\G�o(�?tj�_,Қ���y�f�bQ�R��$� ��G�)Y�[�n�֭[ �H$L�4e�<�v=�<��>2c!�Gjj*�.Z����pl��o~�៵h����iA�?}�>����2w��tHM.7����FeNECG?��@�;�31��.�(�S/H+����a��d	DE[>sM$�fg�`�b�ݩ��o���BP5�/kU����ص]1�D���z�u ]^�ŵ]�7�`�����vC>Swx;\۵<BZ8�vv�,]�gN�DMM� 줲��>؈G{Uwj���T֠SG*s�0+���۵=�ےk{D"z]��������/<����O�Yg���o�駟���������ZV��$�̂mU�J��n^��$.�������_�{꽥� � � "�,ۏ�:]Ǻـݐ}��6��s� r�(��͈W���B��7����s�/,��	E �x2|�0�[����C[[� ��ƍ������PE�]� �x1y�T�,��{w�p��߾};�z�)�	���W)1���C���������ٟ��]���Bۯ��$pw0�n��� �`�5q�1 ֽ="�&Ó,��pTTT`׮] �Cn�hL�2% (7���=��Y'h6�KU<bz(�v�X^�.��È��b��.�ˋ�aP�&l7n�H�D�Ll� �v���ŐU_���4�,Z��{����,:	�p,`�����㏣������
��v+�vc>���\ۍ�����s)��[���[�ApA������;v,V޷� ������GaݺuI+b�4���B� ��o����e��pmg��-l��؀)��p����'� � "��uԡ�dj����B{�Z�ڦB��P3��	
���x�/��������ouq�2D<�;K�������1� �inn��m���C���3�oh AċE%K�{�v2�u6l�O<�����Kop�����Xs,����9��)���K�AM���.����7D| ���)�B_s��P��.sq{�O��nezAх!<��
�ƂT��� ��=.YQ���=2I��k���a�w��b�mF�/QShG�ڮ�7�B�(]�un�>�˫ ����+�ε]_a�����o��������9رu]�A8���wՀ���l457��Z���t� n��]ۣ���A�e�Ć�Y]"��E��ȇ�k�,�C?�S�O����3x�{�3����b�2���*+K�`�b�2L9�sF�?�7��� � � �2-׍֖fddd����/������Z?���e��ϲ��ݫ:��az�,d�$Q	?&M���c�c׎�$�#�1�>Ý�w`՚�(����JD<���Ŕ�p�Jgp��%>|�W�vP�^|�7��ͱB���K��6��̌��Q42Md�H��`ƺZ��rK;�C_\���Aޱ/����H�D�CɅ���]�f�p��OC����tm��D���)��R�9/�W�A����!/X7�S&�WT��KC\�=��uTI1$j��g�1�T0[6m� A��ݟv�܅+W �`,���	n��5sa�>M��]�%"x�h���/76��Q;�'�k��,9�6���g��[@8����˘5kV������1���Bwq�A޽P	��9#���zK� � � �D1?�]u.i�z$�X�@`����~	�dcoE����>�1�8���L/����f��I��?A��`�$|�%˖"k�\�r�.^��7��C&���w�Q�N��ބKb����+ |7�*��B���ںE�}�hH��P��S��xGuo�M�n�� t҇R�tr��t�v��_��i�&ܻw�3`��y狢,�k��z���#����k�V�G�B����J@6nH7��<"���n���W.�W,����%"x�x��E��n؋�OwP��L�2q�S\عc� ��#���x�̙7�5�j�(E�&n'l��(6@��؍��sm�ZD��H��$�v>���R50z����h�K��_�����B�߯�@k}�5L�J�&6�.�ܬj�m���_�wȍ� � � ���(��ܕ�b�3P	��|��8ت��8(Y���<'^��.��ѣ �ü����
��%�����]�]%�Z� �ͩ'1s�L��u��ID�IOOǜ�p��)΀c���a����ǲ|�1���o �X�L�MM�t�r--���[r.��Cw��b�OL]�M7�@�Tq�J�q� =�/��F;��s�=.2�3&F��.�������#qm�jl\%����k�>���ntO룉�c��.�'�{N�bH�;s6���� �H&.]���&ܷn-�S�tm����ѻ�G�w�G&X��W�/ŕ��>�(^��@86 ���1j�(�{����W~�aA*�t�)r�>ՠ,`%k��\n�ٍwR@AAo�MCg{��Tm�K��z p(3�@���=�dxe�o�������IӦ� b�w�_u.�;�ښA$W._���qx`�Z�=x��ND̙6{&�]��֖���۫c������.��vc�V���X6Ɗ��P�����{��8�3��IV� ���pW�"EQe[�eK��ܖ����ǎ��wt�an��|�ϳ����;�s��ZIJ�7p�DQ�DQ�	� �}���UY����D-�
x~VU'��s������y��@?��7��i��B�{�R�>���0�,_2��=� UR��,'��|�g��ӧO�ƍ �Ał
�۴�,��n��$~�r���VXk����v�~��'�>�l��;���?ˈk��,)�t�x�ܶ�?����!�"<��={�֏���A���z��L&X�������N�S=�k�;*{��N֯_����p㫯A�3<<������ T07��L���|����=]�%+�M<��9~L!�B!Yd��Q�N�FX�ܡ�jT�A��/�c	�9��Y��fk��ʺ���o�>��a�s�CM�'$e�exu�wp��qR�G)0>x��a����q��Q�ID_b��m8u�8H~����#jjj����K�M�c��{cY�"w���xl���7��d
��ڊ"�<Ei��TЅA3��I4�A*/��$R[Q(
ͅ��M�pFc����m(.N\��"k�k��Ĺ��w-�v�X�v��=^h�3Z*qI�5{�Ե]��.wmr���<��%΃];v���sx��B)d������g��ס��$�����v[��vؚ�ڇ�4O]�����+6ۮ���'�����?����>~��_'�w*l��OM��:1X_�'��I�w�[&"��ť��9	B!�B��X_fb�I�O�N��.�nu������������e�C�y�l�W�}���Z�-ES�b�I�V�坻pp�LLL�B
���~>p���uܺq�d������Ԅ�O���GL�۳g~��_�+�1��ϸʴdް(�7�\-M"rǰН5�d
��-�/J��l�%�T��|V�T��*�� ��H~d�彳�G����b�Xb0-�v�l��N�X>�퉢�]�����rm�	��2��n����Ů�xa���8~B�B�\`||W._���;046���Iq{�\۝������]۽�0�]۝hiY��/<�s�ς���͛�jS�w�V*b�����qA?%����čA��En�Bcx�%%"�H�k��j�ΒB!�B��֖bL������8�Cw��ļ5Q?�|��4�>���<`��;==�c��@���=��LR]U��݁O�����!��9Cq=k[����?0 B2Ŷ�w����h�'������/�"k䣁Uf�+��*�5�r���4k�9`�����#�ho,�W]S ���<dQ�����9H%��bj�'*���� f7�����[wn���E�u@�v�ص��ێ�%��$��rc��n��m��䳬���bb��w���Z`G�2�ɶ���կ�=Ч`������l�\�ni�k�Ҡ"r��,����D�
�vg��o���/c��Ey�����
'�L��M��C�����P9�!t�D�U��=:�$�����PB!�B�m�c+N�I�}�T�C�1���s)vY�I�:�X��m�l^�����q����`պ5�^TB2E]m�oڂ��|J�!d� r��~�-��?��^Fo?��HfXTW��m��{�6�z���K�={/��6�2���Xz�=(�1���.���ҕ���X���5S��$�P��gT�i��BII�+q�=@��`�A*�c�ʌI�nՃS�n���>��#��`��%hji������ۨ����w�M�vc�A\ۍMA\�ѹ���y<�c��y��%�w��5����Zk��D��a�vC/���w���O?���!d."�e���?�'o���؅|tl̼�ˊk��|�\�>w]���e޵=���=�������k����O@�s��A��?��.]��σP�߯�QC`'�>�L����>:2������$!�B!$�hZ�]Rw8,w�l��_Ja��r>�J0H]�m�1E�yBII	6<��d���&<Ӿ�����2��5q}{�W��W����B2������}LOѭ:ػw�.p7���XF�0�1�S�n7��qsw��c�Ǟ�Z� �9(p�3�o)�4���P�z}ø��h�G��2��L���ѣ�{�.H~�L��-����P�����̵=)7�#ub�	�-�s׮�qzRk��K�f����vS�n�gݵ=/�2  ��IDAT---��gw`Wh ����������?}[�L���H���_Uۏ��>L�%l7��&=�so�u����h��M/�et?���a�LLL�U��[��PA�<]�
��]wX�d����*M��v�2����XW=�/��B!�B2��R������B�']�J�$�5������=_h�/y�l��?x� ǎ��mڀ�
�	Z���m�n�E!sq�s��a�������o��q'I����}-��vD=���׍����=ch��'tw���9El����A��[��=���)(p�3�!�H\�|�}�f?H�ωA�C{�\�{;gg���VbQm��$=�v�Kz�]�e��x�Tl�oʞk�T(���P��rѺ}q���-vm�|q�Z�⎝طg/���A!�q?��{�����? RY�!�(���^��Y�g��=��h�c�/-+�k?�>>z���������~�;�	
*5��Tc�*j�ud0���_���%nw82�Vڈp�i!�B!�d�5U���H�^}�1�f3ƒ���r��	B���y@?��/~�ᇘ���]�@Yy�lh!�`Ų�h]�G!��u�=͡����zN��}�~��ٰenݸ�ɉ	���={�����=����D�n�c�'��$b�'�����X��uS���!(p�#*J�0�߅�H�+a�-lפ_*���U�@�C��08eE8��<yD=�ܸuK�U�_���m{�)nw�G]�n �k�mC q��Mqx]۝��Ko����Ч��n;�D�s�\���w���p��45c�Gs�2��>}�!^}�UT-����`V\�eq�˹��&��]۝�عk�9���~��'N��W^)�A�p���V�_��A�V��g�'�˖tNH����{�B!��QF��+�%� �C�Y�f�%��r�����wOI��g��S���A��lIN�'$U�`I}#�suB�<���I�|~�~_x���%��X�q=�]�D=��~��ߢ�8.	Η�_:�M�3\�/��0��rs���M�D߼t�7ւZ��@�{���с��gwxT�]��.)��v�`$�UKi&��P�� �>��LMq��|`պ5���,��I��-�"l���K���\ۓU�Ɋk�Dt�ˢk�=�������nۃ-N���sm7��[7nƉ�G���B��>|���z\�><�ؚ�k���eB"V�HGܮֵ=��`=�>�܋$��o����
���"�ֲB�
��Ml��<��]�O6����-�XE��Gk��M7!�B!$c�o,���0���m�mgc����4��rq�b�s��B[���}<x>Qς�J=wHH��_��zp��iB�|���s�ȽdU	����k7��ͯ�����Z��oGG����#c,�5��Yc�'�k�m����K���C���1V&��=�h*�H�ؖ,���v�s�ҥ��b�l�w�C���a�����G��G����v��z(�vȄ�]�!�D2O\�M�e�RѺE��Ի���q9\��KK�u��۳'�u�B�"�[o���bhH��WSq��h�8?q{�D�����`�v���׵m�v=tO��@�"��ݻ�+Vx�� T�A6s�f~�����1X����1�	u{=!�B!$S�/���ӈ�D�$ͽ�vc,-i��7��O��웙�.w?�I�s���#L~Q��_�6nۢ�߄�C���(ӊ���#cB�5B���Xݶ7o�!�E���߲	��^ Qχ~���1���c� @9!l׵��9Ck���_�\7�;} ��<�4�/1���5He=�]�T.�T�]9�dKt��:��C8�vQ���%l**�ύ�&���E�����um�}�o�og���]�>�vm���\��m�曻�ř��D�L,���q�2�vY�]����f����`����d�^LOsV!��]���[XPQ��1�L�L���q����44���{���gB�t���G�"�����?�D-b��}����ì��E��=�~Խ]��`sd�LO%rO�1`e]3n�p50B!�BHf(��������B#?(q�2Ɗ�t��š=S.�n�3g@�#V|^��������*���s�A!�x�v����Q|{�6�-�֭�7׿����Z�;�G�����3f.�N��F�c,�O6����&�֮������D�[6�k�"����=O��R��i���H�4�#��Y\,N�A�t$U&q!��l�<8e��O?�C ��6mt���X��r������>����ԉ=L,�Y�vY=��>�"Ϋ��W��h"NK�h���g~��6{��G��%��-).Ƌ�=�=}���@!�ξ����O��/ޣ��zY:��a��abú��#nόk{��l��{�fGp�q�&,^҂G;A�"���o�F����B����hbl�N���ܯ�l,3�pc�<#�n��q��B!��6+�1<4�����vc��e�9��W��&��`���՞�e{�졁N��y�V����Xֲ͵8}�!���9}/��&�&q��2�}��-�q��4�Z&&&t�;�7,dw�p�����x-�/Ku�!W��EKU:g@҃�<aI�F�	���%x��̹�)�U�]�.�n�C�_Ygg'�?���½��L����yn-2��<�mv#^�(� �(ϴk�m��`�q�qm��M���.�w�m�pmכ)qm\e��8��ك��"�b�ھ{?ޣ߸Bq#���}���w03����������26[�����;c�9�7�������Z<x�;��޽� �f�s���;:����67-�CR�n�2���u{-!�B!$]��Mc�ے7tN��zXr����9�@&l��������K+�}��' ꩭ����A�lYҼ+Z����	Bqs��i|��W099�GO���кz%����@�"&���w�����|vgϥ1���]�W�����a��#�� t��	�y@$�����r��E����C��.�Q܁���/*�r�̰o�>:=��%�X�a}�\�MSp�!��#^����G%���}Kc��v��ZM��]�ĵ]K~�
r�ڞ�b��]�vK�%�6Y}��Y� n*^��8��5	!�x#�����?�+���X��q���.ͥk��~YdỶ;i�ݷ	� ��X�J܃�矻B�:mw��*xRe̍�)2�=��RՀ�A��B!�Bңd�ӎɵ�>�<�|�g���*�M���0�r�'N�����AԳq�2[�zy+���!��q����꫘��BwO7	��;lxf3�� Q�͛7q��y<���y)JOEƌ����c��E�r��Wfh�`�/րj����=�����8��+�K��]���\�Y%.��@�I\��R����s�0��6l@Y½=�E؞�v�����#�����k�`]�k�{��$�qn��S�!�k{B�8�t]�ݓ����]/���C!�������������������Wn/�����\���2lW|z��0��vmڀl	����o�����<x��O���ڸ�x!�+������ʍ��/�����F�1B!�B�cqUC��(++��z���'��V}����̱�h�G�y�l��d��� �YTW��eKA�l�]��׮�Ⴧ@!$5G���?�.|~=�� $,��Z��g�cr|D-�?#�A���X�|�o_ؑ+4��F�:���e�gC���ۍE��762{(p�V.���x$� U½]���s`���w��"��M�th�C�_�x7n� QKqqܽ��"nw���\�m�rm���]��h��k����|a�S��vmw�W=�x�-��v�:a{�˙^3���o��-��k��j�x�{��8q���!��azz�������:�cj:�<�k�v��P���ꚳ����� �{��^__���u���������^��
�vc��RirQ�ǀU$��Ë���P�/ !�B!�̖����POQ����?��#j�ի�} �����3�Y�~��B�%Z���ѣGAԳi���쨩���m;���} �q?t���x�7�q�,��B�a��v�"�Z����ӟP]w�1�\�n��W�,y���q٪k[k8z$(p��F{��x������q~�|E�H|�-���6k.	a�9�%�,ȝ�*�PAii���%%%���&<�wI��TP�%u�6�
m)�c�����zLQ�Ġ=4N�xow/����T���񑆛��+~@�O���_&�����>�"�(��2��m������K��S���e�[��������./���q��m�`rrR��/�ѿ���e����X�;��ק�~�Ǯ�~q���K�7G*�]|߆��155�����!���a�O��B��v�j����]>p!o�$���gltT?��]O=#�n��0����8~��_d�}�W%��ݻ8qԲ�n�z�4��`4�����A��2�os�!p7�WQz���0�֍�.�X��VC�OQV܊��|�!�B!s��� FB���XEvc,�������6�!��Bth��Ǿ}�011��o�1�'��U}N����n�8�d�W�T���ÃCY�{|l%#��Ψ�ǋ�Q6�Ϸ��9>1>���,�����,�_�۟=��;>�hEh���:�s���+\[e�����8�t��'ר<�D�Je��n��R5���;/�=U���;���^x�E\������W�[#�.^o�@��|]C��[��F���!�Vy-מC�����y./�ȶ1�������n��}�g���9A]��"B'�&>W��]1-UE�/3½�>;$�R��A*����pHN}�g?R�C�D���\���1!��'U������t�/>�m;w���~��n�� ���t��(�m�W����_c��u�*�@MZ��vm7�o|�%�n\����-ǝ2�2Q �޻u���(���tm��/�V���K���M�b����X���[�n���*�!�ljjRR�ݻw�b�
�B��U}�B�.�����J�Wy������;�⚯��.+?~�e˖)������G����w���\\��:�=t�}��@�ziڮ�w��t>|�M[6��cϳum+�����r=7��ux7˄����}''���؇��Q��{��T ���O��;w_}�����X���:g��`���1h�����ݱܠ�������~�f�!�B!��)/������D��J�;��~�v��A�-V�<��5,�6a��KA�!pW��?@+�Z1����q��+�
���*���~����ֱ�s�}�j:p333�qB�j<Oh�k�
��]|�)���B�y'�s*E�Fݪ�*?{q�&p� [�y��E����l�T8�j41�B����c��PW]c}rB�
T��}4�w�0�w�|sg����ጱ�&��D�F�:����?6Ѕ�e���etޣ��4��ڄ�2��e
">_������.���> �@�ҽ�(4�z�xq1W��KL�nܠ��uٵD`����v�J�����qM��܆���&M+5Z���g)lO��%���q21z��v�g� q��l��D;����L^p��W���T:dB�\B��p(vo$Dڏ��$��A�".Ll�B��;̽�l�~�*D�A�J]^o��y�N�m;��'�Q��^|��'��]�-�P�^fPF7���=a�pn7��81H��,��6n!�B!���ٖ�D��Y��4�r&�5ۄ��#E��#Ih��kN�B.�/���+W|����XS�˪@���Ps�8�d�/����M�^���4��`�"�!:k\ܬ�n���Z��?�.Χ7^����h}}����ʌ��6A����FI�Kձ�C�.��T��؅�Y�Ω����1��ÙB�g/�7�~q�*H��{{z�׿�5>=zh֓��d��%���������v���U�����\��.�+�㩼�����re�[9u����[�Z�������{c�İ�ޚZ�)�1i���=���cc��\�K�j&���qU�A�El�o���e��Vw���$�A���`�Buf���O?Q�����L<&s�tm��{	���b��y�<�k{ a��<}�voa�۝��{q�g�f�u�y�����I�v���764�~�4|~�*!�d�����K���ft��J"��{��ҵ�u�y� ���f��v[Que��˗�@cS��<Q�޽{�����U
�]!l��:��Ӊ�շN
݋��UIa��/?=$V�R�&�B!�6K�F0	�7�c��v3�n��Y��*v�2�rR(����b��\�ۉ��۶���|�;����S2!����s���/����N�����+׮��s@�!�5B�w�w�m��?̶1���՟5ӈ���]��(k���%���
�RQR���2�^��R7� �u�t���]�m_z��P봐�%;;;q��Y��n_���2Gi�\�=��β<um��~Y=q��+.*�ˑk����5�,��;
��.X�`!�5/֗�"��y���+�TWc���l	�d86#����9֜��=�^p�#�(�|�U�����@�����>}/��r^*eӍ������4.�w�va0����`]C1�~:B!�B	��E19�n�g�t�sf5�r����Y�B7�J/�e��hD-�eu��e $/>�<���s��N!�������?�g/Q�L��x�,��+��cϞ=����\A#�g�����c,��"3��9C��>&��@f�
��R��Xf0���I.��� �]�F�p��}�߿SS�D��½�JP��x,���p��ZC&\��(�ڎD�!������k���\��C7����f�����,�i��̵]<+-)��͛���BH�8w�ެ�ח���J�޵ݽ�t�Ac�µ=��ƥ�y�3ؿ���2��
�]9t�.p�m�ww�ٴѹI܃�rN�^9ͳ�.l}��M�� �B!����o(���(�+*��&��Z;S^	��&w?��\�%?~O��3���MAH6�mG��.}uRB!����{���ĺ�k���o@HD?E��.�9���y�]�vt>0��X����ٵ�=�%:ࡁA�.jƝ�i��Pஐť�-�va0g�_"����V�T�`mV��6>� ׁtVM��UX�pa╗k{\�l=Où���]�����;��C�ni�G=2���k�����<]��u��k�f��n-a�Kvn{��������c�����&'019�,O[��]�%�ȵk{Z��4�P�Ov����@�q��A��?�3����ׅ�0�x� �n��rR%WK�V���K�M�I5 �B!�������d����qc9�8V����X��Su�
E�tG�	��Y**`Y�
�K�cay�]�
B!����_⹝;�t�<x�	E$+׬��Ϯ�y�D�F�s��]�m^c!�9��h���֒���+?���ƺ(��nVP������S��s��t`p|Y���2w�A*#�Z���f���_�ڵk jY�q���ߵ]s��;���;c��칶�c5�vm���]�ʹk{"�ϵ�-�w���m~�s8r�0&&&@!$����{�����/���}rQ�"�,��{�!㱅��&v�Ǻ}��� Fu�����!�u�ʫA��1x\/��E��;����Ace����@!�B	F�D��\�<��˾J���;�I~Y�P0�L��e�/}��Q��vq���:�-]�cG��%��\p��9����12:��~*5IjDf��u�v�
�:��?��?���B=o����X��Bg�ڜL���=$��3�Z���wEll,��ؘ{�A�A����t���ͅ�21s����Q�4^RхA-KW,â�Z_�v�.�*���)�����-�gߵ�v<2��,=��(2��E��f��C�[\�5��C���m�l۴ϝ��� !����i|��x���
�:H"�k{�D��(�WZV�_~I�5�����{�x�B��ۼ���s#R��܍�4�
j^KFl�֋��	8t�B!������zQ^^.u}�2�*J���X���·�ub�Y>1Z��A�xя"w��Ҳ2��YB�P�^�|f>��	!�䎃���;�ctl��bM�Z|}�:&id����nttt��^��|`&���]��c�&���]���7������nT�Uax�ZհPஈ��S����`r ��E�����Rŷy�[�(g������C�@�Ҿy�[ܞ����8��947]�e_o�{S��[l��"H��u�A��pme�˗���C<~��Br���0؏��*:�'JC܋e���c��X��gBp,������8~��r��1������N]��
�ۼ�L��Í�ZH䞘\��
����U�@!�B!����o�_5ʚ\�c��� �v/�, ��ݗ|�E��Fc,��Y��Ŕ/�Ԉ��+/}��}��-!��q�=��~|���c�ჼ�����b������uu9rD�!�=��X�P�1��c���c꠫?M�d�����;�Q:9`.3t��s����U��KǺ%N!@�&�ҥK�w��:����d/̩k�=6�k�D�n��<��қE�b��2�hx��)��k��m�]�5��XX^�Kg΃B�:?z������U�����ڞ��wx�y���4ڔ�Xk[+T`���q�����t��������2��׍!�|���KZ����*�{��c��m)�9�O!�BIA-�0�BT0c�p�v�>�$���ܝ*�e����ٳ �����ׁ� q�w���@�BT011��'O���_��3 $k7�Ǎ/����4�>��XUUU���v~/�>f�=q�縴�2�;�*r7&�['�k�O��џ��R����a�'���RC}=�%�	�\�ܽt��=.{����P�'���h��`�̳a�f�E�\��%9��v[,��z�f���p�>$��QH�y�㊛�k����0>W��Ƀ���������lZ��!�����+XҲ�e�7����ӵ]��`��ڕ���v���';033�C�n��B�t�e�T5��A]�+�I=�*mcc�X���.&[	!�B!�Db}�сni<�1��oc�1�2����Jn�/~������Q�ʵkPV�U�Hj6�߀�7�E?!��C� ���lX��o|B�(�����m���M5����y����yot�~�Q�>4��Ț�-[�����[����Oc�/	�
x�9���vG|��3@2�̠U��{?���L������-˗�_�Ե�^&��pmw��5i��k��===�v-�k�~8~���2�k���W��$â�k���۞�����!������/~�K<z����场��>�>s-"�G�}�X���E���a�F\��9�.^��G�����3�0���m��'OZ:��Wߺȱܠu����{����)\�!�B!�x����c(/����c���T^��u�w�0W��lݝc,���� 456�<R��oRG!���7����P_���� ďu�S��?:v�.p���*l�s�3��˱��]���l%hy�ݥ�D02<���b��1V(pW@K�(Ɔ�]\IrKR}��:g��禘� �l�O�>��<*++A�P�ؠ�ӆ��tޔU���k��c�ص]���U�+.�k��=�gQ��|����[����ܵ��n�v�ٖq������BH� ��}�!���?��G�΍.iN]���fKD8��]ۃ��˻)pW�p�?p� ~����B�}Iz�A*�>���]��`W�����ޫ@!�B!^�����D�՟c�e&��}'�ܡC�n�c!۹���=��ܿ�.]�{�B�j���j!�C|G�m،O�}B!�C�ɓx�7q��1LpE�C��4/i�㇝ j����n444����dB�1b��4�C����G��n]�9�)�E��������N/H(pW�h_ a������J��
�}���/���l
��l$��Hq����>�ʵ��!���v���õ]"D����\̵ۡ��䱻]���/�P� >|B!����0:N���v��ӄ5q���{�ҵ=xl����+�t�2<�wDN��_�>�x۽���`��Z��>w_[�ܠ�@�1X5�׃���Nz�xA!�B���M`&�Z?c,�jSAͱle-�3r�~�����W��]�� �q�z���qh?Wi'��|C�O>x�|�U|z��c��v
�bc�򗿜�X�9VPc,_m�Ĩ:̣ñ�+@�C�{�i��`hp@_fй�� ����b�nq��!vW׌���Ln��3�P�� �ѣGAԱz�Z]���Kݿ��黶;��Brdյ������kΥU4���ˆk�����ϊ��c.�DS]=��B!��ݻw��e1�����u\ܞ�k��a>���Up,6�}�5���/��������>�<��e�<c�I��N����^6� �נU�������>���B!�⦢�C��()-�:�K��i�e:��_��+Ih��v^�sn04�Rˢ�Z,��$�w�¹�g111B!����8._���}g/�!^�,[��j��������=����O���g���K��}w��l��OQ\�SL����1v�ȗ�%œ_���{�A+.�v� U|[�6�%g��g���ӧ ���>~�?ϕk{�ܚ:6���{���µ]3�����0˲��.��uo�������A!$�9{�,����(-)��d<���{�{�l���!n/t��0�Yrmw�nܼ�,܃��!��3==�O�����uW�M�u !��l�)t*n7K��j-!�B!�8��T��B8�iǸ�+<sp�jݥZnЯ�Ν;�v��:�lh!~�]�O=Aww7!��/O?Fcc#V�\���n�/V�_�Kg8B�ΝÓ'O��ܬ�V�Ξ�Xn�e_1ͽ�Zʼ�E�.&lnj*ƕGS ���=�,҆0������E�*�[\7� �񭵖ƙ���P�:::B�d�e�+P]S��s��.���n��=���"K���z��K��N�x@�v�_nѺ,\ۍ?a]�m���69�q�3�pp�~]�E!�0������/~�{��k�G�<.����\���⋋#x��p`ߧ j8q�.p7(�z����������?@�\%���d�z�1�k@=!�B!�ɒ��ޑ 9C�r��֜��,K�3�kn0SBw�^(V&j(+/����.�QW[��E��8q�B�k��W_{O�{�?�Bd��^�k��bb|$�LNN���w�y�`��Y1�
l�%�oK܃�#����)\	
�9DӢ��1O� K&� EfR=���R��z�,No�ʏ|qf0��:�nhϝk�ԉ�ܷT��ڵc�Q��Fyn\۽�SV����ڪص�_ ,_��n���� !�"	x��|��W���q�<}��0�9�ӵ]���۟{Gb�X�ϟǣG�����3W��M��3He�c;����=���@��&<�$NB!�B���w"�#ghwp���}����G��DC����|�;�����k�~4!2�ul׶طg/!�G��o��}GҀ�H��m�*|}�:�N�<�܃�_B�pu���ːǵ��7���&�Nw��jAVf+��j@�A�{io(���8��+R8�[Ov#����z�⽐j��B��2��T�/^�ÇA�P]S���by���ڦ	�ø���oE����rm�8�;�i���k�Ȳ?� =�����)��ĕ���aQ-��2D�R��e�:�?@u}��z>���E��*���=h\��JlںW.\�=bb�Hڿ��#T�Lݚ~�'�t�}�[�0�,+�M<O��`�R���A��!B!�BH�����QVVp�gs�&]�ٹU�U��]�]1�|������K�P�8wW�[B���/���GBH�133�S';����p��9"c��u��ŗ��W��ӧ��ۋ��:�u&rx*�~8M��ew���}hw?�����j�&YC���.[��q��A��=�����Lw$� ��%.�R�V��ևI��T93ttt��Q!k6��N�"�B\@�n�C���":w�:�k��#9$qR�vg=鸶'�е��[k+��eµ�-�w�E۷o�BB)p�����ܣC�;�vyd���g�����+6���θ�v��]!'N���A(�A+w�#����C���=�du�r����X�e �B!��-���I_Мab��)Μ|kN�5^��P���C;s!7�W��cǸҜB��.GyE9����]��100 B!�G__�c��K����� �ɂ�J,^�D7P#�gllL7���O~�W9����]F���Ksk�s�&X����tpO�7L����M��7	�
�sH�t?F-.n���.^KZ$���vr��`&�4^<?z�(����u�J���� �+�vHE���.�;�|��]o�!��ˤk�S�n��̵]r�b���M��q��ELN�B
���AUe��$Ǯ�i�3�ڞ��|D��k�]۝��[W���	]����3g�d܍�U�V2'���@U��O�.{]�����{����c�Z��B!�B�QW<���9CS�n:�Y'�5��rp�c��O!�S!&�u�n�{;�SQ^��e+ph�B)\�~v?|��<~������C��	�{
��ܖ�1�s�碤s�!rO��S�bELc얲QP�~J9����Eq�8��e�*Ѐ����r&�-��Q9`�ξ�^��;w�u�*��%�
�k{n���횵6��Y��[ږ����k;q�����`z|
���!���gddCCCh���Ӟ����rmϥ�<h�k�W쮗^�G��H��'����?�K�z&�vbݬE����N���{����B�>:�����; !�B!$���S߾�s2m2i�tp/
էI�$��jnЯ����ϟQCuM5��@��ﾰ�!������#X�d)�!�+�bxp$�����WUU��=�7�}e���p�����eyC�?o����� �
�s�Ʀb̌Π��18�y/Q`�������Dŷks>,3��}	��c$s�.6ѵq����:��}HE��x���6y��]���tc���5�µ�8f� �&n�����n;N�k�f��~F��C\�6�]��� �B�O�>���8JKKuA�A�\ۥ��tmV��}�XU��N�l݂O�����8H��UB��d�Z��`5��TԼ���`��U���A��bU������B!�B�ʺb������ܞ�Ni���ܽ]�:��E�2
-7���۸�-��ׁ[6l��W>���B�����ʲ�_�.���+�d��5�z�2H��uBO��of5痩��i��m�wHc,i[��Z����� W5���4�?����1=.wr�<�mU^.>�p�X���� ���u��15,��E}�1��*�������d��0��y��n��S��)"O�3+�vs_.Q|"*�<.�k;$e���'j����[���|B!s�O?����]��|�s����У�tE����#nψk{��\��[��l}vΝ>�{:::R�1�Q(�V�y�T�8�/7C��+s����]]U��Jm$��2B!�B�� [�#7��7�2�$a�mX�D���`.���E���������@��ښE�,-��@!d���ߏ��ZTWUc`p �Xi[��.�����#�����I�c��.��Ԙ�m�7�c�9B��7�)�9�=���AR@�{����d��r�0��b|1S�.h	;+se����۷q��5�oڐxfum���S0���2d�v�ݽO?�[���C��9��"xM�ڮ7��ڞ����d��ɏ�T�k�H�qI��n�}<,�k���˖,��{���!������4<����u=ql.X.�ϥ�����
�}�
�1::�S�N�?�AN��a�3Y���A��uҨ�=���D/q�&���ղ�B!�R��`4	�3�����Ͻ�.2dY��PyC��3���g�p\B+V�����Xמ�?�}{��B����x�7���A �ki�rܻu$��`�҂XYLP8+8�ۗ��6�[֟���l��L�|]�#ԗ�������-���}�̅A���pg�8ù��E�:�/���{|���=I��r�d�pa��J�J���-����]��h�9�'��b�]����Ԯ��mq]ۭm���g��n���n������ڞ���w�]�%m/))AK}#��� !��e�<y���Ge���$J�����YsmO������_�k�3nqK�._��������w'��
ZO<D3�UK�X�p���)n���	�Ep���B!�2ߙ�N���c9Bc�碐��3yo4w�$�s�~�¥p$9VErͪuk@����z	�;N1�O!s��}���z�9��x�XY�n-��E�p���91�R�t*c,3.x?;��u�߃���1��E�?����%��Fyy�t�JvBk���e������_ZǈT|����R̞�z�ЅA+V�BIi	��v���H{��C&X���!n��_�OO�6�B�`��k9pm7��rm7���gp��AB���8~����1<2,�N���vmO'��];)pW�����/��/(.���@Sf���[���T�����ܽ�����X@$A�"��@!�B�ǈ��b�p��3�c%�&�W{v��*�xy�6Zn�/� j�k�Ǣ:
8��%--���Eoo/!��]����r|M�x��467�zQ��Ar��3wٶ�d���򑜈�9�~�S7<<8�������Z=�h�D��7k�"dO&ӋBX���`b��O�X�����9��S��u�������ȵ�C�̵]V��8�vmw��)���,�����cȺk�}kC]�߹��B���ߎÇ�ŗw�Q�cK�4�c�H�wV���;VO����k���6���155�[?~��W�b۶m3�4�}şG��W��#��WK�#nQ��2������.!�B!d��^��:D�~Y�m�e`�Zͳd9�B��m����܉�֬!Vĵh��t�>B��\8?|�M|z�W� 6ZW��Ջ�Arϱc��?�)�G��z&����XN�v-�O��׋\ۼ������K������!�XE��*���<�U����Uk�)��~�j6��:u
��� �G̮Nq,bl�k���{yP�v#6��=jJ���ܸ��"x�{=�eڵ�������5mi�btp�B��=�`� ������y���.���-��xY�oYy6=�W.^�-��ELwٶ�hJ���V6P%��8��_7��[��2p5=,�Ț@!�B�����c���_��fX����/J�nM
��;9�V����v��e}������� �ʋ�=���N�B��@w�>s;�ن�W�"&��W����03C�o��}�6nܸ�u��e,��9�P�X��C����Z��L�n�6�	]k�7�gM�bt���}A>c#!b��C�-�cWI�u�j6��g��am{{�Ea�ʵ=�I���x�>�wm��%q�rm��އ�]���{���z�ҥ8�!d^r��A������%_E��(�^���;��m�N��"�[������|h�|=�{_�r����T�"��D���[c�V#��h���sp�B!�����H�+��3�:¹����=˰�]I�Թ�B��m;�<�X�b9JJ��1������8���@!d���ݍ�PS]���~"(�(G�t� �[D��̙3��]�mn�M�Mf����n�O�7L�����T����qq���,����(/��]n��k.3h[rPsX��pc�q��Q=���z�2�B�.�Be{n�6¥@<T՟�c�[Uu�>yj�O222���N��s�%n�z�L�n)��NNOIE�1��6!�k/��^624��;��l�v�L.��3<8��%mu�[�ڃ~L��va�B<�|�z������1���(�[8��ttT�(����$*�]\o�o�����cW]�������������=�8�T�?�֊��|�޾����m�J�x�9M��� z�{PV�>'��<�]$cn}�m����*�^������r��鍝�S!������p�z�.*���~/��%��c]KK��{�a�)�z\�[�U����U������c����� �B!��C�F�~�5o�y�ܭ��d�<�Ù3ķ��W��T��
��h[��XY������B�#';�Ə���C�A�AۚU�+B�����-��?�k�2�rN47��~�`K����C�}XTр�QcyA�{�YU3�'bqy3OV�lk�������ݍ�ĺ�d�X�m�}�?~��K��U���'�u7-nƂ��1V\�]\��{;��Qص]v������������!�����.DF���f=�����r�����>���Y%�~� Y��&����U�m_���_�^����*e�Kq�UU���MNN*=���Re"o�B[Q�8n����[u��^���.�s��{�$���_v�b���M1�N��.¸�K�SS�(-+Eł
�}z�7���Op켏{y�wVK�k����Ů���y�]f�����$�������o��u�x�<2��eg�t�DY�DYGG~�����@S��1�J�C��#����S������'�p!�B!����B��_�sr��d;ۜ��o���(�ܠ_�Çq��]=O!C����VF��&�g�Y]�dp��&�|���U6�2<8������q������7��=59��ё�c,�u/nlҍ:��ef���~ܾ}[I��H�����J�Wy���D��7*�]\g��OLL(�0v�u�2dS�ً���
�*��w�?�_����x�+ku�����]���*��W�;/Py�1:<���^�����5���Q&Ӯ_�cT!�s��W��������?׍�jk�N�\\�����ͱfk�e����iIM�|���=���Р��=�Q�2U��8��35\�Q�e�
ݓX��HY�K!X	N�>��$za�D�@t�Ŀ����V6�^վN��01��ş�']��]�8��K�l]��5�ㄫ��F�Q6��Bq��\��.u9�J��g]�aQ]]��Q�8��sm7%�	�{R]g6�ɣN��׹c�a�}[�dmw���m�ܾ׮|��VVV*�����j%u��1h��~q#�5h�����c����PU��cW]��]�`���W��c����^U�b�l�ʖ����q?��_�����2�ۼ�"tKaoy�~�ײdI8��4���?�޼��-�������o��������Bs�~/�!l7b��\͋'�<�m�v��"Μ<�tQyo��{��.�� �N�a�)��r��������;���N�n�JtT,�� B!�B��CLx�&��	r�6I�<p�0Er0��-^�"�s�~�'N��E�^�qLU�3Ch�Jt��c߸u����ݛ��b�J��񃇨ZT��Ʊ��L�����z���x�Ҝ�+ηm�7�??�D[[T!Ė��y;qݭ��QR��cW]��'O����_�@屋q⮮.,�<x� �/VfΤ���B/��ب��|�ο��k8s�FFG�Rw_w�~��'������z���z�0�=��_��ŗi��{{чƧ�{���>q_"V���<�r�nc���n6�X���9C����yC���e"��"�
ܳ��`�Խ�s	s�����BPQ�\�:u*}�	���^��:�I����wmפ��Q�X-h=n7v��^����z��}?�D�.�vg�E�u�%�bN���N��\��|_ض/�\���	��L!��$��_ÊUm��띕�<e��� 6��ݷ� qY�ͦ`=�8y�<VL�\�f5n}���b�"&��H��B�8Д�z�ĸT4�@���Ⱦܠ��]��><4��M��O�B!�BH�����܋�},Μ����;,�ܠ_��s�@� �	1���.�t?!��Ǐ�{���Ǐ�A��U����>��/	��l[>�g�����:������qq���JͰ$⢉�Xj&��g�5�%������C�e}q�J����Q=���z������ ��u�J��m
��o�3x����2C�n)����p��sm�Ǝ�8M��!Z���[��ʵ�^��,�|n�}�ڮ�o�����Ï@!��%�֮[��/D�vqgnE�qmOI�]�5!M�z�XQT�n�{f�3�+@�4q��E���y*F�]=n��M�9K��ܓ+���|���o(�ɻ�B!�2��[P����x�P�<s�.c��
R�՞���,S����2E�� �o1ћ���&,T��,�/6�[�_~�\q�B��F�,p��-�[�_�n���u����-�=Zqq\N��9�L�!�R3����shC�+?'�;����Pʋal
D�Ydբ�I�/wl�T9��!�L>�vb�#�g2�Μ9Î�"V�l�!w��hy�LH���n��B��[�?�]�݂}{���n�h]�ׯ}��
w!��9�?~�֛���P��v��s��&�����u���˒��=���K�.�wٶB���4�%�V�GX���:�K�� !�B!�����nmZ�|��_�|�9C��$�z���_.�Ο?�����C�vbPZR���&��!��o��?xㇸy��DDg��6
���ݭ�mݺu����+���Y�cYs������ ���b\��]�Y��dc�6o����J]�Iz�,��P��\��{�CCS��8���^�v[��k����r���K�s��no�۵�k�(?�Mu�p�!�'������Eii)�'��Y�g޵=�"�|um��՝��7��W�����J�/)t��x,�U��y��k�s��r�ց*�C��Pl�t�#�B!d>�T>��ሴ� �����v+�����&��B��m�3i�E�!��+���K;w�tG!�'�;N��gw���� dy[+�^��{�1����]��Ps�nc������Jهv��f{��;��2�H�KL��
ܳH�Đԩ�ӅAs;1���\N��`���2`%ܢϞ�M�
Z׬��k�'S�n-s�г���ƻ��̵]Ҿl����ݽ��q��ז��8s�!�/�>�����yx߾a.��k�<�����^�鸶;c7?��
N]]]hjj�_���l��S�b�A�q�=&0<Ћ������B!�B�ҩAL}�ܡf�1�ΤyC,g�О�O�;�d�/��iC�	�$s,^��ee dQMF���!�)�+������@�9��T,�@��f<�|�[.\�������b3Ghbl2Ӆ�P9C�������E��h��r7�g���';��봗z�/�fhXN����^N�r��5W�u?�Ն�������=m�e}\�!�K�M.q:��\�]ù.x.\ۭ�5�E��fM�%������j���q���ѩi��p� B!ވe��q-��Ȉ�y:�����gA�J��`�����d՚�(+/����џd���)�;w?�я�&e��!yg%���x�V`���pf���������r��B!���9��@_�?q���cY��󆎜a�r#�|���c����|�� �g��V"xa�N|�w!�/Nu�����*�8B��;�G�ń���j����zߵ��1V���]9D��}r�7Vy�
ܳD{c	�#Q�I�� y��~�ۉ��%;�ˀ�ŋ�L��բfѢ�+�v] n/�J��p�>$�A]ۍz\��ʵ=�xoB nۋ-�.lw��;�O��R��������8�̆Mؿ�B!��t���Ż��pm+8�� q!bϵ}��vQOqq16lބ��/��+W��w'�ࠐo���l�xͶ
��@Ź��ʚ(nt�B!�2XU_���)����'����2ł{2��4P�s������½]L�&����K�-!+W����o�U�	!�/�1�4/_����t���m.�9���366��.�����Dp�6hW:���������`[���߱�Q�TE�98b��,��2v��Ig\H�\�8������Iy��|��ԀեK�@rOۚU0��LK�ε]*��	̽�c�,=�v�@�g��]e鸶Ǐ=*�<0���)i����zt>x���	B!A8u�$v<���v%����е]�����U���k�m~f�
8u�m@'_2�c��r���@�UE.w���dc��b5��B!�2�YU5�����_�����p�~���}$���!���l�|�2H�Y�b"Ŕ"�w�5fM�*����X�BR�����7ߠ���%/]���x.��w'����˷����2ǒ<���]���kk4t�8`�2KTFG0*I`���w�v��yXќ�����$se�J�jϝ;�{ZW�
��.uI7�,����0^'y�%�V���no��Y(��d�A�C /ڑ�v�h�C ��>��F�ڕ+����B	�Ç�\��$�'����H΄�<G��h����cκ���,VVϊ�V,�����0H�x��n޼��k�zƨv`�4�];�۵�����AE��1�zE=!�B!s���8�Nm��;��^1*�Ê�@+{yðd;?)��={$�,ok!�m}�/�ЂBHp�^��-6���/@�7�W�R� g���A�[��⢽�%Ϋ��1	]�
[S,�(��2a&[b��,19�﹤�|v��������(��.^drPʏlX	��������܄+%�s�v�gܵ]&��/��������m��ݝm7۰�u%>�u6ru!�2w8|�~�֛���1HA�v���ѵ�3>����Ѧg6�ܩ3 �C�{\�pk֬	5��O��t��V9�����f�8��P]ր�q�?B!�2��w%�}��\��R��&��K��-&t߿OQL�)+/CSK3������e���!��G�aӖ�().�����e��e�����$H��ꫯ��ى%K�x�D$G��Ѩ��;�<ٯw�}L�l������P��j;�g���FGFP^^�q!�;Nr���\7��\�_0Gi�ǕO�R\f0�X��*����Q�`�.�v��#����)�w����
o�h����*,w9�[��µ=�'x�]����{e�8}�6!������)*�+0:6RD�I<[��;;�]۝�o�@����������<�
���s�sP֗��rls8*9\ܭ�T�ފ��P�s88K!�B�\��T����.�t�<��\}�"W�$P��P�k�|��}���������cff$�,Y�\?g������ �B�r�dv�܁�s��g"������� �C��Ν;����'s&G�M�?5��)������?/��&�;���PRT�IvamP�����N�Ay�k6�yr�N�K�n�,����By�����%Δ�t���3SHn"sI769bø�����%����_�m�;��um�	ĳ��G�� �umO)6�o��S �Bf��c��w���{�\�º�;��vm[���rii�8��`�Z޺��I����)�	C��K
�d�A��h{$6�'��.�^��ec��B!�2�i�� �n�&Ib{cy=��/I;`� ��s�o�����I�Yֺd~S_W�������B	���f&�P]U�����˲+(pW�0w'��#̬1���,s>��ۖ��L��\��=��=> &�k(Ƶ'\��
�Y��l�E�U�GQ�/DJ���,��]'��چ��a\�z$���ա�:�<��k��L��̸�����k����n�k_Q�W\\������B�l�����;����C��:��rm��l9�#Lh�\ۣ��p�*�E�7n���@rG__�_��-[�d\؞��Z�*�se�U��i��KZ�b��i1�c!�B!s�%�Ә�;����˛����K�74���>N��a.ȶ�^�5�+���󍋛A�7�nڂ���!�2[Ν=�W���8
2iY���źI�b%,k.���A1�pu1�NsJc,٣Ȧ�i��V~��U3����Y�dz�K	x;1���6H���ra�Ǩ�R� /\���@rK�6��":w�!� 1��Z��5�2����"/���M׵QwY�\�]mפm����v��'=�c�mj_�3'��N!$}Μ9�w���.p���*�k{�����7�r9�|_pI&sߗʬ����Z�ny�d�J�H�{�Όg������qΝ��z�c[[�e��k�U][֒�U������ 	 � ��׍" &H"���'�tm�~��5�#���l�0���.)-���/���rJ2���4 �
Ύ�	w      ����1���5��V��M�:h��U�1w��Y��1�{�.�����s�[�1H/K��fk+2�<   �	�x��O�ss��{�Ԓ��h��*m>A :677icc��\����냜#���[}m]w���ۨ��ܡ�C�1�sQc����@������U�Q���l	�v�>f�>�A)պ������KmW�ڵ]��*;�ѹ���&��� ]����+*�v[K��;��j;K�>��S�Z��CL  �ش[Ϟn���4�W&յ�G�(�^���l�.]�L����1w�ܑ�G��FpA+G�C�������fpS��˥�Nfi�N      ��||�pm7�*c,�����Gq���+�'(�$�8���m��_�@ �|��w���v   ��՗_ҟ����/��������G�Gݼy�._�I�0�w����Cr�j��q#���ꬹk�ża����X@�0��Y�T�T,[�R;���g8�B�H��I��=(nܸA Z�f�i�����ۅ�B�p�!����vm']R�g8��k�u�<)�y)��y�qm�{um��W�;�$kV���H���   ��y���&p�,�n��X�k����۱}J]��=f�Yz���t�k��G	�n�M�Ȧg$#�,�)/ Q\��@��O/�d��'�2���      ����,��J4:Zt$�U}��M����e��Z�k�E�9�۷o��\>GK�+����2m�x��%   �c�m����"���&�NV��Z��FFAQ���_���<�y@�(��4�9����{۴��:��쏢������tR����si�y��GX�.Z�"f��w�Q�JA����7�|C Z.u�"	Ƶ]":���ڮS��=��i�]��:yI[����yj\�9�]j�ݶo�?�+P��L���   ��{��1�./���������P(������U�wo�����>��=b޽{G�=�k׮%F�V�L��*��W^|"�ZP�����2?R#      �p��\��(��ɸ�5r�FR�0���24�A��$c��^�ӗ_~I ZV��Q6�%�^>��1����/   ��믿�?��O�ۿ$�N�1���
m��$�?���t}�s��:1_��yV�vŜ�)v��3y��7���W�tc�C�f~�JՌ<P�tbp�0xsb0�ZeE�>+6-D�ѳva݇k�f^�6�v���*yK/�!���]��W���A�]�ڮwD�_�N����&    hX�����v�U���	�}?J���z���{<�k�ȅK)�˵�A4��ͭ[�Z���*��~�ٮ���pI�J�+�7� �����B���W�       ��b�F��1�,�����U��|��ܡ>@�A7>|Ho߾%-k�H/���i��S��  �����--/-ӛ�o�����!p������ܤ��{�Ǐ[��uC���=����}za�L;�g[Z���56p��H�jB�Ze�}qI���*I�J��GPJ�ݻw�Y�����.�;�����E��e�Q2\�e��"u��c?y���:ϐ\���s�����@Ф0Z���	�J%   ���~{�-�����~�LRO%BA���p�U~(�FFF�ҕ���ۇ��M����׎�8�I�c��Z*!X%�J!&(�A�����j� p     `8m���HfK��Rc,�C�z��Y�ۇ	��d�[���]������������-   As��M��_�������3Y_������7n���z�s}��ݍ~ukQ*'���w� v��]�f~.j����@�0�#����R�2�/r�p�NE��̆��B��F�i���ٵ�YF���\�me�g=;�S��pm���2�M�m�=���F��?�F���N   @X�������;ؗ�O�k;��cG>q�ޗ�ݷk��Vytm���!p��/��"�v��U��_��{�s�i�fF3��       �p���f}V.ҙ��ܡڵ���\�3L��U���D�����a���.ғ��   vϷ����VVi����Q���y��~G :�ܹC?����>�9B�u6%��KiPM.}|!_��)
����qs��@� sc:+��h��ف!�u��]�.e?��>�A)q]�Z�o���@�8���]\�5aC�p�������*�����$�#���|�rm7�U�ݵ���k� ʷ�ۤvm7ʊ�︣�C*��   ������\�cgo�,É�O��wmo��X7Z�v��W�#-�_���O��{�E��G��`�)���U2�H�@����$���{��rw      ����zB�¨ÙM9Vҷ�'o��k�Н=���	D��:�����KW����   �oݦ����{�a.��G�W_}e{�=�u�:�*a}k]w���-������?g�e�h�R>;G�:f,`@� Wg��9�8�nIm� �07��'�qu�Ş�$`Ÿ{�.��l6KK++�
a�Ñ�t����\��V��n�������by]&�'��ڮ�+]۹6���ѹ����k�y>
Q����ý  @$0���_3�tm�P��ޠ���u���iii�޾}K ����͛t�ʕH�I����x��,Xe����Un�*����^/!n     `�x>Kک&up�������=��:.yC~�0���A/_�$-��k���WޣG�%    l^>{N�����&������5���M�������n�k�>W���i�
v�/	�y>7���b��N������*�e�X�Fə�vso�.NE��!z�P�0xN��$v����s$�ϭ��T���2޵ݢ}�J���µ](s��5ތ���9���e}��;�Ѝ6��ٗk��}��]!�'�����n�`���U*   ��i��<5?G�GF�v����x��k�X��G� p��H��wPo+�]��N��_�q�nY �E��pp/��
      ��u�7�Upp���(� ��"�ża��C�0IW��c��7����)���$�N.�������   6L����'�����Y�ӓ�P���o��������煵�!
��~6׷�b���g�����l}�A�1aA�dT?��$Q-
�m�3� T�d�QO�r����u���'-�/�/��\�;bj��;�vN�m�͵]s��ޮ \��gb�Z}~�^]ۭ���O����   D�7_C�����]���%X�k�����{٣���W�_��	Dǭ[�(�z$�>v���Ry]d+1f�(�      �tF%n�qޙ���[����Y�Bخ@���u�~'�Y=�N ��.����  D���-��ӻ��ce�=y�@4�>3�bwٺ�ԃ�a�!t7���n�<��<�`�=�eƳY�J�t$�f�pJ�R�Y�r�n���V���۷	D��yn�A_���69�����K��5-b�v�y���.�]��&n玧rm7^��ۚu]    D�m�~C���+�P�pm��\��W�x�v��s�T���)�h`B���=���k����P���s�5��K��:	�UN��`389:�b~�J�      ��r$��w5����pM��T���FEzn'���s���^�{;  �H�q���c��_�+�����{԰��gnQP?}k�i���.�k���xs�
��`� �11��ӓc*FM�����S��r���wb�+j���y��-={��@tL�����D[�ΐ���l[�]�ퟑN�(]��N�s��vᵣ��;�g�n��F���W蛯�&    j~����O���>n+��*vI\�{�M�������X����W�֍���M7x�����X���un�8.K!X%۷l`����F��,k>gw���e���     FrDǇGT(ly@/b�L��rڵ��'�u=�upp�����/.H�SS����V   @�`�X��3��#�����f��\���7oR�T���g���i~嶎=o���2M�}lo�ϼ�d����!e�i��^��xo.KT��=N-(���e|��QGZ�	}�V̽?ZѲva�ŵ].��<#�3Q�-sm�
�%��g��zv%�Y�k��L�^(�.o=������vvsm��>96Ao޼!    j*�
��:y��E���6�*��v�{����@�!�o���Ö�}���y��b�ʪ�ra0�WR���%n���x�0?      ���y�3�&�e}ǒQ�=�tI��7�8�l�6�#��X^]i]� }��w?���&    j������1�귿!�.X�xay�޼�"����Ağ~�ib�a�i.�w������7�H���x��7�ժ�>��g{5J;���X�2�tDE7�v?Ir��~�,1�������V��ѣG�eem͗��.��	މ����J�tm��9�w����@�z+]ۅ���ڮ��a�����.�ӟk�f+�����[�tne��}��   ���կ~E�ӟ��W/�|ֽօk��vY�J��W��%�r��}iy�
a�k�3�|�{\���qc(f��=g	      0���5(Sq�ޔ�����_��;��<�@�0z��&H###T=�P�Z%    j؀ƑL��Uk�v�	�{t�>߃Z���h�Xe�v��\��]�k<�a�ͱZK�.N=ۣ��{@Ld*t&qa�%��1�~8$+Is]�e���w��&�XZ^�ܿ�?
�t�Y�k���BpI� \��7W`�uum'�c�ǵ���� ^�v�h��v���)v7��|X[^����s   �����z�)BUjأqm�R�&�v�drj�5����;�p�֭�4��	��z8p���-�l��A+bv٣����t��      |&�:�2Μ!g�e�7��)�~��.�c�^��"���U�T�Ax@��N~��ߡ����   �����/���|����5�t���J����=J(Q��?2�����_��g|�b���23�<�"[?��
����H%���
�8V�Z���0>>N��F���bb�������'&'���'����J��tG%�{�C��s:����U\��muy[�˩T*�
w����r@��c��
��޿}۶�׶��)_q鈴�fѻ�o���[.�9-�كG����ȓ���b�����666b96��b.l�8`�ξ?�r�988��/��f� �s����z���%�<w�Y;>>n}�����,Bq��0������WZ];GG'���k�}描�iow������n�����׿QU��Wi�����?��g�������I�c��7[��ޱl���y:;-)����>	�W�k�؀��ϟ��˗)i�j�i���d�'���O_���)�n��     �a [/9��]��r�^ך9C����X$�u�Dސ=�m˿����������*d�   ,9;5Cc,0�L��Pq�H%��!f�œ��q�W������wM�y�.�XBܠ�3�S����Ѳ�MuQ��xa�]��p\�$O��q
�ezA&nBp�\�%�k��㡗s��;��kJt�V/w���V��ާ>�f�S��˅��3݋�{�N�޶��KK�!� ��`~�\\��2����ߺM׿�qOm'�L�vѵ�lS�՝�7��O?q�ǥ��ɧ���?�ҥK��_����Y*���}��i���+L���K캋&P�p���������~�صq�{����ަ������K�����y����c9>�?ZXX�mpA����~�3z��R�noo�^o��k]�
CpmW����~M���O?��������G]��i�W�v&l�V*�~�|׺�{��i���}{��wR�$�I�^�u�Ν�g9)
a˸X�|�K�"v�"���׬83����      ���5�����`�s�B�6!��H�~��I���/_����݁4�byC�������Y�}��㾎ͮՃݽ�qB��������&���~{�^��%�Jg��[YZ�������cai6bF-����ۋ��)7gb�`�{7�<w�=�οR��r|f�=��L�0����!�g���o��Fǋ���#]_f�`���	g���;ψ�>�trJ#{�{�p�og��}�}��8������O�Ȼ����X_������ܢ���JX�[��i�`s�7$י�������ww�`���~�����$�[��Ī�lSߑI
t�u���#-���)��v��&�G-q��K���n����le�<�.�_gs�vv�8'ׅ�:�t��T}������u+����O�5�+��A�N����v�$/�s�0BǇG�   ������u�۷�*��Wq{�"�~�*E�rex_u�ܫ+{��Q0/����Y`X�D÷�~�P"2h���d�2����.V���7�%x��_�����     d&F2tvvJ�¨ҽ��b�7��V%һ%=T	�8�l�v����%<3�&q����'�&1;����O��{�)�l��əi�˨��c���{��\:���ZY_�ݿ�����������l�̙�w���t,�O�{���[���h4�A��L̜��|����&����6�{��=��e�(�~o�ʰ����~�/�$]���ۺg&Jq��|���~������D8�X�����k����Y�gtt��IX�����7oҏ���ԃF���tx.��_�_��N�(���Z�ӆ����,ig�R�pbp��_�H7q|p������K�?�o�[aB���y���S�����z|G���ќ\�����\ŵ��;��~��׵����l�̶K���������+   ���{�飏�c
�u��]R�k{�����O��݇`ݯk;O~$Ok����]F������_�����+c`hkQ��O����sA�\Ly�
     �!��l���j�;���`$���E�~���$�(o���>|H :ص���L ]\X[��O7   H
L伲�L�߾!��ϭ���{��QK����:��|?�S(7�r���>�[�0c�
�FC��39z�[�4�{ ,�5/����&f'م�t��	����v'ɑ�<x@ :V��Z�uQ4�ݵ�+ٵ�*K�k;;�����ǵ��.��C|O���v�l����	   H
�w��`���lkZGgYQ�\�Uu�ڮ��ӕ�߃�=B���9�
�� B
�q�;��K+X�}��՟��� ��]��ևP      ���8Q�"IP�^�}M����n%)��Z�@m����<�;�� =\����?��   ��p��]�џ��)c�Xl9�����N3IWA�=���m����1@��K<7I�x�R��0��RY��V&�� �p!���F�I}A���?B����g]�\��=b�W��7K�lI�V�ڶ�%�Bpm�I�F.1D���;��Ѻ]D�>��@�o��smw�ݕ�S�ŅEz��	   I㷟��~��?��/�BkĚ����zw�v���k����k�6��ɓ't���X�M`�.�.x������28��\�����Ϛ��       ��2��PYq��g��D�����[�H� ��	·�~K :�ޞ:
#*��7{  �t�~��F��Uk�v9N�~��`���Z6�m�N���������};�ny���"���s�|�l�Ni� ��N�#)$�v��])d�vl�[�j����8������trrB :�W�h�Kx̮���	bpI��W��ծ�z]ۮq��}����v�\Ϗ�~���/��   ��qxxh��k{�mRW���G����γ���
�����G��0���k�"�{[4�0n�>ޏ��[_����      6�z��.�X�����FWlyC�[�3�<�<{��vvvD����t��w>��7n   �4n~s�>����~���}t�Q���+z��5������仺�v�A�.�Zy?�_�_�=.3�*P���= �g�����<\�F��{8J�`�8�c�A&�����)���ܜ]��~D�my�].��zе]V�һ;����.�D)��e�trt��  ���f�_^���ǺH]���'\ۻ�����rt��:��xF X�KF\�a��bǥ�!`%�M���1 	T�J%�-fh��       �`R-[����ۭ���!u��G�7t#���G�D��-.H�ctttD   @���ۣߙ�&�.0�2RX���Çt�ܹ�ЃA<.{.�{�}n���=oH�~~/9�F�� p}1Y�P�D�¨�sV��y��6�뼻�>ѮX�"��
~����A :Vέ��iF��R��,P��N;,wQ��vm�� �k��
ܵ��&��^x����+��W�}N   @R�}�����M�K������z���um燐W�vq�/]��=Bz$�]�?�н�W���u��ޏ7�I�������Y�     P&FX��7s�lI�]s�N����`�����SD�0Zf��(��H�VWi��   �ʻ�oiq~��w�H�B��f��p��@4����&�ܢ����j��7���F<���r�y��8m�{�\���r�(!9-wR�3�C�ca�1_G0�%)�~���cyu���S୓�ƞl�vN
�ѵ��_O��ƶѹ��$>�4� ���x�
����'    ��{ȓ�c�f�T��S�ڮ��k;+����.k�������ݻ�h4Z�3F�"t���e����b]Y�ݳ�]�b��X��T      8g2De�֌���<�=oh�5��$�y���pp��e��kWާ��/   H*�oݦ��G�����})�����ci���_u۷���~�V|Q=@]�74���z��w�昵��L����(�@��'�E�2g��v���.X�*X%�u��v'9����9+t;.��	��ݻG :�W�5�F�\�ۓP�k��пk�D��E��j�Y�h�M��l�_�v���ֱ����E��    ������O~����զ�<M��A�߫�=.�v�peu���g�k>;;;���I.\�k?�����[�N�ʵo�$-��/V	q�n4Si�3K      ��ce�(S�8���.$�ct�
K�,¼ar��9��cai�@z`n��r9��;   ��7�4c,������A�k���
^�.�{;�{�*�L&#5��d4Z� z�K��>��T�"��������*��#2%����W^�xA��)��FL.��مYA�ݫk�U.�׵�o[��X i{�v*]ۉ���v��wm7�.�[�����A   @���ۣ������ۄk���ǣ��������iu�m�xI |�ߍ͞u�����н�M�ݶU��ߺ؏Q#���מ�,��=�(7�5F      ��c*[��b@�J�Nʁ�Z��!��G��k{_�~�Z@4�����ӏ>��7n   �tn5�>��ݺw�@:�}i�lll���>���v�;�W���uD��(u���r}xO�wS�������3 p�|�LUc$���5�\�|��;N��8�$�.�Ӧ`�x�,�,S6c�j�rmw:����g쇀<:���.i�]��k�M��9�n�;��rm'��]�vM5�|�u���c�Ѭ��\Q  /�=�əI:<:�L��R[���z~�&յ�������\�t�y��i(�MJ��ؕ�R5{�]��|^pue�/��)A�     �`�m�)���Ͱ��9��P���t�vٺ���#o!ӳ3-Go��'�����   ���f�����.��P+�����Z��2���?��XD�n�[��c��˻�;�󆤈���eTg3?�PZ���OՒ}zq�E�-P�p�a߾{8*�	�?N :VVW�c�M�]ۉT"x�_�f:�;���.m�\��ݵ�lm��K�v�#��dmĵ]����6���:��_�[7n   0(ܼy����˖��Q��֕{�]a��˵�����[�[[#�=��'E��q�q)#`��������������ͥtrBYm��z�@      @4*%3O�O+޵O��d}�ֳ.yCUB�%��W�� ��d����Ez��   {;;4=5M�������G3�b�^��"{.�j�E�ۋ}z����z�+��~F���9+��ܭ�M3h\��Hp;.lV%?�Z�낌�����E��ڮ~�t-b�vG[a{H��r��؆(\�ݏe������m   6R�Z�t��k�TD�"�v��vym��v~�������ȎW�ʀױ���µ(���7���q�%.� yv��S9zyP'      �`qvzB�\�S�Ж7�&�53?��uI��7L�@y�hYX\$��]��~��&   `P�}�6��������������x�@4<y"��"P�|�P�R�W���k�@6`�R:i�a��
�}�8��Z�J�Q��*Ub[��e!��[$!������-�bj��D���QF�z�M��Y*Z���{pm��%�]�]�n����9�˵]R��&����G������  O����"���I�õ]Z�����˵��M585=E����ٳgtxxH��ӭ׃���q���f�4e}�â]��݉�-���     0Zy�Z����G�vU�[���@uސl���&!o�P�<�ava�@z�6�H�u�'   �J�
�<��0��@ :�`���"C���l�?+���\�^��۫��,�X*�hb$CǕ�����d�����R�0��2:"�.�p���u���Ar]�� �gfh�P��ӵ�#��T��=��i�߮�܏k�ޏk������pm���{-m�b�3��-sls��y�s�6   �ƽ���?~�!m<۰�G���,�O�]���jT��Ы��v����t�&�[���3�������	��lɷ7��;/5s����jv
���zݝ2�e���       ���T�޾d�����������$�����ڦ��c��� ��Q�'������-   ���=������]����4�G�T�T	��Ç�I:z�$
ԃ6�jI���˩���5s��$[a���hm:C�ә;�������T2��u���]b�cX�)�gA�j?HQ���Lm15	�i"C���:��pkm�Yd���(k�`�����W�����g�͵����\�e?{��G�i{{�   �A��՚i�0��pm�ϵ]��z�����˖�]�p��ۅ�f��gQ6���B*T�eX�7C      ��a���k�9��'�ż�8x�y�a��&�7,���a~�i����_��   w�ܡ?����	f�I�4;?Oo�^6��W�����}�g�r�����������zM��*N�q�2�4F��	�}0��SU�𸋋�T�t������#`�6>D͠9�3��".��4����ݵ]�Փ��w�	e��U�����f\!���m�S .�Ώk�c_Q��P{Y��]�$�A�|�N��   T?~BS�S�z�u߂u�u�9���ۧ��c�umW�Ӈ��Gq���*����܌��Q��)�\X��b���su:Z�K��E      �\��}�gQ�������C�P�7�Ǡ�ٺ/^ o!s��҃��l1c   `�`���,$�ibn��0�/]�40�ޏk7�2��BT�o����>�y��\z���m�#T����5P%�P�\�m���"�@,Kb����D��Ғ��[��nWP��|n�K�ڮs۵7�����,>���\��O�ц~]�e�v�����t�"���   ��������O<�ǵ�O��]��{�7"<�v���>���K��f�d���O�J��]��x����_��/��Te2��^)�      #�2�$��]�>�<�yC��}��q�N3s������s��%>_   ��w�hzj�a��
0�P���KNnQ�S''���I5��ݖ;���k��_
��9�R�t�uPT����`�i���%�ݮ�pe���3<H�l��l.G3�ӝWy����������ؕ�f=��Ei��Vc���)����k��NB�*v��� �:�NSܮ�������drtu�e��f�+����   �J�ѠZ�ҵ^8��5�µ=�=�W]ZY�-$�#�ɓ'�׃��}{��]Ӭ��B=Мwb 3P%� �.g����Y��       H<z��I��o�ж�|��yP��ٳg��]s������G���?   0�ܻ{�Ο;Gw�}@`�a� :�LZ2�#P�︖�O��X���m�~��]>P��.[;k�e���}P*7/$�*2.T�]��}v�@)�Q�6KZ��WDa�ťE�d�d(�"o�;��������!��J�v�#ng�I����v�\�.��mm��i����k�}��Nz��3v*w���I���#tt�Q�   ��_����r}8������ܫ+{��k�������k�G��ũ���u����2T�:�A��]�H� d{6;��D�^a�      6P��U"�9C�AL�LS~$O %4���   0�T�U�e!�L��Q�����cᣚ��W��[�4Iʚ�+���)� x7����R9;!܁/f�Y��+T,���[�@V��^7�sJ�#���	�#d~a��$0�v��,�ε�cۉ�#k;�//��f�mD�fەu�cyqm�vJ���x�\�H_}�9   �Kj����r��+w�nR\�E��	D�`�'�|K)L�v�:1.Վ5��!�Px!�!T1�+|}���d��dw      ��b�*�*�9�#:���i��
�ffn�@:8���2   ���=����:�w�
��m�hx��!�j5���`�(P���jQ�7S,��-. ۟�C,�JT�iT�����Y�ʐv�=0e<��0
C6bC�����0	�^a�v&� �0�0'\_N9Q���Q �	�Cqm��k;/.w�������~;E�����   0�{�Z��(󺭼\Z걞�nH���� ����b3��x��yK�"����1�gF�����oT��,b@,����     ���>�E��Ǿ�8.�m�\.���y����K�闿�G   ��Ϟ�'��)mla6�4037K/6����C��ڢ.���A�-�D�$�[u�}{��\�E�.�X���n���=2W�)S񗜶9�u�#��1/R늷���oP(��,P�񁝹���3��g�v�5qs�L�-���xsm'y�I��h�F1��s;��ڮُ���d2tV:%   `X��ݥ+^��f��+pm�����%n�Qp???O�l��u8\G��f8�d97؅�f_��������pE�C��H�       ���(�f���#o��q�@l���	�@:�kj40�  ���~ϲZ�@:��jt���Y����!Pb߬���4��A隽o���d2�L=ޥ��{�L�4;u�G�g���Q�ū�h8V�� ��#��ׯ	D=O�L�J�ݛk���[7kr"m�����zDζk��л�m����7A�v���u��A�_�?���
=z��   �a�իW��s��C�����[�
���˫�>������}��@���a�+D���L��bԕ��{�X�ZG�"��:��l�       �g"_��Ϝ!����˗�czf���3?7G��m   0,���hrb����7�GK?�X��[��c�}p�/���u��@w2��~̱24�O� T�{�@U�h������ �vq�#5��L�;6p��
F��o6��6�`&��z�2�s�3��,�L� ����ڮn�L��ŵ�!n��.���bqm����߾�7   ��Z�Fz���jx����um�S7�v�zn���������{D-H�s�$����|��׉{.]2����+�;      ������n}�v!�}웙�h�����H���������g�   0,<�ؠ��O�_n
��4Z,�Y�D |T:�$��z۷ l�N�]��K��{��O��N�7��V'�p�?�@��#9�JU��$�@[�����~����i��aN+�����K��Ե]!�����Z��&'�õ��v��v�ޝoCԮ���=Q����Q�Z��   ���c�f�T���ٵ]�PO��@\�����[,���-�A |666�ڼwi��]���R����vW��U������~�/0��V=k�N       �d����GbyC op�L����e   ��R�D�㈳����Y�z	�{�2�8.�{/������~"��u��]�.�sČ�
�6 p��vfKB��u��dImQȫ�0�D��}��������?N ��;�:Rn�k�W�s�ۮ�s/�k�ŵ�&��ӵ�s��bq�2�v"i�bwj��]������ŵ]<�񾍏��λ   ��{w��ǿ�)m�~m+ϵ]R
�vO�Tu��KK��������imm����s��$,�H�Vq��`�����rvz�|��f�      $�z��U��=oh�)�7�o6�ߋ/D������T+   ��ѠL&C��#nff��3=E�q�y�$�_�z\�X��5�����(h7�|���Yy�D��x�rVrMD3D76���l�N<�2!`�g�F]���-1��v�*`�vC�M�2޵�] ޏk�&�N�v��P~��]۹#+�Wtm�&n�ʺ����[�_�˿   0l�)��h����~]��ԍڵ�K=U]u[=��#���-�3A0w�s��%^�ľm"waq��U��X�ʥ���h_X�}����S�     H:,o�D3*�5����߼yC ����^�B�>"   `�x�t�ί�ӳ0Vvf0032؀㓓����Z7I��^���%�vu��9K�)tw���K��f~����{����T�tq���m\r^�<bB��gs���g_�̍D���\(��ium7��RGP�+�k�̧k�Cl���L�f   F*g�t�um�ֶ�\�=�S���v�C=U�z0R(����ku����n�0���7+s\���<���o܌��z� >C+�     �t�G4�T*T,�[�7v�,o��ؙ���=�..Ӄ�w   6�={F?�� pO�s3��Z�ҫW��>��_/�64�|ܾ����f=���%�����N)��TO�������d���P]`D$<�A*�%�y��2IN����ׄ0�̈́A����&�㻝���8e�j�"!���7�v���7�"uQ��pm�0���ŵ�^o��j��m_���|t��S��"u[�I��aS��5�p���"��õ��@V���4O����~D'k�ݛǋ���{��繳ABq}���޳c�}�����ٱ�����7��\�� ���8���Ϩ01FG��B�d[*�E}����תUr#�v�_s�۷k����F�}��Jɵ]dna�޽y�}�2�nWX�x�sn�"͊^�ZdbT�D)�h�[��x>;
�      I�L���{��yC!�����}�~��@4
-�H4  `Ha��ls8 x�'&(��6
X�mss�%pw����_��҄��κ�Z���-oHB<������4����t���Kc�N��g��"�E<��'��������靤����[�A���ߧW��,���&�q;���)�x��V&
��m�ʚ�b޵�x���KOُ!ݝD�-)pEl��Q[�vx�O�9��q<�Q�|!�M�T��٥G�;���qzF�ǖH�0M�λzx�MNNѷ7����E�������v3y||�=L�W.�[#��������M��={�Y�5��
�<�����󑑑�oN�y��c�yq�γc��I��e�io߾�>��v�w�+}|�~J����1o߼�k�~���������޾�K0���.��P�^�}vo�g����U�0R��ޞ��U�.��}xTΎ��'����bF?߶�>�.��[&�po      �����'ޝ��{�yCqP,�ۭ�c���E���J\1T�s�������Ўͮ���i��p����;0f�����Yl�^�T�����O�OЍ������Ȏ��QO��,�:�qǔ%��]��}��g�+���B�y�,R*�b;�ql����8�{v���q�ާ�3��޹}�ʧ���#*���g���]L�g�,�7����ǚ���z�;/�{{C�������e�2x�E�9��p�����{i+�Ms,� yQ�̖���;Ӆi�.��´��N��ET�*��
�`#~NOO)H�{�>��~0��k�7N<n�~僫�އ��]������j�k�y����������ݵ�VOӅO��l������7��+�폓ҵ�ٮ^]��:�&����9��e?���w����d��O>��^�����������`�*���-��8`�����c96�������R,�g����u���{�:���gc�B5�s����3366F���?�sg�Y�4�����-,,�(��g�VL�o|�����������D쾕����~�S��]۝��r���;��t|՞�U��o��X��_[_�p�n��W/��������3��[�t��4�~�kj�^P��5aiו��+�kj�I�3u��      �b���c��x]��&R���8o��_AC��@�"��{lb��Lx�R�2-P��p=����1;�i����_:�=�6R���!?~�����q��yO�{o�"�y�����q�Ń����W��t��z��atǏ�w>����x��&��p� �{k�1I��Pͬf�/�ܢ�ҳ�4iRѩ�������|�;_G�O�I�u6���D�Au��nIj#H�����N*����X���^����K�0;;�zE�2���f�Qfsm7�qmS�-�1���gB"�fu5�Q&k��Z���m��u"idBr��$�Y?r�:��M���&n����6�T�Vy3   I�%��N,<
��"x?������'"�z����ա���Odn~�@40�;�b�ȓdw�^�W���uDq�:X�P�{�ә�T<D      ��ԩ&����H�'����F$�y��ϟ>c*s2�kV�o����}va��C6�9���*�NK4>5Ic1��ۍ��˥��߽�:���ޣ�Ϟ���hd�g�LOOOS\�y|#n�����3'if ��� �sg��l悸���দ�bsp��g�t&r�g>z����׮���w�?������L�����D��X3�s�s����pp���n���E�9X�E�Π�_�؇mˆ�~��O1���_�s�rog@��y�R���X�$`e<e�"w�rIoQ���[T���LZ0�m_/^� 3�3�6��mN���B�Q�M �ߵݱ/�k���l(߆ \�u������k;9��Vh�����)��@�N�=    ��g�ra�vv����wmW�k���Q�����������{�U vvvZ����Ůu��+E�
GgN��)��Ur���(����A�     @�ayC�K��Wn�ٶ��^��8 ֶV� (&cāh`�-�L�   ?�z���3=3C �6,NZn�-%���mP;_�ꟛ��5C�u����R�� �tI��u��mT�#%��f	Te�vˉ���`]�n��Nr0�딅'''�)-@�L�~�;�o-@�v~?*�� Ж���rm7��6D�ڮ�ֱ�o��������'   ;t���t�>\ˣ��k{߂����Gh�Ph�@�4z��-,,�*0�mZI��c��y��S���.�Z�	�!&       �d�e���q��.T�۝yC�����2��г��B[�^   0����������^p�lf-6;�1�[�.�����w�+G����r�bސ�+����y�d�4�\�����2Ή�(�/ޮ(V!}nM�0e�۷o9m�02>1N��QS	޹Z�x�[_��ߵ��Cǵ]"ZW�Br�%&��m7?NѸ�������sg�ѵ�:?vv����,}��o   ;�����U�ݟ�]V?R�v����}
��
A�.��=ө�������AP�0�V�l]s����ɬmV�b���x����D��c=D
      �?j���^�\��'�|����v黤8o�^�j5��F��������W���   �a���'t��З��^�&�)���R����o�O�C�s���]b��=�\K�to��g��3?)M@����Y�Q�R%��N�=�2����R%!��7oބz`137�k;9�um�H�.�!:�v~ �p�����	�H�o_���{�	��k���&   ��Պ�u�]ەM0�v���1Ѱ��@} ��blJ&t��Z�{�ʸ�w��f��K�0�]�E�vO�'      �T�ʔ�f��Xƣ����;�ud3@�����O���D���/�@!7�r�   �6�Dq��p��Hl�&�?��ڢ���ĘW���/�$�vY���
�X��!�4~`>
��r����'���:x##���,H�)pqb\�T*n���IF����G ���;�'w���~]��u����~��{um'�ߢ�]-R�	�[?|����nP�P��]�   3o߼���q:>9	ŵ]I�޿�<�v���꺝�1��w�ޅ�_=���΍��ҊHkk�6|__��2��]Öٱ,�b�*      I���Z3�es9ǀU�Y��A�D|��ڷל��_� o�095E �h  @���^*)���n�XI�����m"w5�Fg�n�%�%�W�~�r�[f�Ŗ�1%@�Ѭyqے������X�2هA���`�;;;�����	�Crm��J���۵��J��N!��q^-�]�Y����+�H�]?��d��G����   i��Ç��?�1�H�µ�뱒��η`��`S�� U��S+�]�Rv����A�|�S��;1�g
�     �T�3ds]ScY�B�@�7�	�S�7k�5p295I`�-����   i�tF��Q*���9M��A$�9�s��r�gc;�L�k��8Ck��B����c���O�Ƴ�ո�3ɓ�ݝ:��qg��F|�(C�*:����t��Џk{�����n����$
�em̵�l�µ]*��m��������O	   HGGG��e�R��{��_]?݁ \�yFG���7o���f�T���:}s׬];���*��C���w"�;      Ief�y�^�;�1�I�N��3���ʺ8����Z�5o�T����F�����fq~��>yB   @Z`�{�_���%0�����=*T������Ͼ�9D��z���ܡ3o���"�͏e pj���j���]l*�6��V�2+JV��ۭ���{P�ޘ���
ăpm�]��P�յ��/��֕�v��i��������.��rm��'������4�R�D   @���+�+��{=�/�}߂u�u�ۏ�(��P����|\lmm�?IP��Jˮ�x��0Es��֮',/)�B�     @R�.4��+vc,�l�g���]���l�לagI0Ȋ#o���[�0��������O   @Z`��^��;�9#ܣ����`�-e��&M*�f~��yC�v6S,��,���j@��ɑ��̛��rY���27epJ���3X��=h p���q�Eꌨ\�u����T�n4�^f\ޢ�]���\����|��J�е��#�Q��  @�`.��|��ժc]�N�pm����{=���~���4����ׯ_������u�w����U"ws��H�&FL�z��`U;� �!��n�#Z��CU      I����IgA�.KP��^������ڍ1s��5q���;�~)���q8�?��    a��v��I�u&u���kn����|��*����iw����ĳč����mIl�A*պ������-�@>c��Ϗ�ir��rm�������2lr���vq_����gLW��]�p���n�K����N�յݠX��Y�F�  �.=|H}ﻴ�%@Csm��=���	˵]�:;7�{�����ŋcmG��y�S"?�]��q����(s}�iu��     �dR�4�ݱ�bsI�� ��;�<�ob�l��fz��$����o[�RA�0"F�E��!%f�߷V�   �6�:fr����y���?c��l6�z��U��Vi�5��7�����yC��\�n7��Z��4�^�O
Z���+tuq�'�5�zc���8��b���u���c���!>3�3���k��˵ݱ/_��6xi�b_��b{Tۅ��n�Y^\���}ZZZ"    M���4�}2ҟC�ڮ�
�l�nR\��z3�D�	D �L]�pa�T"Ҁ�!l������j����}68n]�%��      Hy�F�1���>��K�����.��+�����Ak�319I`�Y?�FO�?���Q   ���˗���J/67	/�0Ɗ �3<99�����u�,~w�[j���f~V�myCu��܂���V��� p�I��wS�ncOb��m�|e�m�R��~�{{�f����𙞙�<��~\�u�k;_��=7����Ե�YG(s��7��A4�}�]���Um�~�&�ƨT*   �6�=J�Vϵ]V�g]��{?W��lzz�@������n�:����$�+Y�S:�T�-��J��H      ��mԬ{x�'��O��i��yC��;�K_�[7J��!����	����<}s��   Rǋ/�~���9�S�G�u2����q��m�*rW���{���e��|�8���[�ȥG���3�L���w�ywpo?'�l2+I�4԰/��G��sb��q����� �m�k;2��3O��d���N⾽����	ǳ�K�-��V�'z�Q    LjoS��k{?�p�v]�g�aӏ[^�T"FL��C��enD���w+>``�͛�h��2      ��Vo���!���6��u�o���sW�O�,7��C0�:�����a&�e�y  �J��*�s�L;��(���w���ի�0������7�q�g+o(����F9�`q��|���L�9�yubhc�L5�B�j�7G��i_���m���#���a7��2�v���pm���\�M�w���2�z˵]�_IYK�b���"rm7D�e�j�   ��rvV�\6G����P�S��^(��Q���'n����31g������TB��:i�]��k�d�pbw.PU)�       �Ԫe�}�Ù]��n�l��=j�~�chk��i���7��h��'0�@�   ��gp���lTt��m~6-�µݹ�\+l���3?ט�==3?C��Z��z4�N.�v�4��Yg�����~?�I���@Ut�@�Z�.X�tm'��Q�v[|��K��:���n	Qt�v$�G�MR�z�v/m�(��R��   ��勗t��y�~�α��A�۽���\u�;>�{d�)�t�;@V�Kf��:�*Peݫk�x���ئSΦw/htRF�     ��Q��)#1�j?�r�\��&n�d��F��a�0Ɗ�����%�ɴ�   @Z��|f3^p?���_�����>le�6U�L�7Eiw��@s~�"n�<��Vr�O�*����񉎮H�S"�ٵ]D�"tm'��D$�۵]�˶�ͭ�"/��q{�6q��F���9���$    ��|������]A��k{�'��f��RE]YMi�Iq�H�\��5�Z6������V�n��[E�蕲/	TA*2��f]{�J6c{�0���2�m      �D.CT���PuTU��I�X�^��=g����-b�^���7�cp�f�����6   ie�y_9;3C�
C0����=2���"������� ��Frl���s��kYB�x4���"$R����ו�-�@UX�#P�v�@|8\۹�+�X�
޵��Nׄ2_��n�v��r�=�n�o~�   i�\.S&c����ڮn� ���+��ӵ]R455�
J�p�KM��6ʴ�RפS:gg��a�1�%,�p�1@��S`��#      H��l�Q�p6����mV*\ڇ���=Y&a����	��^�� ^έ��7���   ���js��]\��}����=*T���ͯ�B�*T�5g��ߙ�k�:��htRI�������Ӆ�=���`�9�ɦp��T%�m����86F�\�+q
����D�2�k;WOx���zw[���+�N�筝���nַ]���n�x�~\��c����k    R��ݏ�յ�_q� ���u�g�!p� 6�*��
~{~�h�D��b2��!l�����=p�\�x      ���"�p��y�}�tJq3�o����	Ⱥ6��v��ä�_�c�h-�R&�!0�������   ����+���'��|>O��<U+U႙���g~��ڟ�f~feS��T� p��T�y�4�y�t�:�)��T���QQ<r4�����!>����gN�z(��2q{d��rq�%V���+qmo�R&@?�����;�C}���u��   i���=���õ=q{���:Wsbj�@�looS�R���QFTZv�=q�8���8����o��o�:      ��D�y�^�f^����,��|���O�$��V*r����������#�    ݴĭ�v_[�����A��R�&{��Y��r����#�����c��Q�'��`�#A�]��
D��TVY��d���'�h�� �������=��KD�Ra;_dkC8���l������zsm'�����)\�%mj��1j   p�9{��tZ*�^�k��v�k;�����9::���cO��u`P�]�ޮ�8�,�z�`�,�0�m       Y������Q�ԃZ;6m�}�#�y��8��35}����̸`�H(�C�>�@�   �$
��0ּ�=܇�=l���R7��-��ʌ����KA���^�5�@�x��J@��u�A[�N��O��:ʰ���#�۷o	����d��h�qg������/�v�p}�]���"���   �v^�xA}�ݖ��_��JDޏ��o�vV��0���`�� |�����#� W������*:U�p���`�Hw      ��h��4�o����f�0�U��6� ��Y�)c��W������16>N`xay�ӓS   �N�Z�|.G�Z��pR�}m0}g�f~v�˶w��1 �-�`�5h��iw�欋̼H�ܕm��t�J������+ ��	É!��ο�z���+µ���ί'nwݦ�v���PG��nqqv���{�   ���:�86ޟ�9\��u��tmW�B)�o.�p�
э��pW�N�n��+��m�K�U�s.֐3�J      ��P�ڍ�x��^����/h�P'���+��!�� >�&��˹�U�z��   ���zk������M��f&�6����i*g~�*t��r]�|68Q�\�@�$ZS�{wpo��4��*[R��s��~��wmפ�r��y!���Nr'ٵݾ�ו����Nܱ'���ݻw   ��F��ZlD*"���o���������"������!P)]ܻٻ�����\p�Mܮpp�Q��      Y�5���;?PULL�5;�~K�P� ZM�7�q�����7b?�;�1�W���E��G   ����-��{߅�}�-��xa�m���Ѱ�w�g�Z�Ϯ�tup��XȦ�o��F2�K���GY��ic3�kk�H^�0������TED�8&��ڮqE6�v�흝��u܅��xum��-��k;�_�T�U    Q�w��k{���u#vm(���!*،[i��� n競�VĪ�`=��� f��@�     @��i������J�sי���FS$�%�H�	�888 5�l�!    M����(�{���(�Q��kI��9��I�X��ֿ���0�$17���=�?� ;�߁*S|��bN�U����T*�6b�6tC"v�����yumׅ��(�䡻��N'���tmw�����n߮3�E�7G��
b{r�Q*��|�4�u   @�z���\!y��KǊԉ�O�x\��6a
��`��^�=��+q���BA�.	�����      $��^wܿ��V���0�}�[ZPQ)�.R̯��
�Q(��	   ����h*��=:�`��:�b�(rW�����G��{�X�0Ki wd�nsTk?���@����TE�hK�����.��kB-R�	�ܵ����ڮ�_���   ��ĝ(�vy��tm��"*�v~E6����U��2ȁ*�y#&e���U��*���+b	�:n����      H�������A�>�~)5�B�0:�1b0�:    R�����8n��̳|�����f��-o��4��l}&E�s p�T1����c�M�#
�)`�v��]������]�S/��O�MH�y�;���(t�H���7I��]�5�u�9�   ��κؼ�)��;��ȣsm�'��n���"��T)����ciybL�j�s��vmK���&�Y�������      HZ�2���߭�b�Ј�;M�4IA܏t���ӏy�I
� ��F��>�@�   X�wq�����HKͦg�,nw��+o(�se|��=6X�0��t�ePp�ii	T����{40��\>'�����*n�^�Jq���.n���������}��!�wm7���l�Qr   @�x��]�z�N�$��pm�Y7^�vU���c���{�Q	K`/ƨ�AT���
w��=�`�����
�      $�F�b&�����;$�:�DY�Q�c��ݹ�7���h!��A�
*��	    m�ad&��FƑ�H.�k-�f��~�kq�g���l٬���5����{,�����sMC���^��"e���&�m��|>�������l6� ��b��>|Dַ� �v<S`)Ĺ}��v�wg�=xh+SȦ��o��f/h�tpЪw����M%��\��vک���C��3�m�tyc\\�e������Sz��M��9m�z������*�J��1�<�j�J�r9��f&@���q��� ��z�y�q���e��q�;���8�o��z+I����١��#�q����U��w��t��ݞ�W�%O0a���;�>õ�g��tg���q�k���ޛ�I��g�/�̳���>���[rK�|���w����iw�[�ǲ{,�#�j��ե�+���Ȍ�8�	F�@�#H�A>_);3 @F1"��}����,�fξ̺�C6���?��;��q�˹Ee��p8����7���_���!d<�"      @��N;?��Hu��zᬼ�3���W%Ņ��6�.�9����}�\֙۷>�Ã   ���#���G�׿A=a.�,�	�E��s�M��r��`]U;4���y�:oȷ�O�� p��lqc��tO������lR��	2�M0��+Q뛉M\��oa�7n�ѣ?�@)$+�=I���I)��W,l��Z<���ӧ	Gt��\�SOc���x�v?(�{�����,�'T�	�}���z����Ŷu���O?�E_�{������Y td0���۷�L�y��M��zN�g�~��'}����z���յ��	}ٽ�w=)ux��wg�|ϳq[D�~\��ڙ�����}��[6�p�������w~�w���p%�����OON��gOu���]W��>�}r|LO�>�4VwxW�����^��w���������>|�������M\�-�(�Y���s�A>eL�=E�p��x���q����!�j�!      �g:+���aX/��In9g��t6�ڥ�,�-6���ަ�p��`0c ��������ܟ������~rx��5����N΂ݮ]prtl���8:��� ����췫��-=��\��7c���#1e�_�И����kg�yv�̐�,���}W�L._{��3�&W��������>o߿O������q������a�����X�~������k���%ɇˇ�﫸+R�s���z�͎���%�������������9�2A����$vpWݘ��hɁ*�q2i7?�_�@[�Sf0���*X���us�?�����7�)Ru�//)���_L�B<�/�:m���H�õ����:e{f/��P�u/��긄�]!$_���r��m�;�Qt�{A�׈kG�K�/=�����ݻ���AD8Ha"'���� �\����U�L��^{W������\�&\����fT�=����>o\�ۇ}�
к|����H���q������g[�� ������L������h{G���3f7��y��������8H4����:�n�z��Hro]����.�i�y^�v�p�Fܾj�e���i����;�]���6]M���      @�_σ�\<L2�b~���9!d7�&ʪ��(&L*[�Jx��]��p�.=���V�~��7��ӏ�o_��ݛ{Q\�6Lxe����?�3����qGe�����ٳg�
�����̙��������Ύ��8]^;X�{��=z���/_�7,����}���ݻw��������l�����~�?����|���W��{�����1��o����}k}3����F�"e�y��d��]ܣ2}���q�_�/�^�+����)@���ٌ%��7�|S����nX��+8A�l�%q�Gf��B=^����~�X/\��~j�X�n���ɣ����~��Jr�K�Ƶ��P�N*�����}e������"   �'ؙiIyZm���
���3�V�r�pm��s���I�@g�E5�
���E�"w�=�y^��k.D/��      P������O�$s��NɹAZ:\�$t7�ra����\����Ϯ�a   �,��>�?�yC;,3_�onQDm�ū�9=�p��7 �'cw��m��h&,yߞ�db�Y�̎��*��-*U�����ȹ@*/ZH��tmO
Г�<��~FQ���Ke)���9������]��O�S^����F�ΘM�   d����x����YaѮ�i��ڞU�l�v�n�7Uv`w��
�]SN�L�?�i�A�n0���ۅ����vgM      4��`�<?1v�I��_��>g('���椬ݙ�yC;�;!�����}   �t��Xk:=7��7�u����[��u�U��0�=e�7d����kN52�k �!��)u;�L7~�E,�M:1��?
vbX�@���9��	@���.�M�;b�Q�k� $�����.���J��Q����e��     �o���U]۵*v��+������ʇ�ט����&Փd`�K�'��xu�8fO�x^<A��;pp     �:lt��x^��3�5�k/>�����DE��?ߟL&��:]�    �0�PS��Ev`�X�`|]�՗Co��7Ê��۹8���6o�S��Ѱ�@�G�[$�c��7eRԮz.�L	N� �b[�_\\(�n�oϵ�Br&�D
A�\پ�k��<Ȟk{$�����?�6�   @����;� 9*�v�k�%X/ŵ]����H�ڀ�3����e֭���g����v��EU�굪�       �K�෗H2�P�?V/xU�N������bwg,�srrB�|  �9�   I<���L�V`�ټ���Dus�zq�X��;�tbɰ'��{�+z��m�pR] �lrND��v"��H\�V��H�^d��	�///	�O�� ��I��um���]���Ūk���^)R/��]#�O�rm��-|�gT   2�g��ߠ�I�cP1���������um��E�[P&��`8�:�L+ͬ=�<17��uΎ^\!��P���=      Ua�s=J�qIgE�O���H=P��0w��H��vC�� �w    	�kM���6`F���6fչE3q{��n�z��>�ƹ�TS,.o����,W p7d�+�����I�%��X
TUiBw{���e���D�Zq�,l�D�NH.���ޑ���vŻE8G���z=�um��^��t�   ����)���s�;\��ߵ����5F�Q���mbr���R�*���)�G���     @e�D�U�<�y݋�s������3�VӘ ���!(��k���/�ì    ���z��n�1ެ)�>Ʒ6`:O��s}�'n�ŪDQ/�����yCw �n��n��	Qn-�V)+,<$�e��n�^#sGB��/O+�V��5BvI�>���ubm{�풐��wm[ԞS���b�D	q���f�O���     28?�~�W�k�����!nw�ڮ�[����E"�E8�7C ���"����>/�;��,J     �����bWpE̞C��x����ԨJ3([�Y벃X@\��lmmqQ    �紵�Ig���%�ځi=�1���nf�Us�U�-�z��Q��;G�!��\��7�8Yn���W���� �i;t��V�� ;͵�����'���'�*A|)��A=Q��[v$�]ң�u���5��	�u��^'�7tm�w/
�766���   @�- S�Q��ڮm���i3�C>�����m�)3�e��ֽ칽b�<��'��ږv��x��      @�t[�|	{ ��Lɼ�j��dy6i՗�Uiw�4 p��*�eg{�X   �������{M���ln����2�E]�д��a��X<F�7\����^��i.p/̉�<�T�[�V�+����\����RYȭwmOuW'o!���u��1���K��<��|��E�9Iu���K*���    l��^��/���Zy\�]����"Z�����x<��#��x I���"��%��bt!p     �2������S������ �����t!�+ۛ��pL    �h{o�@=�$r ,��䪸��$�T���H��z�"q����3���k/V?�&N)��e���U�`_� ��E�E���Y$��k;�k.�v�pޞk�X�ͯ��������+L  ��ٌ�er2���4'q��pm״��k͒���O��{�X!Y��E�	���q��      *���RZΐ�G���&S�u�]��d��%ǹ�;���Lc,    	�~���>�z��4D\��yk]s�&g�(D���ý�v3�Ș�����
O�
Ik� ��{���:mYQ�L%�����.<��vw��i��������ڞ&��w�T   �@�n�ڮy��9�!n׾�>u:]�e�%p_�����\��
��EnR��b�ߦ      �A��Gۂ�����k�������zTU��=�1lW<PO666
   u��j���ԓv�X[TA��2�-c��?�_����o?tz�T8�Z$x�խ��ڎ\s���!L���	�x�v����r������4��I�{��|)�v�r��/?�������e�vA_   @���]du�v��]ە��uqm����VSq;N]l�m���5�b)4��H3 �a4c�����g[��6�      T��������T�+}�b*nϢ
�U�B��
,�T��`%��e>   ��a�u;]��wk�aޖ�[̓3̚Wy�~�/���e܁��݆�����|ERz�w�V��/O,�0>�E�����]�)w�um���ʶ]۽�v�sZ��]�P�k{t��%�)   >'po�k���������"�^�@�4z�f�J���C$�)�W?�      @shyB�c����K����z�1�
�%+�p���:po�7�%    @u��dmas�V��4?ły[Z.��M�5=e� y���t�f�������)�X��� [ʧ91Į��{i�v�q�F�v�@�N����v�S7wm׋�m�e
���/����u���ή0�v�3   @�l6�^ݵݼ��uӺ�]ۍ�I�f���<�]�@� P���y~R���!�     @eh]�ϧ�'t;?{&s�7�C�    4��:�ƹ3�J'k�V��˕G09Ts��ɝ�cu�TCZ|rY�h���Q�د��.Uv�;[.��j��\���R#���+�����q��k��J��TG8�?!\OI�b/��׵=!�   ��l%q;\�+�ڮ?�N[I�`�y�Z���A8?@�0�+��Қ      �CN<��{��9A��Oe�#�����    @��\�sǘR�N��u�-Ff׺���_�V�924�?�Ғo�7KB�jt�z���\;���c��ڵ]U��k{F�+��/Z�����t�,���ڮoW>&�k{���3    �!}O�ھ����v3q{���Δ��qm���nl�hNr�Aq���K�{�'     P!�8��:�񥌄�v�d}�����`�e�N�Z�#�    h��d�ic�k��tJu'�+� ��(M�/ĩF�D���]x�d��E�J�g,� )`�f+M�!+P��z�^t����5b�Rn��*��+�W���/�s"�\�iQ0_�k;�<a�   ���k�ڮ��޵}!!��Rq�cVp���� ģr��k��{y�      �J8���a����~�7���>w    -�'�ƹv���ݕ�ܧ���7��e ��	X���w����j�Jsm�R\�%��R��j���T�k;Ie�Ӣ�w����    J��ܕ��S�6=CL��󺪚帶�z�E���u=�E�|0o�F��NiE�Ųi�      nH찔7�'��6�n��ua��3    @�x��`�g;4:ohl�%�I�F�����.6�s�^C��D[GJ<����5H�H�A(a���=�H]S��?���I�r������uumW֡�\���|�#   @�j���k{ �^cq{^�vS������|����y�V�K��-6ҭ��U�     P�Ni��ZVN�@f���ÝYoW      �y[:iW�Д���⑿|��3.�nv xv`�Y���]��e��(��M]ۓ���,�v/���sm׉�^x�b_�k{R�ηS�k{�>bT   @*�Ʉ:�6M[�5Ƶ]�ĺ���k�O�>��Eշ�>��f'�dm�     �
��3P3V1�B����f     P?`�e�ۊE4�V����Z��!ѭ�%�j���s��}��m��l^�k;�(-�۹���%%w(l�_µ�����>�ye;庶׎�   �e6��_%��!�^]����B��d�qx�\�yZm�l�T��^-�[�r��     P��s���OJ'���m��Z<X`m�C<     �c�a�{�r��"h�!p<e"�zcV]@�@���\�M��Q�%�v�NX�.��-3���   �c:����pm�q^���pmO�� �0o��JK�1�     �2���sO)c���1p      ,&_Vh�-���I�����E�B+͸�!p7f�L2�U��C�k�v�-:��ھ����	�b�L�v�ڎoE�B����*��2���c?�b���+�����Q[r!    x�[p���k�Yai���4oXQw5�v�Nvhb���;˰!���      T�<��RWc6�����    @�h�0#��m��l/�O�F��8�t>�X�t�h��]�c��\�.�U�k{|J
���?}��k]�=�A!��T�k{,n'",   ��0���祮盾�e���`Km+ PU,�;`|     @u�R�˴c���6S�.ͩ0��vī9�+    z�=Yk<���y�Er�Ư/���]��g�V�]�k�T��ڞ��k{xNĻ�S�Kqm�����pm�1�   ��f>��#Sq{u]��륹��XP�k;_	Y;`a2      ��x� �M0���)��2    |O�*���F�O����!p7��Ce���̵Ԛk�,Ҷ���I='*��]�vV�+޵=)�O;'    Ȱ	���1Wwm/���L�^�v����R����VN6@�*/�     P��(�>Vh�ٲ��Z-�M�   �`�Yg�X����H���Mi��P��b���^�k{R�mѵ]�/�'i���Zյ]QV�k;��   ����攛d�µ}q{����r\�źH�١�n�      ��G$�&JX�uma�3    ��xX�l���Ҕ�� p7��Cu����ϾX��V�n��NI�5'$W���"ɑ<�k{xNJ�}R .��+�'յ],Ksm_�it�j���<n	�v��    5��۟LVvm�S��庶���w      @S�@?(�?� �����F��G   ��k��v���.M��A�n��1��}�@�n���ݡE��=N���k{�%=͵=)�����	ι:B_�t�'�NQ��r����.~�,��>_}�8   ��m�<�%��k�ھB�"\�5��>�"��g>U6���X2ߓ�     P0>�
柖@
��9a��    =��,��m���M wc��!$�*>/��v����[z�>X������y��>�L�g?���I-����5(R�ˇzRm���{�O��O?=�w��,J�K.8?;~�y�J(O��g��� ]כWo���cv[�z�L��.���c�bg��?.<}rr�(��`0���sg���驳k�����Ņ��ٵO�Sg�.����ap��\���]���w�}�~\�����}�M&'����{�._{�Y7��>oٿ�p|Eak�<��d���7�����r͕��s���o���n��n����k�����zZ�Z����ѿ��E��NNi{{�l������}^U��2)lJoؐX��*      ��vI�ņ�V`�&W���*;���wO_[���f`�ߘ��8�w'z���b�;��*�\����.�	�]���!� ���3����.m�m��!e}�5u�b��B�\L���.`_&����t�x�[;������k�S���#��k��~���;�ߨ��r����K\��/����E�U�um��?|N�'̟�b逮��}����}��	����+Ta��gϞ�޼yC�nݢ~���o���ٵ3�%�޻w�I�/^���O��+\�w����{��{.py����mmmY��v����۷���'��~���ܹ�lq��מ��������������Q��U�k;����~F��\�Y���wS����~�&�	=x�P8'�V����?��E��g����Ee����`n|��A�     ��0�rɘK�Źʎ3�\��n���C��l<�_��j���prt��%np>�������k��}����q` 2?.`F),�
f���5wi���w�?�ײ�+C6�A,�r�WWWN�g�;뻉�L���\��l��L��=wtt�Y��+�~��B�gc��_~M�p�����NzG�q6��ݟά��=�Ɩ^M�=�p����$�?9�Cl�fC򆸫�ܝ�d::M�R�Tܦ�+<�o@��7���䲰]/$_Ԏ=�>��ۓ�m�2~�\�u(QG8'��Rl??���^)$׉֥2_ѷ����e\;-\�)�^���	ۅ��#   @K��"6+L�nV�L����fuu��!n״iz^�^�vq���-(�C�ơ��K��f��      Tѥ'��;C��ĥ1V(4q%:�}��}��O�����o���޾|\��+��/�������S��_�u����������&v�裏��s�U�̜�����������w����>���M.pm�Ča=z���/_�7�.۸|��w,[\p��]'�7ِ-���_������������3c�*����[�f��;��X����湵�>˝mll�8v5?��9�HB�n�J+|�B����S�����^3um7�k\�=R	瓎��]�9��\'l���B�%��'������r���:    H��ti<��]]���*X7����Nʺ�\�՗5/�A%`WɈ��X��0P��0�     �:,3>��0]]
�m�     ��Hl�U�mkm�U���6���5�	��7�p3�Q��(�P)����lʜ-�tmWG��k�(�(ߵ]<�pݒk�J�_�k{�1    ��Zfߓ�\����uum'��*˵�o����n�u���?V��xF�#� ��=      �A;3Α�NoI����V�-b��f���Y     ����Z�{�'�b���!z�����ԃ<;�/pY���k�(ZW���K��S�Ϊ���1wm�w�+���'������4�   � �{����f�;��\ۥ�q0ٲ�m�ķ�/�J������       G�q\C���������   �L���09�D
0�>�#T���		��e�q~Z-����7R�l�0�*;��W���wm���C�rٍ0�I~i�vE^Y��+]�5.��)��
��
���9)�Ay    (��E�smW>������0\Wעk���ނk;_w2(��*gcނ���Z���      �Qχ����G�ik[A��0�aG�Z��!    ��q�=o3��/gl������k�,g��Sz|K'�?Y�B�k��xBŹ�3�O��.	�=OZ@dٵ]hWю�k��^�k;	�H|���Ν7�G   �������3���ZŻ�ӏ����ڮ(]O�q.(���������ߓ�Bz��     ����}2�:$���`�,�;�0�N	Ԙ&�   �e�x��L1εB��������7v����=��C�n�LvL�U�N���:eͳ���@��%P>㫫x�fŵ}Ѩ�	[��Ȯ�|��]�e�k{� >Y�_.��k{Z���Z�y    Ĵ��I��++j���}�z��tuM��Tw2�������z��{�틇p�^��Gm�k��     P3���9���s��C�R��"����?5a    4���\T]�^Dnr�i�<���9uÜa�c������!�@���UR&7xx��Y�ދ� p�T�>۟�e&$_ŵ=<�+[Ƶ�?Gc�v��X�k�HP��vR|�*�a�V�   Z<o�=��k��0���"\�M��Uwm���ʧ��0'{�/�3$����     �����)Ɣc)51X��!yC;La      j�t�q�ʞ�U�<+3�g�?�:������	���{���ү��Upi�P��Ɍ:�Va����K~�z��3]�I�Zn���yU_tK����*�rmO�7���۵�{�Ն�   ��j��yWum��4���k�I��u�]۵���w+4z�f���ew�<�YE}�<      T6>���YJ,�������ք�s�=��0��e��W    ��k�������%�̮3��ɔbv~q�"���!��;bSQ��Lb�&���mHuh=)"����	�a2�P�;�((׵=n[)nW�ծ�|l�ڞ!Z��ڞ���������2S����Uuf3?<\]]    DB�,�ھ>��|]l�m������`� ��ח��!�     @e�r��,S,��s����S�r�=%� gK     PG�7�Cּ������+�Қ�)v���x=	wc���@�N,��Z'���[�*r_�a���A������.ѵ]�6/���ڞ}>*��T���]ۃ�|^�"]ۥ@��j|E����   
�&�pm/I�_�k��x����T>Х�p��ȡ*��|��=!�0gF       �L���m� �fMZ�	�?&��f���Q�V�`�-   �D�Ŗ��l6~@��a޶jn2���Y9q�� g(�9n�m��!WS?vXX������aC�[���L&I!����	q���8��F���ڮ�K���Ο�ޑ��v��j<���:::"    ĴZ���Utmן�y�����L��A�|�U���H�[^�M�     `���@�sR��!���3����s��L�v�?Y�3��LgSj��p0   $677�rxI��`�c�*����M���l.��F>s�gn�;�5#��!���P�xnm���U
9�
�1�{n� ��ڞ&n�]ۥ::���̢Cu������w�X�F���FW#���%    ��NF��'pm_7�v�Jv��E��=D��{{҉!vl�)�=��=0�     ����z��H��}��C�_U��a�i��dB-�޵d0q���S   @�~\\�'l|�P��q3̳�x@"�(�T��L��UC���2��D�>����fl�q@h!6*�2�A0��t:4��b�LBqWp;%]�����e�UD6]��c�'�'�q�Lҵ]��ʮ���O��pD�;;    ����`!O1��\�>�$�v�C����9i��k{�Z]��ءW'���M��u�D)�Nʭ����X�     @e�L�s	>o�\�k�+ա�dU�<;�����d2����>(����   ����w+�y[hh�DLf�������������b��UC<� p7d8���Z܍��N��B���(����`aۣ�-` p/���0����>W���ι��r�G���um�(ص]����S�^�k��T�p�΍[    �����Ǧ�v���~�e�����0��E�:��߯+:1,2:      �>��z��������e�;�u��JN�����mnm�L��c,    ���6�9> PO`�e�:/LNK杧���9�d�����\2���~E�jՄ:q�6��&ĕ��P(S���-C���9kby����
pm'��[tm����v��{��=lgI��4q�*��]sN�y�um����]��C���y   @f�����^�k��/ee�s�4P�k���e\�yF�!;��!�N�N��      ������g��紂v�LSt�j�xeU)7�F8�\�s]w��ԓ����=�1    ���_� PO0������e��������]�Hx�=5j��P>r9aw����/�7��h�Mi(n�E�������0��KKvm����vmO��tm�}�:��=�k�\��j    Dvv����}�3��l�p�jӵ]Ӭ��}Eq���[�k����n5�,�*ωA�$��|��C��       4���F�.!�_�|��w�� U#Sh�|9C{\A T[���&    ��\�@�;?ۡ��Q��5����Y�A��H?��c�*�3F�������o���r����3(Q���R��5��bw�B��8 ����]�CL]�}Eٲ��$ճ����.ӵ]��Z    �^�O�	��Y76W���z�v�����
AH;��Ǚ�s�*9)��*N������Љ�!�*      ցaV�M�ļab���d7��	�,Fа"�3����3C TW��)u��3   �;��!찵��=���F�{�a�#w�q�V�{~4�F�LڝvꪈD����SyTx`j�����%P>���$�.ϵ=��%n���D*q��k�ԗ-����)�^q����!p   ���G�q���y����z�����k��ڮ�:�����N��P_r܃�za|�k�<�-vI���       � 3��[�D��.q�{���I��-wu0q;�(�1@     �F`|k6_�Rް�-e�_ۆ<�V���/��s��|!W�r<�& �{:�*����J,����Q�*��H\(A0��0�.�j�k����ȵ=^���c   �i�ظ�\��x��u���k��
w+���o5h�����Wn����S?*W�������܉aM      4�`���	��屾8�O�V�#|͜dM�ۋ�-���7 p���     4Ƒ��v`:O�d�N�;�d��wf��^�Njr�g�.���B��&���f	7��	q�3)\�(S⪘U�����!�ˮ�ĉ����\�#B�ԎPV�k�ܽ���r]���a�"]��Sl�[�0l�A    �i����"\�M��并��˴�uvm��k4���l��o5��@ռHw�'�+r3Z��Pџh       �`0���X�+�3٢{�A��oo���E��L��g2�1^�?/   �� �^o��nf����C�q�"g��B�Pz.nO�*3<�E1p��=�N����Ѝ!���Rߐ2�_���,k����m�s9^�
J�ȵ=ֶ�����]ۓm9pm���}U�v����3��͛p5   8d'���V74�6i�,�v�x4(�f-HNT��W�$�
2�+R��=4%R     �p5Y��Iqf���u�_�,n�jn0�]cY�5w   @�Ÿ��[;���X�ӭ���A�\_�����34�<b�Ӧ� �{ڭ�i���v⢛;&]���Q��]q�u�w�T���|?(ӵ]�N+��gԉ������=�'h��ӵ=,c�?�t���  �l��x�(µ]�@��4�vCq{IךO�nVw�v�����q᜷N��8F �����zb[r��m��4      ����t���ũ��w$lOI\7E\���yC;\�  �3�ш��~`�   ������@}����{5�j���>��BS��V�9���\ix���I�, �Lp����`X�f�����<��tmg(��M]�5�\�e}��	������U��Y�{�9ђ��a���~B�߻���/�K    �N��Ksm_Aܾ�k{�y���QWI�uu"�������gaA�U:Rcܯ�@��~��'      @���:4�ƻ0��ƄI~V�Z�<R��6�Z��`���C�Uj���}�����k    ��۷����@}]b�g�uA�.�)O�Mf�fX\/	�U9C.���w�)@��ߋ_.�M-�S\�n#�5!4ugpd��r�B��0�h:�R�n]a���9��u�B�k��8U�n�ھ8s�����g;��ג��.����8{<��hk�E   ��������i���sˮ��Z��s;�//n_յ������6��|�,�wU�*��'P��A*V3      �j�j�h:��%T#�D�����)V2��k|�����w+� ՙãCzt�.�   ���wn�/���@}�0����Ύ�����v̷�Kܕs{NG̻���1��a=��Vw��o��r�9*#�&����z���cQ��H�n���-v����,ѵ}�w��]�))_ڵ]rcOз�ڮ>��\ۅ㮋�|�   !7�nқ���B\�U�õݬ#�-�������ŀ@�T5Pe�2U±r���q�U      �-{q�u���0�����'����3dl��
W���r|rB����	    s�wvhpqA���9���@�4i��oڬ[�.�����4"�pݮp�s\��vs��͹�����V�-�M���X䮉L���C�������7Vwm�K�����v]��~Q ^�k���#�jv���L��G,�;�a   ��v�[8Z�v��sm_�����D�1��A��^����!P     @=�Z�x�N�|A7֟��#�	�'U"w]�`�4a�s�ilC�n��xL���I5e6�Q+��    ˏl�:���l��g��k�"ͷ��w?�a�-��-�'c~�9��\i����U���`��������Uڭ�d��`ss����\ t�vQ5N��m_����c�d�vm��z:Az�k�t���I~-�qm�w�   "�H�,��<a0cq{��<�V��4�����&�׉�//.	ء��*mP*�,�D�*u�
�*      ֈp���?�"Uݶ�QZ�����3�r�MI'���ሶw0�-M��      ��C��MY�,�[���LO9V#��UZ�לE����`<kQ�spo.U�j.ZO&��U��ʘ\�UYg����7o��0�2�n�L�vr����EQ�����}M\ۅ��?��n�   4���F�!���k��n�v]��6��_bIk42P�,�>����f�"wYC�	T     �.L�v<~'q�*I'��|nn �S�+A��U<�c,{0!��N3��    h8X�UkF�!;d�������yp<���#H���yY�<���7��=��6��U喃~�+�g�B7fC�}�6�Z���o�����u����}���'n��C�޵]|�tm��WWWt~z�i�'RI��\�Gz$��������Xj�\�������$k��/��d�J�~B}��P������)������jъ�kg�<�q��_^^�;`K��k��9W�O&g}3\�������嵳��3�a��5p���~4����s���ί�#��Za8��6��m'�6���Lo��?8;7vw��_D��˜���Ճ��̺M�<�y�d����ɉ���s�4�<�7n�>�� P�+�T�s������b�8f�;      �c�/v~&1�����7z^h%eq�^�����v��Ԙ�X    �0�LW��h�q�-�0_K���8�ǟ1��v�����%��3���=��G[�`=��O:�II��F\��0��L�/���C�j���_����*�^�\�^&4qտ����1���h�P<(Ҹ�����΄O�oފ7/'�W6�����UH)<9>&6���U��PInvN���oG.;=9���_��ӞuX�P�s'��B�������@�w*,.�����Q`��3�/�����J�����&^����=τήv�py��]���N'�q���[�}��oo����:8:�%�6Ջ_\��{�<|E�vS�{����mj�Z�P(e�zv�{-s�|u��	�ٜ������\��]�-�(�nݺ������t��.o��
�K�7k���     �c�Ue����Ry(1�,˺�ӎ���Juqg;�r���Z</_��j��{W�����7��㓹iE��\pq>�~��9������yS+�p.����>���\���f�k�r��_{����A`�����}�̙�!���Y�.M ]�w,o���������[&���O���_��]��{���kt9��S�c���C�c|vϹ�[�Q�yݹs����*�x��������y�0��MG��ae��Ϩ	@����أ��c���7�ue90�n�Ď����	1����ࠔ����	�\�g���U��O���{�&]�tm�cA�O?��X �s>7rm��3��Vp�Oo^��W�?|R�k��v�Ne�����(�De����O��a;Ͻ[w��l�p��=r�l6�P�M�l�������%��g�����+\�w�lQ�����{.py��g�Cl������l]^;���W�����MP]��g�$���G�Gt:���[7�-���svzJ}�qf]��\'"7;/V���?���Q]�����O��{���R��kN�v�{��)���d��rn�FY�
�h���gM�#:%UIq������0�G�@�/-x      8g<��E_�E��X���(U&�u(�ں�6ff�Pw+K�biL|�0���,D�vߟэ�{V�f���'g���a׽��C�H���֯����g?��~��/��]�.}e�⸮�f0����Y\jww�I߮_{����<�[�����w�q�?��{ޕ9����]3��7���u�i���}��:|W�w��ɩ�1��8#��7��햛�����K�c|��c����Ee�yX��h���D�8@Z��i�C���)�@��8��*e��H�jP)p��P��J%��UpP(��P4���_(�r�i�	ѶFHN�]�ħ	ă�^��=����[ �Nr9a����m露���{�>�ՑNU��|���5������Lq��^����  �n  ��IDAT �mn޼E��pX7��\�j�dX��t�G����<��4&�W;������	�A��`��V�U�/��x=�����_h@�� ���     `]�<�h�������:f;?'g���K�ܽ5�-�y($2�T0������U��3���b�n�k�?�^�G�����;]��>^����G�����v߻�����g�T쳯�������"3csտ�����L����5ؕ����.���{�>Y���>��^�S�wq��v6�`�g�t��X}�c��]�����|���>���<�p��}�a�0-�m:�Ͱ�T��D�0�1��.&5^�.�{�G3�;��q$�WM�6B=u�*!tc�(���^7�2�۷o(�p��u���(�k�P�8a{�@<�k{�?��{��G|���BJ^sY����(�8r�   �D�-n��KD^��� �vMFuWum��u'�??s��aӸ{�n��+��� U2P%
�S�}��Ѥ@      ��ńh;�r�TC�y��� n1��G�r��:��l��3��K�bpA��0��v2    ǃ��v� �s��Ma��2̧�b����
G�P�.�+���1�`ܜ�.�\rp<��A�9^Ȯup���bPkފ6q���=/�!�ځa���dsy��>�L������Z ��W�k��������\ї��]U��r�*   �-����d}�.\%�_M��Sߖ�ڞ�g*n��K��v`�4~���n��'�L��a�j�w�^�xI����@      ��E����M�d�g�^\!s��� �AV�w~f�X�|��r�    ���M�\`\k��H�J��Bm��X~.�#�����1�,�o
��`<����7C�=@|c�7b�����*�;Q�T<{{{�0\��M��.˵}�c��5��'�6qmW
�C!yѮ����Bv�q)�v�8Sa��n�Iާ��A��Ǐ�/�    ��0���l�x�v�)��ȍ�jO�������*ܺu��A"��^��R�┸������`�|�A      T���O���z�O䅯IS,mB\)lg��Bg��"��� ���3#e�   ��t�]��	�6�]	��2�4�"��P��I�C��}~���G��4���z��ጚ�9���4�L�`C�;�}.0��v@ws�V� p����|!p/ɵ������\�E�wm'ѵ���s��g�۽��?E�^�k;W���>��C   �
[�up|�|�a��Y�0��v��e����^�	�S��H�����a0W峎�����(;H�����0��ے��"~�?�      �Z�\^����1}�N讛7H	l�����v���e2��x<�_���;x�pxxH   @y��!�y�O��/.i6k��%��\-��u:�0q��D}Ew�;��	�$�������/��a;D�*������U"v��� �*��A�n������>.ϵ=C ԥ�]��sҜCQ����R��B�
�zX�Ե�/�N����E   @Sy��1�x�J,,A�n*l��5�W׵�Z�{l3h��`}E���9>+� �x\����]�ڼ(��n�`dW4      ��l4��v[X��'�u;?�[��u�V��s��7o�$`�������]W^�yM�<�/���   �&���#��_�;���]���N���<o�;^��*����)9v�K����e;׏O�1@���V�+��P���C�0��Jv���ba��+r��U<����K��������$\ۥ�b]۽ص]#W�{q���N����.p]���i  @s��ؠI��]��=�r��4�v���k�����	ء��4�@�i�J�DQ�8X���ɟE��      �I�z�.��&�I�[���5g��Ur����bp�{�9=;�O=%   ���7�4	�c�c��aY�Ue!��)=g��J���ۻEe��\����S���='�V/Le���8����3X�%+ڋ�W��[����$\�Sw��tAz$���/���mõ]�w��n��v   �(Z������j��F؝K�nV����U��������*����-��MԋHĸ@|�$P��:q�P�S�׬@      �D��[i��x~>gu��ynܸA��՟r�   �3��-�vp9Os�w4���*�h�;QjA6�nw��7��='�3�iHT�spO&��*�����"\<�c�N�����\�v�޲��~���W�߃E�����L]��g/��R��M]�úY"���(p�   ��>dcJJ�W���ʊzza�Q�"��D�Zq��9��+��>���w���|�Yg�>��p/����2~�O\�ɏn�Tq������      ��x����} &�s��崉d7v~����G����)��T#�   �߃�g��5���\���;&�s_Q+�.�R��a�0���R���='�Y�Z�ʈ�{��7n|��a���ʋ� ���N�⾿�O�\޽d��P쮪C���ĵ�Vvm7�Ǯ�gu��M��SM��tm�pՕ$Z_A����"��5�N�3�H   @�w���
e����z"[[�v���	ֳ:��\�u��߿OU�Ѷ�^4V��sٹ����}�֬լ@      �=^�r�X�<o8���pʡ1�r�34���"��t�o՟�hD�.b   �s�>Ů������6`�R]̯th��F"��D���q�K���d���g굩I@����E�aZ�Jn5 mC.܌�Q���~��/�*3�S���9m�A������&�1u�=#�����a��
�v��T�k�ԡҵ�TBrJ�G�'�������+��E�����l8���V��   4��}���j�m��t�
�vsq;��o�������(�~�Ow��u}ne
�{H����~tK��'�O�      �Ʉ�9�IIg"J���ɼ��9.����Y#l7ŵ;{0�{�ӡ1��AP����+�s���5   `�O>�����@��a�������V�l~�v|�pY����DjG��:_�I�1u�c� �99�"�$�@�p�rN!��[�����E�!uP�0w@`���3���m��8�v?�k{��<�_ڵ=!ʷ�ڞ�����ƹ��N��;  �Ʊ��M�W�\c\c�v�~5�:\��]+;�3$^�������0��ڭa��>*�ىRp�
R�Q�JC�Z���,t3#      @�Qgn-l%a</���$�ک-lU����)�e��s��ǳ��|��@�@T����^`�   4��7o��/��@}as����@�<~��z����\�U�st�X\Ԯ�K�ܵ���ߗ3f�5�� �{NNFD��@U�C��=,�׉�V'ǣ'Q)V/�o]T<�����(^UU�k�ؖ"��pm������T�v�8_�Vi��}��ڞ��V+p��F   4�v��kA��\]YQO�7�[	y������h6� ��6�U&�������mpA*��e^O!nWa.��z�       1���1�"�<�3e�ga~`��sx���"��(2��j��y)��3�L���6�6	�f�תЇ   `l�Z{&W�J���f���:oXt�Qg�g�3�����:=q2w�ZH?C�R8�����U�vn�|Ω��rM�*jK+lgTk�Y���m��prtLk��N��<�o���a`9���S���O֑]��kΉ�wm��m8����_��   �&���K�+��]Ʈ���fus֋���ԝ�ھ��}y���芀�Y��^[��G�dT�U\@��(�b��{>���      �����^�+����@7wH5��Y�Y睟a�Um�g�ל����-�q  �����G�1�z3�B��l���T���G}nҜU���9���ỳ�p���v��f-ހ�='��)�6Z�d4C�&:��n\��:煺�Bn߾M��G��U�k���^�k��ܗvm+Ku����\۹��hH>}
�;  ���駟ҫ�oR����\��޵]]���C�Z/�	�l\����6�;��7���0���G��     �t�x�N8�'�b�路�ȹC��Q��2�Z���ݻw	�apvNw�������>~���[   ��G�>�_�ｺ3�B����Eb�P7�����Xa���珇��|ߣn��L>+��~x��oF_���|�g.�ͷ��:�BnݺE���2]��B���@��Ĺ��˩A��B���666   h
��ߣ�����Wwm_M��^D��8�<�}�6!p�GY;lUm��u�J�0F�J.z˓1Y��~�.���       �F0^����$���8����a����'!n/~NT��"v~�����zsxtD���w   ������7���@�����h|�0(ʘǫ4�a�P#�Wc�e��7��}	���jx�8��*.�E��ŉoy����VyE�:��
�f+}����}��k��,Ӻ�+�J���N��|�]ۣs[\e���v�   ��n+˝���[��������.�������m����$W�+�8'�H��	P-:�T쇝��%��      T���)y=/�x'���b�M.T�iq�]���;7�z<v~����ug6�R��%   �)�q(�2�g|��-��7�I�7u��:-q��_H��uixJ��%hw��_^$VG���LZu�'��P:2'r�Q���������|J���4p����#q��k{RE�8.��µ])�V�#��'˔�v�/G��.)�m���\/�ѣG��w�   Pg�R7�L��1�kf��\��ԭ�k;������1�#���-�:�G�91h�T�"���M�C�     @Ua;?��}����j��=�.�͘K�c�~�;?��v��|�;��4L9�TZ%�   �
��	��&0b�g[d-@�s�0�|r����c��9.�����K0i��N�k^��)��!�O��M�
Ri��<iO�k��n{{�<x@/^� P>G�����]��d�U�v��yF�:���ѧ���   j�G}Do��G��ڮy
�/^�^+[�Űv`� ���u
F��p^.�wb�[Q�����\ݻ�M      T���&/.�c�Drz��b� �eeR1��]G�s�,g���������@}9<>�   Pg>|H���	ԛ�xwK�y�a�n���9��4��	ۉ���ߠ���\]�l�H�����Mɉ��χ����C������z��	�8<8��ˇ/\�\����k{X������텺�S���<
���v��N��{'   �χO?����7�ߥ����k�YG���u��tz|L�,�i�W�`T����]��W���NiB�c�q�yN      �^g�z ?H��DD��ryC?�F���w*��]~*m�S���Wm�޽{���Iʅ��g紻w�@}�Ջ��O>��  @�y��3�����@�9=9!`����ޞQݦ�u��E����$f'}!�ݼ�!�K0��i#�"��=d�7e��޼�*���љ��!@������w�R���?]��d[��v�k{���]�)�Ni�틺�\�墍�M8�   �=�~?XإB���L@���q�rD人Uܓ��������nG��9��hn��()~j<@���D���G      �j3]���/VM3Ǌۜȝ���d,�5H�/3%Z��b�ߧ�O��_|A�|N�O p�9���vo�   PwX�pt5"Po���y�X�K����v"}<@#j�bW�B�ǣ�W�ىH�
�����Nت:P%���.�g�&\� �n�a��b;��]�=y/�&����������kT	�UZ��:��A �׿�5   u����ԟ%���j����4��ԣկU>W8�ۃ�U$U۲0�-�������PȞ���~q��s9c��      �ː�ۥ1}�7#9�'M�PN|��yGy������]G�r��w;0��#����#   U��GgT�xT���SvX&o���[Ǽa\7+׭��B�.�-
��5-o������=R'��d5qu�d9���!l7�� �*mC�n��7o]�%7�EY �N���E�*�yY��:Y��j�������+(�n���}��� p  P[~��ҷ�^	ej]�f���`�y>a�j��r������><��ɶx�葲|��Q�m'�!�sX������E����lܼ@      ����M�)�z"��?,�&�bY>�m��e���s����?~L�p�lo�޽{���O   @a$�{��@������W�yC�����=��b��Q��K*?5/o���=��o�R���"ǅ0�-�[��T:�*�Vi�M�����hl��л�K����.	�%q{��z���b��
�e?{�w��   ��r��=��̝���j���P�^D�rD�UܯVW�Z�ˎ��ء����tI~�yT�ށ-�&�3F��Ǫ.a��j      T���G[|Z��V����C!�-΋usa��{��v�1�c,{��!�?_��+����=�  Ԗg�|L�?��@�������~)�V>o���6��#&M�@��~X�ܽ�@����F?3@�'�śS�s�4t�*��*�ȕ�"we���h��ӧ�j�h6k�
WЃ���sm'� ]�72���M��k;���d�2]ۅ��ybM�k{r��ڵ]�<���-��ڢ��   �F�3��uպ��f�u�k�a�e������ת�{�`VW�Z/*��c�����6���Zx��ɽ����X�\]���㓿��u��uq��9�      �ڰ���f�b��o�~� �+TDnqr���y�����J�w��%`���� ?�򴠾�[h~   ԑV��Y�N&t1��P�\�|.K�ބ��J�+�O�J�|{B\���=����o��r��3D�Vn��s���L�L
\��/C�W7o��o޼!P>�����#i{Gc���3�2�1A�^�k{�i/!�^Ƶ}�z��e����^�E������}���   P'����ٙ������8�X�.U<|@�l�ɶ���kB9m�/�$���?<��DN������.��.�      T�w�3j�l��}i~@~���8�ķ2������V��*��p~ZV��0!���ݸ�G��\M'������   �:��΃�%��sr|�9�%�|�ɓ'���a�����J�I�7�ڑ��t:t6j�Bܗ��'��<�bh�U���p�E�*����Si�*�Wm��nӇ~��%޼zE��{�;P�k���òk�\Y��S�k{��]����ڞ�X8��z ���C   ��g?�����X�����nMD��WQpO��f���@�n����Lw�5t	A*�Bt9������ƽ=�$����&��v      �Δ��76h2����� �7$
S��"D7៏r9E�:��[dw�6=	�������o���}����?�9   u������/	ԟ�Cv���-dg����c伡����c��!505���L��^Ȯ
4)n�P�>��!��<J�pZ�\�tW���ӧO����4m�7/_��(ҵݳ�ڮ8�[��]��'���.���܄�	  ����dI�I\��hµ]�Mq���oVq�*���裏���m+����{�q� %��k\?��      փv���3e"��NVS4_P9�e��ù��;(H䮣
�E�������+�s|xDO?~F���{G���o@�  �v0��_��?la&���L�n7z��a�w�$fW�de�۝>5ܗd�w��U���.q]~�Bw"i������Q������vx��5Mg3�[qኮ���`^hյ=������9�F��+�v��{=.//�����   �:�v���_�Za��`=�k�\\�����{}Fm�qm�K p�I�cQi.���=��H�ߩ��ǭ      քv�z�=�'._�����OL�E�T�iO�)PO�ȶY[l�g�� '����	   �l�8#���L`��Jސ���!p98�h;����ȍAvb��A+I�k�� �*�>z􈶷��(x�A۴Z�@|�~�����ǏL�[��[%$O�������뗯�����q᭑�^1��e������~f����Ǥ�ۗ<Y�껗����D&bt�/pš/_|G��W�n������ϩl�A���}���Z�N�Ex<��Ņ��ٵk�W,prr���F�9��嵻���l�.�j�&.�������Eq������eN�p��O��`{���_���kp�x>��<������w�����r�i�S�������ſ�<o��'r}c\W^^����ø0�)$*f�����9�˱=�u�:�</�஢Lׄ4�n�O�����n��M����: -�W��=7ߡ      ��L�^jr�T�)]�Ĺ��%�*2��T-����G�7������ݻ���;   � �^{��5����'�nt!M����@�0��R�0,���z7��`H�9�e�����/����▌D�eǶ��+��~��I����t�s�vEֵ߹���o�(���Έ�M�2&n��?����a�o_�~?y���v�����П�ş�'�<S7�����㿡?�˿�ˮ�{@����Qټy�nݺ]��7�гgϜ�̈́�Lpz��='�����>}J�`BWW����q����=��v��� 8�*���iypy�lA�۷o_�l��ׯ�Ν;��|����g����*E���A]&n�!?6�V��f��/~�o���=�v���� X�q��}�s��3�������5��ؾ*��(���Q�Z[�Ґh.�A<�W��x@�����l�      �>�~�<����'�ùH,lO1ÒY��9��P�W��?�E�1����U<��ڿ����~��89<��̍�����N�N��u#�8=:��_~�of2�����0*��W�������ߖ����9����ܸ̞4ܜ����]��v�9ˮ����I�gggA�M4g
��\�N�y��8_>����Ɖ��y��_.�wt=Ʋ7�G���H�?.���s���]}ޥQ��Rւc�S�S6~qc��ܗ��O����vn5��Ɛtb��ԫ?��w�殐&�b��Ѝ���7o�7�	�"�(�D�J�׉��zi"y�P���|,Y�D}EJv�8Sq��"xR��}�ci5q;�b��9�gp�w�E7o���   �:þC[���`]W/_�UE�y�_}^��ˮk*lW�8�{��=;����,�ܪ�Ӷ4��V��XM�Ȃ�<�����?      jN�Z�g8֏P$�żaXM�FXq�]���jn��Ç�P��ss%<�&�D���k��ݦ�O�c����o���޾|E�7�h˕Q˗_ӳ�����00�x�Dt��?��?��������l�r��3noo�I�M~����igg'0hr�ks&fN�j��/_&*�v{w�ڳ�X6faN�.x����?��?��_��pK���y���{���펽1֋_=ƴ����V�666��})�ua���;_g��V��yãQ3��/����;}����pÆh�]��@��-���>�&LT��W_(�W߽�(\������T�ĵ�O���*)�[�k�'��e���da��=x����o-��������ߧ��o��   �u�g����n�� xl*B_YOe��Wܛ�S��y�~�sUUֿT�g�c{l[�����,�dߑ!yK�v�"�%��]�/�$�g����98      �xޜ�0�'ʄ�v2o��[+���|ar|e����ǇG�	�A������[!   `
ә�_^hǇ�ڂ�?�����������z��W`cs����"w~F�ffdz»�0hR������=�-������Z$�Ƴ]�)ݑ=���]�3��&��K���(����28�r��'��Z�v�̣���H   �����'�������RW0�;�WUpoxR����vm�R��o���G}D���Fu����Ϲ�����#E񀤰E��a����f�      XG�;��g7��{�>o(��!)��3��<OS���U�-2�۷o�{��f&p��g��9��G�E���H   �:�����_��6w����r|tL�O�<1މ��y��Q&yì���=�P������Bo�f��vF� ����58>=*�7h�N�+&� v`� ����{�/7�4��)�hE':�I���TKݚ�3����={�������|؝�}f����}�Lw�{Q��#)�˰��@nP	��HD"��D����f!�EFJ ���c�f]&)�k;�qU�E�x���q�e�.��zX��\�3��������"���� �B���[U�cb��ax�"��	���>�U�~��{��$&������oDG�����`i�}F�\�9 �XEgklnEr�4cqB!�BH�YM	c�f$	��ȍ<�Vdm���e�gA	�n��-���R�|�+���E�hB!q���+��h��1�$�N��Q��P�mM^uC��uк�1Qy�v�XF������ ��,�;�~dn�X�H��AٳgHx�d�Epmr�g�G��X�c;�E�յ��~.J�ڮ�[��3����B)G�;����]�zQD�A����kwC��V<_��k���#���uX2Ѹ��_I+���9q���$Uډ���B!��򢮱���ܽ�kIqU�����X���)�b�{��A|��� �gyis�shmk���-ΧW󛝝!�R�l޼3ss ����4VWVA�a����yM��q[���u��a}�Nա�= s�48�S�*�+p'��Y\I+k����W{��-�;}�8u�L�\۫�O��yl�cP�\�e}����6hӵ���X?>f\"���m�A!��+��ǧ_}�k�!X�k{��Dܮ~�Աc#���d��e�1�T��!�$�u{�j=����RH�������B!��r#UӸv??�]����(n�#��8��P�>VQ�%r/������b�g
�+��~��'�՝; �Bʑ'O��R��p��0��uCE;���qܓܕc}eݰ�
�_�®��(�u��6{�*w���L��xg&J*F|�A�N���X]嬫0��ۭ��u]�AZ.煸������͸|��fl�]�n��һ�;��_۶m�r��B��$uU���݊��][:y�zq�XC��j��=��&c#� �JT��T�W��>�Ȏ��`O\YXYщՍQ[H�tW) �B!��X2괄�m�`/p�
��
�8����z+?�cmq��� �!V��{� ��gqqͭ� �Bʕچ:$	TUW�l|&�s
aP\(�Q7tO'׭fb��z/ݰV�0U���$*
��7���:�c{�vHUr7Y"G���м�ܒW�}b)4��ųg�@J���������T4�v�Ūr���p�XTZ�퐈��v[�W�����XY�[�������3����A!�����*z�}	�K""��)lW�W��u?�y�{�)l�+�SI8�	Ư��
�%FϿ�p#n�ds�H%&������';i^�1�m��5���B!���bj��ƺÚ֊�pL���J�#f�+�_��R\k���+?����8H�03?���LOO�B)'�n݊�	޷Tc���x���e"T/��!�1V��åVˬN,��:���/�P�������WQ���ȴ��擬N~E�P�z1��СC������o�oX�k�LHO�|�؎ߊ�sm�}8c��n�K$�ر�%B!�ƞ�/㇟��u���҉�K%�74�����U��}I��0?7b�������x�у�+��j ��{=^���HD9U)��e`��vB!�Bʍ�y�)]q����,l�'��H�s�)�¸
ԃ�Ӯ]��e��Sx
���ql5�P+���<Ĺ�'p��; �Bʉ�'����wA*�Օ�Nπ�Þ={�c06JMQZ7���t��Z�G�p=��� �U�n
���Ԃ��E��*8�t��Pb)
���0�����p$�1�ߏ��epm�]��pmw��+��um7?c��˞�k{���4Rx饗02BWTB!偘%^U-�7˵ݗ�<��� �T�ך��bGy�*�.i"�JT�,[��p_�j��[|b&� ����|B��w��T�v\$�B!�����$�HL��j��U���bY�V�b��`~�ul��0Ƣ�=�+��O`��m ���e4�4�B)7j�밚H�T½=
�c���M��o��ڻ�u��6W���̵���^E��)pHuCR���v�_��q��zJ�U����[�J8��������W�\��	��q�>Bwm��*׵��66>�3g���w�!�R�8q=�}���CB{P,D�q��ũb��)XW�l�ر�Q���*Q'��ݯ�r43W�Zلu�0E��r�\̤UcS+�����"�B!��YJc�f���ܽ�XN�sl�.r�c'�63X��ݤ�̯���o��$&��(p� �fg�y�fLNN�B)�����H����Hx���+�n��<U�P>�]�9�M--HNUnݐ����޽4�����u�1��:Kc�Ų�>S&N���t�رȒn�HwW��-v���s��[{4�J�ڮ)lõ=ݳC�n�K&ؼcgzyI!�!�B��������E-"�S�T��K���>�~���P2�W�����c�A�����%9n\]�rQ�]w>��K؎�y �7��#�66�B!�R��74aq~6��i�%7xM�d��'���C�r�-�j�J�ё�@*��~ƥ�g��g��B)^;�:>��5H� �IxD1��S�0���&�K��'�L��m��U�(p�\�u��K/aeMRy�ܰ84��.�jx35�Ll�ݻ[�l�r�!�������ع#�k{���q$�k/q��k�뜊����n�K�^����{�����Y����x��!��8#܃�bk�s��5��ب�ŏ5�o��`]q���+�LT����x�ȑ؈�u�wN����Ð��q'����
a��9�M�{���B!���$U״v_?��Ȫ]34��ng�Љ5�`X7�Y�p��&PzN����0Q+���467�|�BHY jյ5H&� ���?��i���JQ7����w��p���� �a���:Wzݐ���Wc�Y��tn�ۭ�n�� .#�/��lm������]��s���I���� ���v�ڙMf����Cr��ҵ�޴����vm��Q��k�����65=�#G�P�N!$��=����wD."W��Ϋt�� �T�����bĮ5��p�������8��r���m�hD9ݰ��'�K��<��7��*^�B!��#KhP��k���-��]�XV�AI	ͱ�Xw4W~nll���H�YZ\������A*�']�i!�ӧOA!�ę׏��_�>��&&��X$��� (i��E�ZU7��)�c�������k2��M�^`)���� ���;a�tb��JD)�W�$��=J�{��tu���鿳�vG]�m��q.q{	\��q��:E���������4!��8"~����HZD."����9��+���Ǫ�U[��8�Xk���0Hx���k�	�&��֞��4�ݞ��cv�DU6��pu]�(p'�B!�,�X�A�b�&]�,U�Њm�(Zk�V����k_KK:��������Do��y��Bbώ]���Jbt�u�0����겏�#Fף����p�=��=�w�a��T���Q��ܺ!��[I�ik#�	������"����3P�h7���<��]�U�\n0\:�>KO�p9�4]ۥbw��Z*l(��\�Q�+�k����s�+�k�3nxl.^��B!$�����\�cu�)L�|�v�� �T��A�P`�?���A����Rn�n��L��}�����yU�������&+7IE!�BH��b6�v�b��G��8�ǲ���!�e�B�z��b~�ū��J�{������� ����Rz2���<!��8"���fi�Xi���IxR7�"�5E[�б���FX.���~�k��B�t��E�����I�D�ډAqa˶�8�C���d����^y����NLL`۶m���]��b���n��\��P]��m��K$ص{Od�[!��|�;����y���pa����b��Vչ��F��w�1%��T�#� ᡚX\N�
��	���cҊʅ!7�ϵio��������S3�B!�R�N�prs��@��zM�������1��@��^XN�W^�X7
�*����gN��/��:!��xr��Y|��]��b|t$<��Y2�6��ۯﺡu��mR�ӭY2C,��]�7^o��o��te�)p/ɚ��jJZ��ve�� ��92gf���� �09K<\^t��������{��[���cG���cB!q���ˉU��܏�=��\%�5�)�rL��=�`
4������b�E������'����7�VM�n�q}�	�I�M\�B!��r&�v_��ڊ����_�,׸���6/�^��V�����	�ŵ�{~n-k�:�����m�BH���55XY]�������*c,ʡ����U��UՍ��j	�%�㦶v����(p/3�z�).8�ŘW����賛K�j�������}���8v����;�p��������æl*�k�zlY��{���mF�8�b�o����|<5=��^{�wB!�����x������\O�n(��/�XC?V%"�=���O�f�y^#C� �!&>�r��$�˶�b��5�Sg�w�,5��k!�B!����o�1?o���4��Z��qG��ݺ�ڇ��Xn�W����W_EMM���^�=LF�F�r���J�yowZ����B!$N[�|�����B�"��8.&V��V7�����{��S����z��KoW:��х*�r\h�|�s��q�ex3���D��
�NzQ�.O��Y�f/ĵ] �gv��<붧�]�]}����˄�A\������
���.�3��󿅁����@!$n467cee%�8L���]u^��������X�K-Lp?��b�c}}}�q98+�"�ב���8�O:����I*�C&a��|R��dB!�R�,��6�Uo�`�p��:k�Yr��b�u8c�(�[�lI��?NaSXAсï�T�{��浛�B�{^~|�	He!&\���X��}6�
�.e�u�mF�qzn��{�d��Y����V�
����)�l�̢(`�A��]'aeub��G��E!�+1+�����"FF��c�N=�v��Ј(����ID�"xw�����*�u���ΰP\۽D��F�}å˗�ч�B�G����P�q�"r�
[�S8�����P� M�z@��y���bl���_!p/&qOtY�Rִ�r�r/�K�]KY��B!��7�+5hi���A�Vl�Κ��swPW�"\�)p���A��c%�@SSS�nL!��a�8�0RY�����Hx#ⰈCMѡgϴ��9 ��N�2c,�6�$�����.�а��^��qq�n�<�r�t�0�C
��'W�|��-� ����Jܵ]��jC"�N����8���cU�v�!�k��+�gc)]ۭm��v����k7����?��BH�>zw�>��R��"��\�b�4�)�+}�
��/5��^$�x/.G�>k2�㞠G�sr&�I�J5�<7n�'P�&�L��E��3Mq;!�B!�Nߌ�W٪My�	ʱ�z2�5ga��k5ȉr�f�P.�򗿀����"f�g���R9|��G�>s_ݹB!$�=w�>��������MJO��q�)�8��_��~��Ms�B�T��ɣ��"��܊��i�������� �*���%�u�t��y�ɑ#G�i�&LMM����'Op����c?��6��C�]��*{c&�p�vg�/�v��8#Pl�:��6C����ə�A�Yܻ{�BH��ر�33J��4۟0\����4����y�Ā��u�8_��4�7 ��88$���0W"t��6��^cxuK����؈�N� �B!���N��M59a��K�f��*�U��F?y��q2�
��Ƶ��Q���_X@k{��!�Ă���6�ayy���{{��q�X1+���a��4ho+�k��f^`�����4Ƣ��X$j��2����)(�e�W�ʌg�K�I���Z�8q��9H8�<�J;z�/�R���+sm�v{<�P=W��r4�]�ak˵�u����#�6��:|��B"���s���GW{iD��*v��^� �c���u��c}��}	�s����Ƕm۰�~đb%�̱��M�y$�;2X������B!�BH��\��onk��kb���"�е��1ctd��k�AꇢfXWWG'���W��T?���O����B���gN��H�120---���͑��P����U��f(5�b�0�Eb>U���pc(l�_��Ȋ�s1*!kT"t?�
������H"�@_��]ǵ=���܏`]*:7�򸶫����~����킢����nH�W���'O�>!����XY���K�NDn脭7_�^
�ZDP����M�󘙚	�ӧO��OL��P|,��R��>�&��ݜ"�d]3!�B!����{Ø�Nn-�f�[^3��#菵�ʤ�h�'rG�U�~	�ѡ���V�y��adl�^}�wB!��y�V|����Bh��G�@���ɓ����>�Sݰ�5E��=7��z���]O�r� Ǻa
܋��Bv���B������a&�T1��C�b�N��K!ɫC�������Y�{9���D��vm�ƹ��7�T���ؠ��p�NNO���S�B��KW.�g����������avX�u?�y��*��yP_"x�dM�� �Zf��LV��s}�=L뻵R:I*�x>Y�vd.�M!�B�F`��q�^?��઻���laݲ�c�O��O\�pq��=<Lq��/�T��}8x� ���@!�D��c<���P%bN�$�!��@duC�x;����˚+X��bR�u
܋ĳ�$v6���0���$�&IV�b2��>�quW�O|��%iV)<}�o����]�a�Q�#X����8���*�A{T��n�W�����Z �{Umv�܉��!B!a"��������j��X=�u���"�b��W���C������=T���Xf�R�%����O��'�e�J{E�u��HT��|&�!�B�L�Ԡ-eX�d���@5��.n�aH�*��A��C�-	���!
�+�g]�x��-
�	!�D�������>�<��Y
�ÇK�����[�P�����uj�NSm��.���X7���H̯h�ֆ��{� ݋TZ,���N���!d-w�'Bl+f�?�$�����,��۳me���n�q.Ѻy���smwoxt/_��?A!����K���I�D�Je��)�=X��k����Ep�X_"x���k�߇��R[[��^{-6���gMPIw�k��=�3Q�˅��3H;���B!�����I'�r+?�c��-JͲ�cG�K'7��B�	'ϸ�47*��8~�H�11=�m۶all�BH��ڵÃ ���"�W�P7�����a�I61ݭ�Ͷ���m+�Y��'(nP�^Dj�Z��<f��dK
�Kz�`��q;A�~VK��+�ŝ�p�|։�����.�������j"l�vm�r}��pmw�� �D������bnn�BH�ߠ����������@�v���� ��<�`]3Nլ+lwƎ�`yi	$<��ݖ-[���\*�>�X��ĐW@R�ř3him��4U�B!�lg���RCV�n-T�����c˄���y&�
�!M~�С��vtt$&�'����ƦF��⧟�֥���Ï@!��ɉS�����T�󘙚	��{���_�FB���[k� $cv��]U3T����1ɺa
܋�bU�t6���ݙ����Y����P
]��P�}���3Hx<��g�;.�wV�g�vC!x)�k;����Nq{�]��{7<6�kׯ��w�!��N�Bw��5��\���4E-X�ӿ�|=���ՍU�u����~�p9y�$*���1v�gfC5d�:r5�m �B!�l,[ڱ8;��甬 n/������fX���=&z�XUU�W?���8q}D�mX��~� �RY�ﶕd---���!�����P�4�>/X7Q���Ƣ6�*�>7��a���;#�5򜑵s\�e��J����Y74����/Vc�5Ie��N)��.�[���YŴ�>�ŕ���_G[��u]]����}�D[}�}�}���OP]S�~\��������O?����&V����;3�����ӣy<�gD"(W���U�{�������̿r|��Z�~��)�����<Z�[��ۛ�.�p}[T�������#�{uu+++XXX���ړɤ���1�����_Zw����f���Td�]�u/�w�{#�(���W��.�HDҿ�[\�Q}�}݉����aK�Z���]������Y�}��>�G�����ޡ;�:���8�������Z(�?��%�����<�W5�w��7�"Y>���%Q�����:v옴����V�}�q�z�{R�鞨?�ݖ�&�ֶ4��PB!�BH�HԴ��&�c �)��v���	��M�����n3���Cq�c�X����>�_jjj"�_���k��� }����=�
z�xݢ�����(X]Y���rd5�d"�k_^{������ĩ������~��[-E�r���Gտ��ﰨ���������BT��(�;�]������wͺ�$l����5�{��>�gΝ�W�~�D26�}�om���D��X+���k��}+��t�[���7�O��ߋB�a<,����k��}�nN��g<��v�4�r�E�ruH��}�ʘΉ������Y�nVq��b7����*k��mSUU�$���]�+�T~�r6�����ňn$���w�ٍ�G��$��P�����_����q��vm7����϶�rmw���$���I}�ɧ�q�Vd��}�	n���3%�g���~�ڽr��o���!l޼�!�<p�@$}����,v��I�bB¾}�Q��B`.~CĵQ����� 777k	SKA��]$����#[�kpp0�sT�����mC[+6@��\�Ų�{��)�Ւ��}� ���N�W���"�z�O��#���k�`jb2�����v�yyT�^������Ͽ�.Q;E��ԩ��y�pp/��Ai	z��P:��Dn�U����R��|�{J21~lI�gVA!�B�8L�֡�HI��~W�2�2I��	��5i/��Za�r����bbLU>M�M#�(��E^H/r���\ZX����`a~>�y�J�%���'VX���os[�&�~bGQÉ
!8�����{V,�~��_�3Ң����Q�k7E�Q�����wET�u�yT�]�-��Q���|�b^��~���c##Z�������B��'#��[Z��q�!�wĵ_,R�f�g��[���7��Q]w^��[�P�ɟ���&����.���6�,�;�n(����L.�м�	Ʉ{v���E�R^��͒���L��M�t���=}�tAn�p�>~��+D׆D8-�{�U�3q��*��<��nt!�W��V�~w$q�;���+����m�v�s��)l��󾯬���={�B����B*��������0�X=�u���"�����s��С@7��?]a�:6�6�$\�d�W^)|I����y��ڱ�S&�MHώٝ��+���f���d4MB!�BH����]�ِ��c���:�q���Xq���w��ق�4B��1��[1@~(�k����K�v�\����=�qʹm�@sDF-bUĨ^��Zߵu���O�V���ĝ/��z�<��Y�5S���znڴ)��+���w���i��(��s&��!�0�پ}{d"o�;�k&4bb�x�Q�k7�/�u�7������$����}��h�o��cwa�ܔ{����E|߶����Ezr�n�Q�ۛ��,F�ޯ���"��
Y�pV/�>�k��f��ayk�5��֟�5�	QA�{��oj��̤ˑ���>�%������rbv�s6�-�*iu��)
�C�������븶kŭ�۵]W܎*�Ъ
���^q�P\W؞nUL p�i�3{���;�F&�p��M|��� �BJ�,��y��v�����S���k���\�׵�J_��p9��kr��r�gx\��M��Rmv1Jʐ��S)�s��[�'��"�B!d��;��k�k������]�.���1F2��������ҫ?��� �1��_����7B����Bc,B!%���		#K�0	����p9w�\�Ϥ��<k�^�r�l9֚!�f������������c�P�^d����.�q��
��w�Ju�g?$�f�ʗ���*��
s��������Ȉm�����.(o�v�ݩ'�'Z׉�OѦ-n��2�v�+E�.�7	�=;v2YE!�d�;x ��p���GX�+l�4_�4��q���v?�������9���'I����WɈ��zq�J�a[�{�aMd�T��Ĺ����B!���Gr�~����s9C,Պ�V�6e��^X7q	��Ͱc�{q���N�{���σT&_}�-�_��/���BH)�|�
��p�r��=l��pe`�f���(Y�ݡ��S�S^� ��X�H
܋��J-�,�jg�ZZ�NɒUގq&2�9��t>=A���A��>}:=[O,�C��ɣ�i�����ϵ=�l�s�R��pm�ŕ�k�3ntr��x��!��br��I���ݻ�����}��Op���U�k`���1}	�5�T}A�~���L$<��މ'B�/�}����=�?^�u`0ۗ��Y�B!��-H�����]1nH�
้��L�l�w3���se�6q��s�pp�1V����afz�� ��pӭk�Gcc#���@!����,'Wi�X�L��c����#�U2�P�+�>Ǆr��Z��~��c�o���d��DMH
܋���NVIfWH�U�6庸��*+�6I�*��7��y(N�J��Ϝ9�/��$<���#nܾ�%:7��m"s3n������ڵ��~��u���θ��U��s���9��BH��Q{����g\���w�avp���ؠ"�u�8U�Z�����{��A�e���8v��\
�O༗7]�w�:I*��==q�>�����ZOT���@�B!����L��)y�0�����2�aH�t�C�^�z�}�fXSS�D�c�0|ч���A*�o�����.�O?!�RL.]��/�}R���L.b�0���*�ڠΊ��ڡ�nh(�#����87����.�N�ցu�����.lopϮ��#Y%��B]ˇ�p:0YA�I�M�B,�A�{���crr[�l�4d�rq���B]ۑ��µ]7�0T�b�����[��_�B!��>s�=]�u��X��ZҤ/�Kخ�U��
�u��Kp�>p��/�K�bYk*/^Dmm.E��RP��v�N�q����*^�&�$B1Q�B!��1y1W�����c���X�%z��q��l8��ȭ[��'q?|�$<�zzq������jkh�E!�����bae	+�� �K��p�����$�_�P�;|�y�v���=>�������v,�NggZ����\�:2�Uָx
�K�� 	��??��פ�s�k{�ܹf���l,�k���һ���S�i���z�`]ߵ���.�Ov�܅��6��΂B	���ڵg7����"B&���g����µ]}�c}	�5c5�Bܾ��De�qHJO4!sa�?&�wU�� �y����Q�N!�B�F�s"��Ȏ�u�|�g�c�<c�9��YV\j}A�99{�,�!39>���9�X�0�������|�">��B!��ҕ����; ����4f����ӧO�8q2�r���G��5C�����sʜ��m������Jd��I������ֵn2���ǒ�̝�D��!����KKK ����?���ktm��C66��w��K��nA�ܮ���������_�
B!$�ϟǳu�v;*�^A�P>_�W�X��\S��)"Wӗ�^3N՗</�z@�E�?~����>kj
J�v_����w��{s�`�B!���j�@s{V�uC���ڡ�.���Y����ns�8	�i��1������_�L�W���ʸ���́B	B{{;f��Ƌ�r���y�U�=}UU�����j���f(�*r�MH���朼�Y;\ۚ�:����@T
�����:tH
�Ra{�����]X�aKT�	��pI��9���'p��]��x�ۋ�il�ؔ~l
�]��R����������W�c7�k{����õ�~@2�D��m������4!��B����܁�.�v�[!��\�+U��Y�v�SRח`]3֧�^���_􁄋H���	���t�槠vbp?G1.�LTW
U��z�ru�}�	!�B!eGCR�sҺ�z�g��!nי��^ ȞBf��ĝ 5L��.�M��A£����
��{���K���A!�A��t�s�ʦ��H���ק�Sq�񕂜P�ږgܭ��j���1V����%��x�kSҋP~�z�܀��aG���Ǥ��,���r��=|���8}c�ϵ�&{+��u�ܮ����.:w����,�k;4��;��z��@!���k���E!�V��]M��K[5�J�\����c�����..\@]]]�q9'���!+j7���*���Dx"�ԮJT-���*!�B!��d��˙-��������1VX�Z�c�ر�'O@�cblK��hlj�LV	�$Wӆ
333 �B
a�֭����d�
gnv�SS �"�Ž�IX��(�κavlI��f��S�񾗸]l�+�k=r�
+����Zv� ��p]��V}q;g|T�wy���q�e���jߙ3gBs�'9��.]�\|�v��Mi%���%lW�mD�vY�vmw�'D=5u�8p� ���A!������M��<�:�h
ƃ�K#���+Ϡ y��Ԃ{�� ����>�Ν��3a��{�1�u,m}N^��c/[�-;���֘�!�B!���*u��X��.zOIk�^�XY�B��1�}w\j}A�9�)p�ߦ���z�r���{x��u|�� �B
���Kx�A*���^��9��vl���B�9��.� U�;_��Hyc)Vx{:Iͫ
�KDMSV�G�3.d"w�s{Jq�{$��[VPk(��a�$xQ�����mmm���,Hxt>}��5�ڶ�L�!�ѐ�����;�%n�ĕڵ��f������v��\�u����;cG'�p�����p�	!�_�z�6����"r��Z�d���ǪE䚂��"x_�{?�����h����Muuuz�W�u�Iw�ò�]��6s�nNBw����Đ�����nY?M��}�B!���N��*�o��Z�9;�P��������X�:FPs�BS�~��i����	�ߡ����i}�C�`?z�ihA!�G�����ԝ���n6bl%�U������k��K��9��ݜ�w�1��f(�mni�� �N(p/�h#7���\��}9��L�?G��)�r�~���>-����A�嗇?���˱wm]�q��������g��ݻ �Btعk��f����ڧ��������XC#������=b}	�5c�7SZOW����A,--��ˮ�ϠH{Q~I)�~2������`D�[*�R�k�T7v�B!���1�*4�n��씭^�9vȎ5�.�	�y�f��H�ެ����F���]�t	����7���������R�<�|�߾�z{z)P$���0�9x����G ����&�'@�E��~��ٲ���ϡǵ��}O6W������ؼ��%��\5�(�!�.;`���R��UI)�D���6��e�&�T��Ν��=�~�-.]��h���+��ݍ�8�g�v�k�@��θ��9=v��	+++ �B�q��E|q�kW���Ї0�8�u�8�X��{��vu���իWm��qHX����r�݉�֖w�+���8r3)Q�!�B!��rM��X`B��Tܞ�j����9\�ӕI�PF�k�^X���с�'O��o�	��������@*�����3g���߃B��¥���ӏ �EW7H����M�Y����vh�*�堮%Z5�*lU�P�/Cmg\�����D<M`oG���t^�v'����r�qHh�x1���O_����a�m��qrm�	��Bt��%�vq���|�����]�!�+��oxl�n����B!ċ��N��}�Z彟�`����u�0E�rm� ��^36��[c���zzA§���X�ڧ�^��&��x�D�غg�q� �B!�D��r6)��ұ�ȇ�P�\�Y>f�b�w2[��Xs��,��p���w���7:���^K��Nc,B!�hjjBcs3&&��M��'�{@�G��k�^X���v�p�to�ku��T�5k�K�ء��D����v,/�ۖ�9�e/h�,_��DUF�.v�~�A���^{�5�޽ �������mM7���{����3t�
tm��IK������ۛ�smwƮ��b�Νزe&&8� �"���/�ۋ����m���f�J�.��F��US��WDD�P���ɮ�Z�_�!��{؈�����c���8���xں��8���.�[��ּ@MM5:�WQ�	�B!��x�h,������%�mL�{�|�Y\�X���`���\#T�;}�4H����anv�mm �͝{����+��OA!�xq��5|~�k259���i��Qǳ���L��V�j���������N-�@��
�K��Ў�ܬbօ�蝛ɑ���)��־d�*�{��R�S]]�^.��#H�|��7����6�h�p���@۷k�K`noL��Qe_� ��|m�4N!�7�?����~b�q�øy�6����B!D���7���/鿕�����RN�
[I����
=�] �s��q�ر�3&�	+���'���8���U�b���}3��B!�R)L-&Ѽ��+�9�+����v����w�=��y�2�	.l/A�hlڴ	SSS �"\�_;u��Y\\�J2Ac,B!�l߾�s�\��}�>�v�±c�bQ�Y��RS,���*c,������S�ˠ�����ԣ�Zȶ�eEoC� ��eq%�r�&��qHh��@�{����ap`�v��
�%�k�F�[�^t��u7vC3�}<�bvmw�K' �vmw��NJ���j�iU:���NB!V���Q[_���y�}�R��`=�of��ͥrm�=Cf �����~��˴[٨	+�3'%sb�?�˽]�(�Kr��- �B!�T5M�XYQ.I.K����O�0�a��uuu�x�"�{�=�p�������������[x�wA!��8����C"���	�+W��W6���U�}&�ڡ�fX��۩�U��,�4p�+����)�uñ��b�A�����5�U�{��z�~�K����˨��E"� 	��~�	;w�;E�R�q��=�k{�/k\Vd�+X�'lw����\���a;�1��A��;&&'q��%tuue�S!�B�o\���?h���ڮ��{��]������j������B�.v�}^�+d_X���=�[-�U�Jm�I�#�k=��B!�R9���v��b]c
����cK�gѻ�R�>��3���Ħ-�A*��=�Gc,B!R�;�_:�M�Fʛ����̓�ϙ3g��q��AZ;t�3M^cn�~���i��z��;��D�Z�Թʠ����M'p��iA[v[gpd.�TZ�.�px�JTY�K��`1����;w��ѣ���A�廻w�߾��˵��h��rm�;.�k��|1��a�yč��.k�����7��'��B9z��H&��J��߬�߂�f����q��k;�b���ݝ�A§���ϟ/k�=8��ck��)�ߪD�s»�:�I�B!�T���ؗJ���e+>\�Y 3�rcdk&q�r�����_D��=��4O;���7ޤ1!�b��}����>!q�H�G8�_�t�,�����ܣ�@5Ô�_�8����p��9����ж�S�v�l����B�������ڵk�G���4�?��GC��.C%n�=���[�@�n	v�����
�!�X��%�)�o��Kس{�mۆ��!B�l���q��Q|�ݷ���������O�k���Bjo������0H�\�z�����~I喰�`q1���%�rb��t�dv�+csk+F�� �B!�TO�8���=!VR���+?��1N\m���n.�o��E��A�F�ݻ��� ����'Ξ.�$zR�|u�[\�v_|�9!������o@�@����y����*v�����❃E]�z���\+?Kk����\��P�U�9f�A�{��C�R�YQ{\��~w���]�*����%Ո>���G�	���j
�ڮ�]�.��G̸����ѵ�y���!��7��ÇA!�����m����\�R�]�߬�ڮ/�WtԵ�G�����g � �K2���P�c9�R��3�N��D��q�,Q�MR������M �B!�T��ܱ�3�Rw���l�m����i�%0�@:ò�8����7o�w��H�,.,bx`;��!3��X1رs'���A!��ٽg&g���� B�}XY^	�7n�ǽ����Cg���果�Q3����Ա�(��*(p/1�S�x%�t�u��-c������nXE��$��+��rHZ�9s&�=::
.�����G����R�q�v���a��[cumw?W!�7J��.i*����ﶉ�)<x��� �R��y�e�,�aii)Ӡ)��-B��TDnh�>�+4���⸶ku�!6���>b�A��U�L��G��\P�-HU�})k�,a�tfL%1���tp'�B!�Y�i[Lz���&�X�9����Z3��I�_C���/\��������!š��9�$����۷��7_B!���g;y����bҽv�H�G|/^�����<����O��v�f�|�ܭz_��˹��|U�Z�)9���g�xu[�2Q����3:���[��������|���U�sP(V?����~�:���?��K2����p���k��ն\۝q��yqum�[��mn~[�oC"����
!�T���8s�Lf�A���L\�3�
q{�#��5�_k9����a~n$|�?�ݻw{Ɣ��]�a��[�{���g�9(����<@2���q�0B!�R�����%�[�9�P��5C���j���1�#[�0�[��".��+W����333 �������hhh !�s�݃�k'=BH%s��U|��=b�Y�g$|�oߎS�Nž��2�Eǘ�! ��VTKY��)�ڡ� �g�������F�:�8=�JT�_�ܾl�5a�w�A��;2�X3��ﳾ�D��O�SђpD�����KW���umO���t����� �v�u&��Xw�8���>sS�Ӹ~�>��CB�,nܼ���vu�V1\�u�TD�K����
���E��N�h��V6��=_�E�a<T����2��}.Y��҂��!�B!�Ƀ�$~�^%��*~K���J�n��r�X&z����uㅸZ���}�]�p�q_w;
B�cc���CGG���A!��زe�U&��@�I�����E�͛7�F�&~kva����׏EU�f#��z�1�}R�uºs|�to����ӱUHœ$�!�Pպvq��MRً�)�Ca��+cm�&���FLZ	�HX---��K_?���c���cma{���[��pmw�\۝�b��rr�O�Ə?�B!��֭[�Z�ᚙu;u�Ƶ�_���Jqm�s^��p���++����1X����p���f؝�������e]K:Vqkh�B!�BH岚4�ھ��Z�v��ʶ�y�C�9��V(#��C?�/^��="��>����x1Џ����x�o�BHeq��U����A����.�h(�n�7>NuFk��Y3���녩u�j���c��6�oEr��v/(p���Z���Đ�[���%�Rz$[�ʐ�z���(��զM�p��y|�� ����������Eumϴ���~�9�D�n����#��ڮ�ƾ\�3�rq����,N�8�G����$����cW�_×�~mk7J��U&��~b�	�5�T}iƩb��p
��=G2�	�;v��2�A����ջ�d�-9eMbI�S�Ñam�2��z��;!�B!��r]���`���f8����s?"�,ֱ��6��ʵ~(��jjj������	LON�c3'~������c�8y��!����ܹs���O�����gld��3 ���؈K�.EZ,E�Q����=w荵���c{���U-��#��=������2J�7ð'�d����55;U�����F��^�~���)p��o�|����ۨ��˶�@\n��\���vC�\����hS��u��>���;��zWKP�OA�^$�?4��׮�?��?�B��F�={b�E(�k{i�tm�3�Z��=��A��\�,N?�e�$��{tD�V�H6����u`�nI<�`��B!��Jgp�[�IW�Pe���:W~N��-�-�1��0݉�
΅k׮]8y�$~�����~��/�!&��8z�&�;���� B!���4��a��b��Y'H4�U�6oޜ}\��A=�5�t�Ϛ�l�m�S��貚�������sB�Kc,/(p��Q��-X��T^�r�7�C��ڮ��.ITم��s�HI��W��~=�8�D�p�3��T��Va��;�urW��%m
a���zn�q���nm���Rk/��S���O ��1ٶ};[�1�ە~L�v"r_�u�8U_�q�X?��f���xz#�Pi�
�q�fқ�c�9+���Z���M��K !�B!�΃�q��*i�P9�VQ4wn�X�B�cE��^�c	w
ܣ��yN�;�jO7Ri|��W�}��{�]B��ܸ}��1�������^�h�|��vlj��9�e�l'{���:&�kcFzu�ǣ����X�nY�8��I*���ʍ!�pf���	,G��I&�.��ڀI�W^yǎCWW�������%������Ghjj��MMN���3WlZ�G�n����&q�����]]Y���:mq;4�MNL�ɣG�P�y�N���_����S5��u��&#C����M͙�aۖ�X\\͑aii	��ш�V֮7�:�n�a"�+�򽟟����F��ƣz�(����9�����!
�|�b����Ey�WWWG��#����I:|���ct>���E���	�ڃ��/�/`d`H+�Ϗ���}a�����K�a�����|<��q��E����C�*��U__�.����7�����Q�13����)t���M�Ei�ʑ��6mںvSB!�BH����Bk�&,�Ϲ��b��]�9e]�\��ܬ�X�T$�1S�!W���6���?��?�����e�����W����U<�|�S�O�i�E!�s����_�uTB��vu!�J�o��ѕ+Wʪ6����Cg�����83^wX��ElK�f�N����虯�n�l����� b��'�����������^Du�7n��Ӿ��� ���³������[�nͶ��ա���'��m����U�׺\����l��D|
۝m��%�F!*��ԑ7.=�U�q:�?ѿx�U�����֖Ʀ&4�����5�g%��_��&>x��P�QN*�OM����;*�{�ｘ\ ��('4E)x��q�E=�,���D�������x���������GCs�4F{▲����g^�[�N�R>[[D��x}�ucSc�X?��oU�����ٿ�`��u��j�
�T������U�^4�{�8���y^b�������R'��Z�0so�qiQ��wmw�mIT+�I�YC|7��:!�B!��O��}m�0#]�YV7�������k�"5�Xg[k
�8��\h���ɓ8p�@��D�ӢB�R�9G���w=y��E�&�{MOLF�W������,j뢑MLON��i'�@����I������ً���qP(�OO���Q &{���"�?��u�hff&2��(_�����f���龣�WG�ދ��0UQ�ϼ����o�78j��KKi��dD�
G�;u��l�~r�+��mog7ZZZ������{N��G�}��}ٿ�8؋r�z�ˌ�UR7�cV����I�)k��CО[�-�x��$?���/ëػ�Z����ڐ�1�OPْU�$U&�S��:]���V¥����m�ė����s�AT����;�=ë�_�����'himŎ�;��Tn�ra;l���vK��z�f�]���wm�~����Giq���һ�[�����?{z���!l߱��}ss3�������_�ԈH��+LĄ�(����Ć�6DE��H��6��>��Q��"	->�����k��bBUT��$��;��؎;��ц��zt4�ɺ�m����Ԧ�o�7m���� �����Ɔ��;Ա��k5|(��؆�����v�4O@�ZU���d
ɵ�����yU��_�de�(���п
�y]�~]��qpf~��o�xٺ��_g'�����	�2���9U
�	!�B!���:t��d�>����+J��C[�P���a�%����V��K�-ꆿ���\qQ	�L�IT�CAX�]�s��lڲ9���م}�"
��ж�#m�Btv�ȡH�^^\���8v��'����]|6������o��_������NOv�Sؾ)���(_{��������UD��E�xtt�w���~�ܹ3mQ���OL.ؾ}{$�G��������_�/���q�5�߼��	TUW�csD߷��G����pZ����}�5>:�񱱒�CT��B��ؘ�����"�EV6FmP���U/��f�w��f��f�����༐ns��|P���ܾ��S��v�f�ܽ�� O����_G�&�N�>��_~/^� 	���|�����.'[�v�8/a{�5�Nw�_a���=q�?|����	������/`�� zϞ=�A-!��򦩩	5uux��ܵ����ԋU��5���}	�5�T}iƩb�ܛ{�>�$D��֭[%wS�S��:�0Q�:�e.=�tWt����B���d��9vB!�B���X7!�����e��k��TW{�����Zfxe����ʋ���~��߇"�%n��>���A��y�s�\�r_ݹB!�}���o��}����S��qㆴ�k�������s��V�,E��1����h$?���bM��:�d�-I%)��
����$��%���P�Ф����7����˿���X���O?���\�*s������jm����S�i��%q�#g�İl�R���
����ڮ�?4��7o���?�g�B)_~�֛����E۶�Bq�ր���rm�o�!��:��ˏ�}?�5�V024�^�D��˗�u����%���������/nwO@WNZ_���&��6m�1Jq;!�B!$��������0/]J9�Eu���=~mrg��~�������uD��s��u��El۶-�dK§�yN�=���hV�$�ejz�+Kطoz{{A!��9x� ��3�fg@����e����}T�ݻ'O����|�j��14T�y�8����LB��z�]۷�M[�<ŉ?:P�"�ӵ؟JJT��;���0h��q:��?�z��R;5���n�G��|���~���Ɋ��^<a{fO�v�c��vm׋�o�~��_A!�<�p���v#�v�j��-�����#��=�N,]�����ڱ�̠;�LP鎩�"vU��S�nYfp"%�=�dNB!�BH����fg��C��f���E�.�D|��nh��+�������o������I�&��;B����!޾�&������B!�X���#���矢eKq���y�,�DÛo������i��ceƀcP��W��2>�2�2Rr��bm���������k�ASخv���l��s�����V.\��]�088>�}�x����ۛm�k���@��|�����*�X]]EuK+^�u���� �R^lݶ�mx��'�8L�zԮ�b}	�5c�
��k߷��--.��.�QWW��7o%U�u���+D��ڲD���������B!����xI6�+B��6���E�O����X^��KL��=::?���(����՟?��CB)On޾���|BTt=}*c�����;g�e#[�����5��
k��W��{Zȶ ���=D�
�[�05�Y�v?^OT9f|�$�,�KTb�������I�1���+H4|��g����o�um��!�ǵ=ۮ-l��	��.?����m���x{���$N�>��1;;B!偸Ǻv�>��N�!��[>b�ڮ��^�O�(Z�,��$\Μ9����E�$��ߩe������ͱy.Qe��&�Z��0�GB!�B���ë���5Jw�����nuz/h��y�s\j~����իغu+���A�gzj
c##���K ����2���������CB)/Ξ=���aeu����uAQ!j��s�Qj�:}[k�~D����c򹟚������d�uC](p��T�SC6�|38La{ʲ���̑A�~�q�.,�T.I�k׮�����|�M��������H�mO�V�k��+X,��!�S.J �W�w�������Ep�R&���_��?��T���ȧh����+c}	�5c�
�彗D�n�k:?��[�n�����_�eշ�vջ�:s%���}=Q���%������@!�B!NkÅfa�53�rpW�-EtS��^�e}|d�V�1�������?�D��_S�N�t�t���k�Կ	SSS �Rl߾����	JD͓��D�[o��6�3��8��c9J��;�LW9����ִi��Ԯ�B�{�<3p�:���N�LA����vd��m�~0-��/�rJZ勿|�2�mۆ�Q�����;hinɶ���n\O�f��P=�4����u��T�����K ��+����1��w����� �oΜ=����-,J���;b�R��5�AE�J��d}�_�_
a�5��y��@�A$����	��V��eX6KBʺG��Jم�9�v���t�Lb7���Ƶ^�TC!�Bq3W���3c�՟�"w�)�Ic,/�"Tҷ0Ƣ�=:z�07;BT�UC��[x�w�H$@!$��������x��@��ٙ���;�16�r�r�N��>����^3L�h�U��\�а���wo٦�ֵ�yo��!34�ĵ=�XY^�[w:���⬮r)�\�D�awc��r�|��5i�/^�Lݾ}��@��O>�[o���\�e}躶G��36����{��^�����M8w����!�ē={����]�~��-��N\�����Jsm�B�h9y�$����������n����}�� _UM'I%�?�$!�B!DΓ�j�:�����=���Rr��1���Q.B�B�oܸ���v��̀���o���Sl�ĕψq�|��x�W����B!��7������� �<��n)��ҥK�5���߷e|l{ _[W}N���-�6�8�ч�0�6#�8���n�۝��P�9���n��#I�8��ݹ�5i%�U�G���"����Y鸶[�T�sW�D�n1,����u����	�}��NNM���C�@?!�ċ��f�:{_��ƱGo2S.��R���`]a��X��y���KÊ/l�Ŏ���OOr	�(�կ~e{���x�ee�?N��a��%��ֺi様�'�B!���H���F$��������3�R�k\����]���j���؈�7o�?��?@���Y'N�=BT,,.���'8��ݽB!���ի���/XZ抾D���
z�w�D�����$�q���S6�i�wp�isU�>k�ܓI���a��w?P��ˍhO%��\nP5�C+A��潅�^D��7^,7�s�N��΂DC���5]]UE�vG�b�J ���b��n������B��m|��o�νo{��;��G�.?@P��f�����їD�n�_퓇2����oF�V��>v�O��;Q��-Έ)G{�M�0,ն��ۄB!�BPײ���y��mm��J�)˖�TW�W�U���v�a�%���_@�aue��$/C�xi�6�ۿ�== �/<���E��/�?~�D���F����h�홱��9�E�����؆u�mY�ُ1�7�����q8��MU�Y:Eq���r�Z"ws�92����{$��
~��,$!��ӟ�����|�G��\�%vmw��+˵]���}���������?������B)b9���!�v/�!��#���E��+�8ߗ�^Va�G���,��@���ٳسg�g��tfȿ̠�s�}����h�zgj�zc��B!��f,ьF��[���m������].�Uó^hi+c�B�V�߾}�6mJ�I�h[���He�������701>���9B����x��~|��� �1��|�$:�n݊˗/��Ԫ������0Z�����f
ߝ�*���c�?�Ը��*�>�G�����ݛ�8;c������w!>���vdȄٓqKZ+��7ޠ�=b>��c9z4�8�����rm�����@p�:f�?�z9>=�S~�� �-Ǐ���,��MW%����!��*V) n�%"�9qK+��{ih�����<|�	j#��V�;�s��i+t������p�#;�=<C� �7�f����{�^�VK��ƽ�ݍ݉�vbw^̾x���b&B3!͓v�Q�>�eZ�k�&	z$  A�{W�ŭBUefݬʬ����/�jԭy��Js���s�)�d�HK*U�x��!�B!�D�^�6e�H�z㏀k܈�5δ)�R�m-&�1�'7���,�1���C��>����悐H���%�ُ��}�w�$��(iiiرk'N^���D������8ǁ|���4�2o�.@U?����^1���|,�K�W�Ⱥ�Y(pw����/n{ج����e�C_|�"wu�*�Ɛ���'�P=��6`Μ9����0�xX^�ڗ/1g�ܘ��]�M����Ǉk��\�Ip�v-=�=�^X�7�x��� ���EE(�5%e�Z���H��vӱFk���<c�v3�{Y��v#���x���9���}{��i!a�FLL����Jj���dc�IS����I�B!��ȴ�� w^��8����l�K5�W����A���a�%&���g �QQ��wa�u��U�ܽ�_ !�gٷ?.^/�#b�G�C��v�ޭ���6'�#!����7����}?+j���h+�)��)��z��Y(pw�Gi�E�>�c���Y� T��Ǥ��$�$I*' j�|̉X0Q��g��@����;����o���=�M"n���Ʀx�˖B�k{<b����b�Z[�|�
446�it#��X&M���;w�ҵb��>bM�nFDnu�V"��v�ۍ�	�vQp"αc�_��l��xc��n���i�*�2���v�����m$o��aB!�BH4��S���6\�O�5'rW�cy�5ƊD<��֭[1c�<}�����Ԍ���@H$:��PS_�U�V���� ��k׭E��j���h4�֡���9/^�իW;*\7�����:��"R�P=����V}����fL1��y�fL�}yUKF�B�*u�* tO��v�!�U	�U�b����`6~׮]����o*)F�˝��p��1LKV%µ]���wm�k�ŵ=<ބ�τ Oߵ=vQ���*�ݘ�]���<t������!��� �<|�.߼&�>'�>�8a�nl�&nE۩)��4,��v3�CCC���q�<+����is2>�9�f�T�d��2�Q��1����HB!�B�1��fb��|u(�)�b�(�+���C%F���˒��=�>���}����q���rl߷�D���gشn=�͛�/^�BHbBٔ�t<�k01�x�#�r�С�չ��x;]���5�Mj =J��q�F7X?�"j�{T�{�:�T��Xf���!��d����^����Ny���U�N�}j���B'�ڑ�mn�>�+V���r�D�����W���9��=�M"n���#��wm?�!��C�jU�gY�� 1�����<~��N�'���O<G!�~<���]w���X����ܛ���8����}V?��}�arrr|�&�p�j���w�M�,�h�v�k��e���-�`*��S�N!�B1FI� �e�M����\�C�?��?+�*7��K;̚�Xb����T�ėښ�l���) $7�����{|��mmm �����0w�\�^B���܂���d���2�j�ڹܡv���Z&V�q�WeN�4˒k|÷��l<l�s�&_
��v #����-�*JVE�K�G��{Ff�8���}�h>�}�(pw������������E�Y�|_����JodZ'�P�=��F�tc-�l�[v�5�i׼�ux띷}"w&�	!�^v�ٍG5Ot�>"�[�{��3u�Y�����0���KkS�ڱA{Ճ
gٿ���k��?>���KR��c��̩ ��J!�B1�Ǜ�I����d�f8������?Gͱ��3Ɗ���֬Y�%K�����9*�`��� ��._ġ=������!�{�:�G�ӟq����γz�j,_��Q!��}��Ǫ����FK�~�K'��D�pR�,x)n�
��N��姨�۵bwY�<��A��H�j<�1���ѣG��}��\��)����K8z��qm7gBЦ��.�í���b����q�C�h�hÑ#G��矃B�=�]���him�%r�]ۭNr���| �Y�c����(���z������ ��\߆�v��]�n[Ǿ�`eG�� !�B!��ù����3��&�1�7���R�n�^D9���1�[�F������a�?~��׬BNn.��8�]������>�]	!��CZZ��ۋ�Ιz�"���N�*=�Y�1�'��v�e�ƾ�q���h�X���$����I`�06(pw����lޔi��lS�u���4#�d�li���Zwc����&��Ν�6�ڵk ����w�>Lʞ�j��k�,����7k�=6bl�����"� ;v��M� �_���
&M�Cy��`������=ǲ0�L���=��d,�X��	�c�?W�=q�iӦaǎI�l�z�����1���&�F�I�op�m��={R6*�� !�B!�%�#؜y�(�&���ci�o�d�e4> p���7�d$�:����A����p�z1:��'O�BH��I�:{��e�ST�>���IOO��s�U�n&^YT��֬�l�^�m3j����,��vǘ�B���t��#u�%���jS��91Dsc���?��b9�ÇS��0����z�
�8�{�k�,.~��&D�m��H����v�z7�'tlooÌiӱr�J����BH|�>}:�/^�;�K|�������o�F��ٯ7�,K�v˓��$J����sb �r��1ddd_�A�K��c�*6�I*�x���fܭ��Ҹ0�e3
f�[Oq;!�B!�m}#ȟY���Ni�P6&��C�X�E��z�@���y�E���F�\�t)V�^��w�8Ǔ�GX�j%2��@�zzzp���m߆�+� �_�a坲���
���x��	��l޼�gώ����p�5Cm�r�^�6�6b�fl��o��"��Q�+�;LIS
֤Jfo踸�;a��B;1xn n�|N2�1Ĳ!p���'tR��(�??��۷#''�� ���!�iwm�d"�x�}����D�eA�M�{�n�6�*���	K_]�;kjj@!��yyشu.߸�{����?҂0�L���=����cEK��g �"��9�����h�7��D%�Bz��Q-�P�^�:$
Q����0���lp�AB!�BH,��OW���:bw�R顱����^�Okw��.#-��X%%%��$�exh���ƺ5 �(ͭ���?k׭��;w@!$>lظO^֠�����q�#����=�z�pݙZ�dRw�=�,�dq=c,��#�!v"�G��B����wy�}�d���9�EZrP{�Dr����KB$֍��DVnn.8�O>��9���q�����.����n�/c���gM�k�� ^��a���>y
mmm ����8p� .]/��`��}���/�"�޳L	����k�o@Ow7���Y�+V��K����H���m�)$j(��*!�HH�r[����sa��aޭg��B!�[S�T��+?G�zC.��0gw��X^�9�w�cEBoǏ�w��]�#4q�G+���אEwb��Ϟb��7�l�2TUU�B�5�����A<}N�#b���A�|��Y


|�H��zN�e����za�M9��d���7깷��}yW}��.��=#��E�a'���=�8/uc�$���~'����᷿���c$����Sضc������V\��qtm7ؽ�X3�?KBAo��*V�����>CGG!��#--��A���Ȅ����X���k�õ��q�χ�.B�+V����	��h�����>��M��
�V|w�%�����~Λ:��B!�Bb��u���ahpP:�Э#*k���X��|�L$�R4�l�<y2��ۇO?��9����X�v51ý�R�ش��ݨ��!��ؘ�`>�f���;7A�Y�^��{���&M
�v���>���s���wc�B�����xQ��
�]��L�1�� u��;1h��nwc�s�7oƒ%KP]]��=��z�
����{�W��k�_-�nr�k�?Ԙ�ݺ�0��?�q: ;��ϟ���c��>�%�!�CL�<r�(n������$"Q�k�p3�^��Y�I/��L3�q̿|V��.��_���q��!G\ⱏX��$�cb�CȉA�Z�4I%�{��e	!�B!V�)�H�tըH.��0w�)�̓��^n���)xx�P�j�u��A
�]@��]�<I�.߸�};v�r6� �b�3f`��E�2z=%�,�}}h��q1�uC��bm�5>�0����y�D���K5��[�m8�������a,����aT�\B]�@����
f�!~��Ē��YN~��➥qq�cݵݪ�ݲ�\1#,�o���=�|�u��4'�/!r띷�O~���^B��o��'p�����5�&�>b|��X���@��p�/qQ|/,%I��Jt��?�?�T����f��B�v����&N� �B!�X��/EQ�H���jbn`,6�	�uV~��'�1֎;�`�<��9��|.YB�r��>���!����B�1�M��U�����AH,<,-�{�x�W�n�:�E���G<�5�Wcmх�����h�KV7�����އ@b�w���gLG_k��ҥG����$V����7'���}�{q��{1��ߧyG_�K]�#�=�?y�a�����u���c�x�M��w���� !�����>|w����G�n��#ք�fb훸eQp/uV�nf�/�>GG[;222@�C��B�n&�H�����S��L�J����x�"����=/� u/�� !�B!�%u�845͜)�v<3��F'�P��l�e6�ic���4_�����>��T=x�e+�#�.�$�_��;��z�Utvv�BHd�L�����Q�NbF��?��FF:%�Ns��	��-L�b_�YG��S�z�\?Ԏ���\]w����t��S�j^M\B��$LI*�L���.�7e���n��G<Y��s�b���x�"�����slݱ�Yِ���F]�ÿá��c��ܲ��&��8pm��3����A'��!΄#���GœG���R�Z����d'3A3"r�����'����`Μ9�����S�$��D���&vW����\F4c���"D��B!�B�!�F��)����lX�*Əh�����,3�R�b7�J�(�f�������~���.�Utq'1"��/._���{q��	3z!� ??��n��ۉ*J�3<L���dff�СCq���p�j��6��=l�x�`�P�f�j7P7̙:�&��«�K��rG
�ͻ1��F�n��T2�����#��D��}9r�w ��.\����7[��ь�{��%����>�X˂6;��E���_(��^���o��6~��o��&�����h��P�&�>�lTn&־�[�?~��f�����>�v�<!]�,��6�x6��2�����ɕ�k�����t�U����L'B!�B�u���=Ҡr��C"�%K�kW�JM5n�����i�������vK�,��͛Q\\�,B���k�"3+��E\��~yGĹ3g���B!j&M���w�ԅ/b�"��+�@�g׮]�={v�'��ݧR���Z[�Yo���=��ڃ��9`��:����0�`:zۛ�UV�Ė�j܍A��/N$����;�����A���>����|�D��܍ݨk{�
~l�[��$�wܵ]�5~�fD�C�x�X������o@!���;��--c-�����eYDn��e�����In���@�;�н��eӏ;f)�V�v�x�b3���%�ԛ7�jZ'���$wt�R��I*B!�BH|�Y7�]�)���?�OQ,�_c,_@�^	���=��N������V�_BbA\7??w�����@!�Ovv6:��ϟ�=?+�%�i>�Ę��ѣam��cmsbZ���u
ջs���5C��g1��vχx@�����E��^Z,��Eqc�o���ɛ��S^3�ѝ�H�X�����/~�؉��	!������$F���O~�W������>&O���P[G��e���g0'�3AA[ͳ�x�|������Y�������756���I���Ϫ=�����:;;���S8�p�ɲ��>G��]U�H0���I��Ku�p�;ݿpA����mN��g�ZWW���w���n��_<kh�;w.N�>���n���L%ikknAEY�$��5Ȉ�|hh�����}Í������*M���������6<�|d|��M�ZZ}c���\�k�}�aY9i�k�S�ց��B��-\�0b�[� ��>B9)�#c&Q5���DLR�%��\<���B!�B�E����NGog�����M��#c�~
c2��ݯ���?�3���@�%��>)'�Ă�}q�<�3�N�B�_����~����cuM2>�����G�A�gƌ>�d���ǘ�v�x�`�Pk���F7�R��s���@�3���.�F�0�MN�]�<Qnj9��DKq��B<����7�|?�яl�U�����8%v����I�����~�k(�2E�.���/���g~���@�x��x���A����Bܾ{�^��5]#�Bܾs�n��j�k�����.^����	v���:�����N�BS!v�9s&�����X�`�B��-Z�H�����m�ԩ����gw����&���ů����.�5�7o�#����aڴia�۝�����������U�����"��r��@OW�o2��ysUǤs��&Y�qq�㇕X�|Y�8�n�=ߚy~\Q�E˖�}�ZĽ�l����z��7�|=88'�'�o��_�ͅ{��-R|<���86��KT��+]�ck]a�d���]�WX  �B!�ďo>2=M�b������*V���b%&�[1�
_E�}�V��ǤI���[o�׿�5�D�E�NM�w�K����6�G.�~��Ήk�=]����Bz�3����v<��v�o�����C_�#�;�مA���|u;�͙�ǌ��D7g�`��N~vq��ߩ�8�D�fE���ɿ}�ϩ��g�E-�����}δOC��N��ă�0�r'?{�������@<�4�N�1���8u�{��T���T�eJ�kH
kn�g���rc,��WR7l����.��;�;u:��[�&�B'�|v��p/��Tcn)c'����b�,I(��b�m۶�ҥK �"�O~v�'r�㕈\�nx�b-��M�����-�M<D��_7&�[p��ߏ��|��������'>%���Ğ�{Q�܈��F$�>bM�n4־�H���f9v��#�T��J�N�c֬Yؽ{wB�Opy�"1h����OTI\%����1�x�����Z&�!�B!��v�5�q��fp�S;�[5�R�����D0�:q�>��c[�s�D��Dw��n�8@��\���'ǭ����ȟR0:�wȨ��ڰaE���G[Kf)�B���=-3�֯GZjjPl�H��)��D1�͙����3hr�͙�9՜9�(d��/_��ٲՇ��{q���O��H���.����/�c��E�'���-�H��Lu�z��gOd�BH��uճ�0��/�Vp�K����}��~�1V���s�=�w.T3T�Q��1�2c�%3��w�>���
�]F�'�<���'�70{D2�Ŀpc��%n�#ل���w
��A�����0s��O�H�����kT�gYDnB�������Po��E�v������x��i��W>� ���7�$�!$шg�����Z�Z�1V'3���X[�#���m����H�W�> q��+]��7�|T@خ}#4&6����0�N4׌ս9�@!�B!�σ��������A4Escu�ݱ��v��}�c-[�7nĵk�@�E|��K�cˮ �
���y����|q�#4Bq
1�c��=8y���Pz�$.5Hba�5��q�ڳ>��-��c������H�ʺ��u���i�9/(pw�j�ؙݍ!|�A���	-Q�h���<�"�1�p����}�۷s����"%�"�ϟ�G|���"������n��ܲ���=]�#�
��Gϟ��w��~�{��;!��W���#ǎ���J�����o��C�v�N��Tzx��Q71B�0?~ܶD�'\*7A��U�1��2�è�K����B!�:S� ���0�
M�U��KV��#�B�X��"�����
c,
��A͓gX��uL)�
B� ���;��{����/���B����cۮ8}񼭫Ӑ�CKc�^P[��F��mf�k[<�kfjC�P�ި�=d�%[���0��z��n�Q��=y`�0~P��2�G�7w:�:[�KHg�x�Dd'�4Y�I��<��#���}lB,"�U����@��֍�س-^�x���k<֨�]���U���vƙ��*�4k�%�?�����?2aE��g��G��~E9:���޷�>a�n�ν���ͪ�^'�i�z<��}�}x����I���͋�f���LK�GNRi7�n�J6F��3	����Ƽ=!�B!�D�f��2�jW8��]5~�*�6c�hE~c� ���1����x��СC��w����z�)�[������k���p`�\�r ����ԩS�e�6��������xp�v	�;5�]�v9^L�˻�
}�f�*ǵͱ�c��� n��O(pw!m��O��.�r����'�dN�D�:��U]D����h����\��%|�_�?��'��݌��M��M��]۽�8����nQ�nU�3� ��{����'x�����Ą!d\!���@ɃR�h�V�zIv�v�����Ǔk{�����3���n@�W�;�fv��ٽ_�{����х�z�*��^�|<e�A�Cj��}Q�N!�B�����/,B_wG�^u�g��MV�OM�P3��� l�ceff��Eݐ8O݋Z4��c��Y �*�y��8�{/n_����fB�x���k7����gm������5hnlqo��6��CR�d�Z96�dm��@�z��,���Z]7ND�����	��wr�ދ�Y��=�|�"x��$��41#t�_(�N��O�$�Ѿ�Ν�={��̙3 ����c�޻�UkV�^�um���ܲ��h_&�tm������̇�U8|�(Μ<���6BH�#�m+W�����>�{�#��!a�{��i������6���,\�;w�t<�����;�skfPjQڄ�j�\fp,6�2��Nè��핓�	!�B!�ѝ^ xZC�Bc,�8�;6�78�	:�k7��ϒz!����X?��}���)�y�<fZ�C�q}<}��n߉���h�X�2�����kW�&�/Ľ���� �@h�1V�k~n]��?F7Y�ea� K��sPgn�%�`��|>��m���������>�f���=����y��jڵ'�p�Ԟ�A�g0����,nLB�9^��:{�3��o~�+�����sF�&D�m6	�-����(t�*�7k������I5>��KW���KBH������������g�DVV��ݾ�����5'��X����:+X����[|&v!---���.�ݯ�$KBA?I��믄a�A�ds�2�YY�(m���B!�b/��S�.-4>���YR]1�״)�F�>���-Z�l~��y��hk���O�p�����>�{z�C��ւB���3�\x��2�'�+����<�9s�D��K�ﾌ�{��G0�VL�����by|����zz���ݥ��NA��Ew�G��tI�~1��+^+/����$�ō�-I(3���%K�����yZ�[p���ڳG�M"r��6���{\���&�k��}���'��q�fL��B��RBH�1}�tlܲ�����s�(X�	��X;~�X;D�n�|K6е�-��������`u�������n<Q%GZf0l�-sb�oƔY�42QE!�B�������K5>��_���Һ�̥��XƏ���ޢ��Eܿ]�� =��?�_��m7#7/U�U ��de��#� G�k��-!�bhp���jS�6���g[<���pիmP��c���jc,o�q��n�?�mOG@�G{.�����A�l��B����8�\VA��6Y%�I��%�G_a��I(#m����{����m��᷿������h5#"7kB�'�n�#X��+ݣU�[��b�~O�?��EQ0� �/s3!$yX�t)�,[��7�����9f]���l�-�,
�a����"n�������(,,�N��]����*�P��u�J_�.KRyu��a��&����Q�)Vʠ�;!�B!�~z2��v����Fc,+�ݽ{�����ӧ ���ׇʲx}�*O�o^����M[6�Ƶ� ��dc�ƍ���͒; $ޔ��bp` ����زe���D�C�S�G^�Y� +�S�Q����q;�q�w��50�ܹ3��������_^=5���C���\\���$2	e�~�ڄ;�~�����8O_?N�:�w�v���0'h3#�7�=��{]�-�e�g�����ô�"���[�㧟rb!���Y�ٹ9�~�V�ͨ���}Ą`�L�����{���!����_��a{ .1�.��DL�5ow�]��:	j�T��������^�8Z7IHP)��9��(��r8!�B!��ō:`c�W�����>''�]���4�fcb\���|�T��c�+K1)7�ē҇�X89�M�fHI�s˶;PS�5�/AH����FuE%�{��W�6�X��5?{D�!�,���ߩ=\'nY�&l���7j= �w�8��O����_|?��N�HM�8����)^���T��3����D�{����<ߒ�?��A���3g�}�v̘1C�nYDnP�����x_�tm�EDn���ٵ]Fsk�s����C���;�B�Ȗ�[�34���I��#���'�eJp/�G��6q��� ���;v`Ŋ�LDّ�
806u�1�иX�̠�Z+
�h&������ENCB!�B���;�ɋ����]��.��V~��yB�T�X�7FSN2�1����w���Cttt�8���������[AH�yV��=�8v�8N�<Ś!!��ddd`߁��q����A�ܿu�7V �@��,V~o�W�⵲V��������(3���L�u'�KVV�+���j�ws�փ����ur����OXɜ��5#��&��PF�I�v���~�A�K�����_����#�fYDnY�����{]ۥ�1�#��u����C���W?���)��\Kq�Q���C�z�-�-�6{�#��D�v�G����:\���.��� �;����1����!a{�g���e���#��x����=c�8>$�B!�$�o2=-Q��'�j�򕮴�v��Ke�%q��7Oc���|������A����'X��2N+!񦥵�/���c8w�,zzz@!n#77����]����A�4����������#''��Q"�����ۯL�ѸeE�!���F��ZS��Yu��~h2X7�
�]����Sg���>b�J���'���a�����8�zÖ�H�$�D����o�>�:u
�<,����X���w����ƃk{X�)�[���iFh�?�wE>��	���@!N������.-AOo������{�(����#Bw�����OU����K�b���I��2ۗ@��
��D��I߽=4��q�,c+&���
����I*B!�BHb�V;��y)a�LE3����+]	S�ڡ�M�E��<����������A�G�ݹv��1=�#����/N�о}�}�Y3$����ӧc͆u8u��y�;ㄒ��A�Cvv�ou)N��}Lr$ZW��C��[��Ħ�𦥥�z-�vA���y�7	Eڂ�$Aeĝ����I��Q&q��dIBY�_�N�>�Pa�̯~�,��ː���h5!"�,h3ڗ5�^,]ۍ��*���
l߹�e��� !�8�̙3�q�f߼���g?����k�E��)���XcǤ;�\�ܽ~�Ͻ.C�*%���̉(#}�Ƨ�ve�JyA���uAol�ua��2�G!�B!��3�E�ԙ�io
��[�9��;��"#�/^�={���ٳ �����% ����乳صe;�rs���cB�ӈg������� �N�+*����:�9s�8^�K���\���\+��:4.�7�RQ+4�J��I��0�b���;���%-�k����w��ܣ%�����;Q��x�NBE�j_[�l��5kp��]w��ڊ���Б#0-"�$n�&X��ںQD�V����x�={���,��чC����hV�\��sg��kWl��X��3u\��Y^M��'��cǋ��i�c476�����;v̱���ɱ`ZJ-l�:Q��k��v���ݣ3�\=��nc�h�t�!�B!�$���y���'=]];4,r���2�:�{���z!��Bm���.����p>222@��k�ū����X7u
�ܢ�-!�96oٌ�����b'��(�{�=����h�dqf�kw�����M!n�]��v�&�����b{֗3�+��w��=�2
f���eXaݣsb	W?�C]��#:1(^+/�����b䶄S�m������?���QTT�j7%��E����`݌ͭ"r{�����g��x����yy��W?���)���@!v#��v�ٍ��N�,�c�c�>���wjJDn��-3�e��!Bw��]044��;% ������ɓ���$t�ǅAo�_^0R�J������T��&Q�?u�R�N!�Bq�/�p�0#�=NwL��*ꆱc�j���Ac�H$��=Rێ;|�eee �  �Z�i=��;��0w�<|��~��BH����ۇ��>!v#&��!q6l��u�\&>�_���S�5\�e�ʺ�n�Pn�5�̬,ܩD`lL��I@EG&�y�GO��,c�Ɛ�
$�:��׏�,3�&{�6����uuu �@<D}�?�����l�~�,ڌ�]��n&�k���ѵ��n�а��=��8�֛�|�2�jkA!v�������Ni	�::u���V��-��V���#�c�*�wZ�]P^r}����&D�Z�e�I��D�ڳ9 nW)��^mJ#b�}DW"KT��v�N��	!�B!N14dO����z���Rǹ�t��HĦ�b6Ƃ�f�+�E�ь��x�wwQ]Q�E˖�`�b'/�j��юc'��ʥ�hmm!���ԩS�e�6\�z��|$!����Y�w���������g��иT�0 n����uEO��u`��B��]8�F����$��q���axpP:$�r��U�%!qf�z�'��Z�$��"�Hm����dտ�˿����wKP��._.0(h���n&֭"r�5a�u�'�mW\oVWa�����b&�ܾB�7���Ǫ��q��˄�V�#�'~Y�'�e0N/v����l�@��Jwq��!��&�M&�H�{ ���:7�cTqr14N��kU�uΞ��B!��7�=ãc�C�X�՟哂�b��i�u��q|�{�CSS�;��;Wob�у �nz{{�ǳ��e�F�44���
�b+V��܅�q��Y��Idb �gw�����e,X� ���O��_|�
d����B��x��[h��0*��G��+�	�I�H�tx����$Kss����. ���6�̠�cPaJ�'���}��_��������|�����_��A,ڌ��ڮ�}�D�H������>m9�3�O�����o؀Iy9�t�N�U�E���8�f�\ۍ��t6��nHݾz��3�!�_�����dqF�b�?�m�ra���"'�d	�@�*�p��!�B!�8˝�A�3k����-����X�6co�����'���+�{hnlD͓g��x!�q=�z�V��;v�ĕ˗]��%��ĳ��m���݁3σ�D���- ���?DzzH��&�{��d�uC�M-n�b�*�Fwo�7�
bi&�O��Ei��vC�{�PҒ��F<a'ˈ���������� �r�^��()1h&RR�/b��VPP�w�y?��A�CkK+Ξ9�c'N�tm�V�C���#p��ܪP�L_��S/��Ѹ��fL���WG ���?����+b �w�>�l�CՃ��s"�k���_�E䉼g�ӋuZ��b���Ghn�ۘ�عs'V�\�x�I�����jq{a����D�J9�V%���8\0z� �B!�'�򔼙�4ר풉�ac��B~d�h�X�#S�<���~򓟰>�2Jn�¬�����	B���
L/���o����g���B���L'j�7��AKk+I�}���.��(**��o��*��5G�bӠ�*k�Z��Y�v�)�:�Rڔ� �C�{��m����S��nԉA~�z��jf�A�����῀(�S\�p����׾�5�����e���$V�]��s愽g\�f\<h�>�"rsBI#���M�k�n1�3��ׇ�G8t�0J��Gee%!�,�f���-�p��m�Ȟ/��Gd����b�pm�߅��J�v?(�S�.ĸ㣏>
k��9�	;]��*�vu�*z�J�ܮ�T�������B!�B����t,Q
�u�a���f��]%nW���| ֕�RR�/b��6e����������e�)��-�@H��Xg����޹y��� ��X�3w.V�zg/]��0s�$��ɂC�� �BL�����vS������B�H�uB���R�Ľ}dă��i�={@��$�=m*�=m:'Md���M���*��ܕG漰�,V��={6�?����7 �A|������_����k3'h�C��V����wZh��߽�Ǐ0o�"��lN~���zL!FX�a��B�ɻV�#&��c���g���uZ��a{���o�D��]�Y�[�nE�8KDYuaP�ݵB�p7�do�I+ɘ;�p6�A!�B!��Q�kLEO��K�V(_�9��]��]�f�ө�j�,7�#�Y!0A�W����\Ɠ�GX�x�fL!�b`p 'ϟ��u�`�ܼy�b�l�i�f�>O��x�$���:�<y�.rss����#%e|�ڍcƠ���b�L��;�G2�ҚQ�O��gO�K�'�/F�'/E�̠�Q.������BȍAv���Ag�1*�3�L.9��.����1̙����ӧ�y�:�l��Z�v+�v��:�	����õ�(VcM�������|_^����zB��y�سw/TW���$ª�ܠ0�L��ޖ��E���+W�G����5O���1�Њ�$c�����̱�0�O��{,5(OT��#{�g��!�B!�;�)��$]�Z�W]3��*q�3o�%�xʜ�̗,��xc=z���oA܃���}��8꫃�H�߹���g���c��aOO!$y��]�UZ��f:���#�w�qr�y�w0mڴ����b� ˨�=��9�{u�J��l�g��VL���IDϠ�
g���^:3DZ�OKsn�w��KR��D�(��jwu�j<��#�-[����ǩS�@��'��5��X���U�Dqm׏�*�4�+y�D�N����(�|��֣��/^!�hY�|9�,{Wnݐ��`�>�3���NM��w����>�$�y��� ��W^�5ܓ8���=.���.pa�*I��P��_��/(n'�B!����^��AX�=�)�gtKS��,Ky��*1�(�!c,_%1�'�1֧�~Jc,���֎��X��� $�445����m�&�44��� �=����-�]7�Z<q��J����.233�կ~U����2��ޮ�!d��F�*Ǹ���X�U�[jj
�׺��?^��=�x�3	3��qcО�"i����|/��.]zP�:D
��qɐp�������Ӯ,Md��������ڨ��+m5g.6a��^㟕���c�}�׾@���x�+��_�]BFIOO��{��ՁKׯJ"��G
���&�>bQp�����(/����Nw!��(����j�ō϶`jʰ�]-r�sb��̠*Q�k�d	G�B!�B����"w�,��5�L�t��v�1���?&x_+� +P;L�G`�4Ǣ1���bϞ=8{�,��9�� /?�$q���W�,ŁCq��yB�Qغmj�p��y����,�d,7"V�Z�p!R\^���z!��+��������^2��G+L�m ���u�DA�{�q�n������`����L��=�DMU�R	&���v��]y���q��h0�%����_�[�nEqq1���u�&�oڈ�sd�.Xw��܍�{��;-44��>����щήnlݱ7�]�s!�Y�fa�捸y�.z��4�Z��X�����>bQp/u�}��*&�܉�V�8qnOR%ąA!n&�"�۵n��=����6Q%^�}\�!�B!������(R
�5�X�L�B����J�fGc,sm}����W�&"�\�s�v�B���q5j�j���A�=u-�� ��ٳgc�����������ϯ��������HKKsĽ�i�{�`�P�!�]=���y=��a+>k�uO���DA�{24i<��ԅw:��6z�S��cnju�*��+�,�"%%�NVڄ��իW��r!?��O�������3�bM�l&�����E�����~ݚ�эn��L���g/j�_P��[���3!d� ���m�oz*.^�M��*"�����5�v�2x z�f7�G܂�7ݸ|�I*�"�����׉H 9���B{�
���#v�NbJ7Y5�^^��V�\!�B!���[�CxgV���B�B��\4�{�A�ܹ��X��6l؀͛7�ڵk �O=ƢW������é�_`ڴ"̜1uuu��#B�C<7�۰i�8y����y��-M�|�F�*Q+W�tA-Ͼ6-�1�N�*Ff�5���>�[[7�5���srsq�nJ�,�
ܓ�[�X�ꑞDF��*���RS� xe	+�ɪNb��$g�hۮ]��v�Zܹs�]tuv����~�#����(��(׏�*�4g&VGi�H�v�ۧ��]�mj���D�Ç(/+!d�3{�lظ%�eh��м�ዛ��`�����@�^_�"�:)nO���������V�1m�4�����9 ��;����1�9��O ,Y�NP��T�x��)y�J5�k���<��!�B!č�:�7w<-�U�QE2����M��KE�ʣ�8�B�1���ד"G4�(�y3��¤�1!���I5�L���Ǐ�ڕb����2q(**¦�[p��6ZX�!.���ew1��Di�dq�-d�eDܮ�#�̟euC��6l��6�L�z���$��˃������=l�H�tr��	���0�wJHuLX�/.�3��III��S�m��o~�����W�`���X��rU�U��u�]�qfbM���n<6>!�o���
3f��{�_��S��=:X ��?����];����W�H"��G
���&�>bQp/�ݕ����щ���d�V����#///�:Q�[���GPЮ�h�*܅!���ޘY���2��p�Xy�.�B!��r�)+��|�l<$��׮�po7c���Lc�`�pX\�f�޽�.�q���ؿ�8M{{�ϵy�u�N���K���&!����͛����;����D&���cxh�}�U�7n��"���m�q%$��fo�ڡ|�T7���s�(K�jo6���$qP���4x� ��<z����KT�%���w�M<X��*g���X�7��T��$g�h�޽{�~�z�ɪ��U����ɾ����?���dggc����&��ScF�,i5(�.�}�}�b�pmׂ��^C}�[/������4CǪG�BC�g�}��8�&7����{���1=�y�������A������>4����N���=d:��D�ۋ��w�'?�ܹs�_0eU���^w,^[}oD|�~�G��zrL�"�'3��x|�|˂{���H��Y�C����^�v1���;y�{��\sF���嫾���YL�Ϸ����|�AR���+���x�0xF�v�dU`l�5e6<��B!�B�͋�al]8}�ac�Hc�HYF����BE�04�U&�1����K<��,!N#�7��F����� ���������B>v�n�D[G;q��h��qb\�o}+�M7�ڼ�-$nW*��Q��d�MS/��#�b��?�O���'�'
ܓ���L������4�D���:2DXrP�.�I#P��ĻM�ɪo|�����D��p��X�����I����_��~��_a՚5h[⩽�c�]�BCsar�_cC#���W4Y���s>�&�(�_}�&�F���C_���Ի5�_3����f<,`h���f*�;�|b_%��1);3f�D��G�������a���)�K�S�&�����	Ŀ�D�ۋ�wuu9ҿ�]|�E��e}?~�i3fh"L\Ǥ��~����������1ԻQ��{fwW7�^�F�ܙ��V��������z75�J�w���A��I�^q��_ i�o@��uю簀��)��8��dF��G�½=???�z<��cuaк�k���y�0q���0�f�]K!�B!�5e
2=��q͈'�_Q�
�+��cj��zZ@�~�n��ٶo�>������a�W��\��_[�I$⻘�����Cff&2�2�������K̩��յ65;ҷ0g���v�'?������ ��.��I�c,�� s��CYi��n�f�:V3w'����)����S�]|n'��-��N���N|ޙ�f���?�����z�"����;��u�H������<������N��N>ߊgz����/�v7mڄ����ihk���HY���u@U=�#��j��U�Eݰ~� �&
ܓ�!�Sfb��VZ��s�S%�Kj��nR�;��ɇ�9�M��G��x��/]���݋ڿ����i��x��C'It��e�{`?fΜ�{�p�"X6�b����q�f�XSn���vE��7o��˲k{�����X�h!�Ƅ[�:��;8���nX5N�l-�����X��5�~�5dێ���_8w>�I+��y���)D�ĩ�����z�ԩ����gw����&��� 77ב���W��/]��[70���",ze�"��}D��:q�l���T��
潦�C�8q���xa�����X�u\$j��;0s����K�DQh΂�p
���E��uut���b�@�ĳ����IN ��k�X"�/**»�;!D��mr�2{h���'����n�:��'NC�S&�!�B!���쟜�.�덁d��ʓ���ͱ�c!4nK�1�Q�0����QRRb���b'p�o'��K�V�j�:ߪ���af!�"55ͱ���=-}b~v���v���E}����i�V4���EM�-����+8�����E.۩��^g���2�q�ϙ;��ǵ���ى�ӊ��{���D6��n�\�T�n��G�ו�ܷ��W8��}������ʱUJJ2��bkS�P��Ɵ��a�X^hM�e��X�U���6=�^�n��'1�Z��J���*wo�IpcP^ �\��v�z�.�nqO�c����g�g>7�Xl�^~��?�G��3_b������L��Gp5֦�jE<hW�����YEL��'���ǻￇ[7n�ٳg �����BlݶO^<Å�˒�����ucm���\�����	���ĳ����:}�


��'B�J�_m�%#�0����ܽ=����PlM��x�B!�B���a`R�l���E�J�4�X�X��5�Dc�KoGmr���X�r%�޽k�����@��8�w@ ����
��.Ƥ�I���C�CF-�Uu�8�@_?������t��<�^�U�cŲ�غu+.^�w�q�b=y�d8������0fMN��g�Y����_��,V0u��9�{����[P�Ԉ��!=+٣my��������t�ã�����	�����ֽ�<��F}����V�x�v�=_�����m`B����s��͛�����o�&l��K5cY=c��cfM1�h.�[�aBC�{S�:�����6sDof�Ȉ��.�!U�Ơ��f����2��҃���-vɪ5k�JV����щ+/a���v���Ċ�-
%%����֦3�N����	֍��r�]�](�|�ů��UkV�����܄�!�;v�@Jz.߼��9o�>bP�mUDnq2�~l������du�n���R�6���1Q���ߟ���^Ŧ@������ubso�_�L������B!�B��Ҏl,��)�cV~3��q��1��6����׾�sqO֜�x�v�u�߲	���Ux��)��ځ��V����B܍xذqr��q��u�ĵ�D����n�q/v���k?���ǔjc�`;�S#��)�>c,Ot��h5Ļ͙�GAw'��=�iB!�=m�Y##U�qii~��r��W�Ƞ��KP�(]��	�ɽ�*;X"(���r/�X�t1.^�{m\�,�]ۍ�o攰Ghh��5���j�}�����a���ϝ� �� ���׮��ٳp����$Q�Ms���u3���gY����d}�kkiEEi9�{㇩S�_O�v%�a�D��P�,I%OV�h�T�IޢM6N��܇�U8�.�B!�����i����KU7�3�
��\��c�Tc��v��A���?���L܇��<yT����A����_bƴ�8r�*<���O@q.����v�=4��p����z��U�O\�ƍ�}��q)j�ަ6����m�0�s�Dm�f���N
��O.,'�;�I��a��)]R]�D��=#�H�%�RG�Ґ�ٍ!,qHP��B�<�@'9�U�L`�d���d��9��[�S�H�u��<��{3��pm7J"ŋ���b���E\k+?BvV�|�-�|�ׯ]!�9DrJ�ۅsJ��:QV�#�����w1.X7k��j|B�D�{��q��˾{
q'B���$q�)����R��Lܮ��
�޵������� ^2VV���vK��@!�BIFZS
��i������\�}uDci��������!i�K����<y��o�!n���	��;�W_Y��Ǐ�Zq1���@q���l޺/�kq��9�v�)VSC#�;c�?��?��V,��D[�f��B��@c����f�W}����"9�k��aTƺ�SP���� ��ga��f�J�
ڥ��90|'pj��؄�])lW%�?�x�2'�V}�))�#v��wĤ�o~�����{w280�_����O���(n�n��Qpo�7������X{>��(���e�1etp��{����[���!$q��Ԧ-���َW/���"ߟ]���$�>b���b�xI&Jn�Awg�{E�)�I�ͽ=� ��ݱ=��gD#^� ��}t+(��gta �B!�$)�^xpdj�aS��C�HZ��+m�}/���$v?t�~򓟠��ĝ<,}����a��f*U���jlX���Y�Z\L^B"337m}�J���i4D����6��Ь��lذ۶m����6�b��$j �K^?Ԏc�v�J�Q��cY��8��uC'��}p�1�R�'�T�|!l�.3>���M[nP����]x���0^I�8MV	w�d�͛7A�I僇�z��vlGB]�-�!�7�k�^�9���X[��h��@���ڪ�X�f.^���.�	�������� -7���v�;���nE�nQ�oJp/s�}$�h����*�2c�|��I�|�2�`{�}E�JW��˪6�z��h�v�6��b���B!���dpH�2-/#�ڕ㣴�13��1V�+�1�J�.�zi�%����o������K�����ߋ7#��7��ANNv�ۋ��6ܺu+��ل$��j�*M���wn����$����bN�p1�����Ͱ�TW4ڦ���	M�0�qU�֯*��ca#���0�
�c�	�A(p�vc����l3��.��������P@W�.���$�HII�dU,�/~K�p0�n~��O�ʲW0}��`�;D�	�K�Z��vut�H�k{��Ok����{�CO._�ā3!q&==��؞_0%奾s���ĺ�[8&��7q��}��n��$��y�*�������k7$��a��L܎��֍Aw���pQ{$�B�{�Yٸ�bJ�!�B!�$��2�W1މ0�W�b�f�Km�%��+���X����5�@H2��ۋ/.]��Y�q��Q��/�
Є���ŋ���[v����d����hkq/;w����S�f �NUU/���V}6�ޮ��5	y��9(p'�����M>A�'w�̔��7-$r�:1h��&�$ɪP�&$�NII�dU��۷o�m�/_q'bɶ������w�Y��.�[J���`��X78���%�:�o,��1i��E����:^�
��{p?<�����E
�	���<�n�:L�9����QE���H��b(6A�,��6��G�!n���=��,\����+�O����\����bw��zS/3�	�q=х���[�y�4��� !�B!d��݃M�����ݔ1�����Jc,=���X���c�X���h��r��}֜�(�>�$��u�mū�qh��(�w��� �ď���c�����EN]��$�u�x��Ľ��poW2Q��k������aX�F�nt���E3��1��NC��8���a�5+�C��ɪ���tq���a"��;C��]�'�+�N~qJI��*�HV]�z���&���'��޻a�%��\*��Kpo����=�v�;c-�<�`��ء�!<z���w� ��|B���~B�#�߫׬���p�A*�?�[� �X���G�������H�RU�u/^��q��������lU���D�%>a�Ulc��["�ܮ��
X��#rU��p��]8:�hːs�F!�BI~�S��i���@Q�c�4��=c,��n�cź�-[�����r��K8��qdff��d�Ae�o{u�+8�~J��E�K�	���ٳ�z�4�4���s $�>߸\<�j��C�a�ڵIch����Q����]o�g#��hbv�6<:��(=�ag��}��=a=���iyfj���+_�A/9�"��.�ިX%�!Y%n>��S�@�˗�/`٫˰b�J�k���5��5Ｘ�a�-V�W#�|��B�~� �zzp��e_;!D߽z�:,X���Kq񪿸�k���ݢ^�����c��@?����K��ĉ��۹�p�v٦��$���1���fUy�3QGB!�B�8��fǦeE_�Yf����3��h�5����ŭ�kضgIF*���q5^u9�X��ܺ���&B�3s�L�Z�Mm�>a�x�#��W}v?>c,%�ahe�-D�KV3��N�Y�ꘞ1�Q�vaTv�Vh��k]�=P�>��Z��^��*�I�����'�ҍA�Ȑ���C���_��z�>Q��dIV��_�%Ο?���A�����	���?(�2%�M�D�Ƅ��q�5k⳺�m׺(U/���E�,nPݟT��N��&:;;�克 ����o��������.����^�b��ڮmM�k���v�`7���d@�"��y�s�&�����}ɪ ��۹��m^�B&`�sc����핊�#�6¶����@>��@!�B/� ��gc��ቿҚ!��h�5y��O���x�R����OY�C�WV`Պױn�zܾy��� �������Qn�g��Sd��M�Ҿ��eY�,;�c���q��/���؎�؝8��L���d��93���{���Ξt:�N:��vbY��K�}-IU*�JU��J��\.?�  � ����"���G�x����� 9���b�����D��+ݽ��<���X�z�Gk�ۥEvn�3�Ҋ�C)��)�v�g3�/D��� �D�H5+�`��ۢ��OZ0��!_l�A�f����]7i%��e�{<q����*7�G���UW]%94��7��_�����/��u�"�D��BGG�e2�Bl>8�����N	�������8�4����*|�s����7TTT`l�O�⦴�7�xf46���Vl߳+���2���Vbszq��JG>�z���br�T�;r!�M�7�X��vBj��Z��tdJS0����b��jZ�х�B!�R`���z�~!?�����X� v�1Vas`Of5�c�D�s��1����u�a��p�i���@I��؈�7nD�`?>ڽ� kH���뽂�˗A�a^���O��y��g_l�6�R�墢�^o�g��a0h<�sZS�@@�W�{w���������Z,vE��R�����E^�	��)��JrcHra�
�%y��d�Sɣ\o�_�*�{�=�K�3g���͸��{���Jڋ�����|ݹ&�bm
��Mn]?��W���0F�Fq��	����?�2_)v�څ˼�!E��1���P?�ǚO���3��v�1���,��NM��4b2�(6_�#^���ε�Emm-H�"��P�B,���gv��y�Z��yq�F�v�k�z^�ae�E0M�*���'1��T�"WB!�B)$����]2��I���=G�X���2�J���X�.�!��o�=}F��!ċ�~����|���108�y���BG)f�,]�U��r�@?>ܹU:V)S�ٺ#�@��	�=��.]Z&WV>�o�fR�����M������jf�C���
������z����ۓU���=��'� &79i��&�Dǥ|��.�v׳h�"|�_��~�3����?���˖a�����������.�wYh�/�ҍ�y��m�%���k�E_��rF*6�Y-n����Çp��,)d����K�Q�O���q�rk��E��[����O�]���sy)��������[o�m�����Ė5�v�䔁�=�aKK���Q��!�B!����bv��Xq7w8c���gܮ
c������ ��`� 7��7�B
���{��sX�z�}�~\�Љcǎl��-��f��¢%Kp��6m���Rp�Q��i������eŽ]�|�'�C�,���0]?4Y;*�u��818-�� H~@�{�S2U���ɪ�"w1\�_$��;C7�&�c�)�zB)[�qbݲ[�pq����_�o�'��!�|�[�����9��`�����m׬�Ӛ�զ�^?0�.ȩ�/>��y���a�����ށ��tRP��J�>\��Z�;zXz*W��d�?�d��"r��#�ꯌ6��9�k���]m���H~#�^z�%Kb��K4e6/q���:�%�ԓ����h�*���LRi��E���aFz
�� �B!�7�xtQ=�GG�`��wFc�L�#c���?�oZ�O�q�L,^���mg�i��y���{11:�=�w3�L
�sڸq�ԧ=ul�B
��3-8�J�C/��SOa��ٞ2���z:vŔ��a�����ڡ���F5���8v���|��d{{ ͪ0��.�~�	_0&f�%	��4�*u�F�ae+Y�̈́�S�L�>]z�����	���?�^x�%�a�
�ӵݮ>�{��$`��}����̮K��a�|�{�MMM��� !^D���֭����y��؇#'�&�Y{��(�\�o�x��yā�#?�#�ā]{�����<���X�~��	�|po�'��H)� Q��o�>�-���a�RI��I��h���e�!�B!�����Fy�%�X�s;���G�~���������߽�PW_B
�ή.i����ͷ�
�M{�bdd���ո���ر}Z:۱��QR������} �Ϝ9s��/9ku�L>�^�1���C�	ݓ5�r�0&ne6곘.���a~A�{�ڹ�������ك����$�Bw��2tc�qdH�dU6���O�w��Ο?�ߴ�9�?��>>�3-�����vD�^wm���[�y���Mo�l�,�Rm���¾ҙ���'M�Խ�FEY9N�l�ɓ'A��5k�4AiyN�mAk�^�X��Xy���J-��{�)�}�ۂ�B�ZO�A[K+H�#�h�$�	�l�Ǯ{{bJ$��F�����0�1���$UM�\t�0IE!�B)l���4�ʫu�1�3�<������oS��x����(-���&�CCضg�T/��ƍ�,+G��f\�� !^d���Xy�U�Ǟ��z�K+� �P#p�ڲM�	��G��\[[oWD�]�v��G@U+L]?��M�1S,�1��}��{{Ee%>��1�o��@�~��[�J�)��~_�''��&��a�
�'A����K�4Y���TF:B!n����?��?�?؄EKc�k-���
%��R��v�kW�����Ѷ̶ɰBQ+�f�oZ��-�^<*^��S�-R�왳���##ؽk]H�!��֯��s18<�ǏH7)Q�>�bi�Ϸ{�g�<b��e�v%�N��m7�����^:0x��|�+X�p!�ە��H����FCjTI�vy���:1�LP"�������<*��v�B!�R�L�����)^?������Oc, �q�v��͟��2�^�c�n��Z�x	n�󓈜p�������|F�q�o����8�u�wn-
C$BM�wahp$�Y�v�4�"�|��煡'h�Ӛ��S�b����b)F��/D ��F�A�{��7´�0v�KW�ʉ��rP� B�ɧۡ�MV�א���BHV-��g>#%�:�������o|�hll�ϳ�ڮZT��6E�&������oI�j3V����Qj,�rO�4U���O݅����̩Ӓ�;� �M�P]�\�Vzr���f��k�Dd�'��Vb�;�d�oˇ�H1�Qa疏�kz���~멧�r�y!��dc{�c:S8Iܮ��R�ۓ�[�a�:���%Q�<E�k��p���vB!�BHq��Ӈ�+@c�,�;��1��h?{�����V��BG�S��ڤiZU���:4�O���V�ٝ�|bѢEX�j�aߑC4o#EG���p�����˪Q�����^���d�ڞT;Tc�9�����n��7G�A�
������*�9(�$��~�b�A�4�A�/6䠺c��t�tD�2�:�|KV9���M$����
$����c|���QVVf۵]��]�M��p쿤�6E�N�����ܛl@:y�X�vZ����ON����zά���#���� <���>��M��u��cz�t���a��#:Ǉ3�Xqm7� K"rf�C}[>�G
�=[w`xh$�� /����c��̼L>�{{��<!.h����)�d���B(�<Ġ)E���?LRB!�B��+�!L�/��.�˥������_2�jjj��i�i"�XÞ�E�_���G:����D!1q���*i����h�8�ͻ���b�Jw�<�>��O���ow�������{�D�PF�h��aXs/��j�����z�B�.�����?ͺa>B�{s�/�����`�5�����!��SJ'M���&:�������7�x�t����~��t�w�׿��x��O&/4-�Ά�n��4�u[hh("�)J5���.�V�m��-�+���%iz�p�M���;48$��@H6�E�֭���p��N�=cm�7����c�"�/�k�<bS�o���z)T�:��� ���k�Ib�̈́����:��x�ڹ]/I��*���!ɪ��rl:�$!�B!��8�W��{�<0�.�F���`h�+c������?����m��s�Ayy9)6�;;�I��7�p=�**q�B'���9�(q�x�f�̚3#�c8t�(�'�AH�2>6�[�J�'$�Zqݟ�v����2�A�0�+��>y4h�+�,d79譈�" �P�^�Oգ>�-]�V~�4i�x�Jvb�L>�r�A��EONViV�dU����J
 Ye�3�=�6mڄ��Q��g��&,Z���~{t�a�N�VbÆ�����Z�����.C��~�ɭ�/�&����NMM����uY��r�ףzZ5�FF��>��L7t��^��ƙ��%Q�����2kǻ�Xk"rz�{1X1]�!l?q�(�wx饗��M�M�{&����b����KR���A'��.'�􅘺\\}!�B!��������+c,@NI%jl�f��q�F�w�}4��#�Ò���{>%��	)F��ư�i�����7�r�UT���'��؝d��.]�s�χ��ͭ�q���;�Cwo�D��<�裒9����ro�ͱ���o�����C�(�iͰ4��u��p����|��gWG ��Sc�3 Rz���!C1р/�qc�%%��	+�EiE��e�7Y��g�E�c�=���� ��w��-�̙��+�'-�&�4g%������m�R��wuL�jr���N����T��܅�p*����PYV.9��kj���I�~^��j�_��RN�jF�Ʉ�׹�^�"�:����t�<����h�;�2C��سmgQ~w��O}
w�q�#I�|pYH�n9A��t��5I�ԉ�p�~U�k�UVU�g�~A�[!�B!���zMcISd>����
7�>�@����r�E;x�6n !�N�+�$�7g.��.�����y'���؝XF�/[����I�X�ζb��= �$8��	=�.�x���z<��3�y^�f=�@�cEEs�C͈ϲ)VP6�ү4�vy�ى�VL��'�C�P:�
i�$j�k���C����pc�I�>��/)Y�JX��(�udP�.�UNF�ɪ?��O�x�"H�#~�?����7�BccC|�%���tm7۬\�������ܺ�X�����
�m�A����Ϝ��WVV��O��Or2���!2��m�5kP[W�`�s�l�؛gW�n�rʵ=�eC�  ��IDATl"�hvV\�m��<��I�����9c疭�����<��+��M()�U"�M�v��
a��>2]�Jf0jPzm��ALU��w��uB!�B��=<<����$S,=c,�h��1���W�sh����vyޒ%K��O��?�!�7h>z\�s/]���(]�.J�@��o��NT�����?v\:��8.[���,FYE9ZεQ�N�mgZ�z��wx��g1o�<�_e۽]y�'n�d��%c�`B�nb��f�������3������C����>�H6�Tn�"wݡ#�/�$��am�V��*A]]^|�E|�{���9�?����k�c�tm׏�Q�F��3��)�76k{�Y�Zm��a�R��Ǎ����S�k��0k&���g$q�`� �;&Ő�@\#,\��W�@�*������V��m����\�Qlѻ�[�͇�H1"����;���x�'�|�V�ʻ�T&�ɖ{{b�:Yeֹ]5Ġ҅!�A1%����"��FB!�B�a81V9%�jc�tu�lc�j���C����\��ψ��=���������ދ��1Ca�E���/^�w~�S@(���}ӦM���(HqSSS������u�>�9׊-���b̕���Ň?�Ċ+��SOeT�K��u�Qc,����P[;L��:�X��1c,��Z����%�-@�
܋��ȕ`�z>BWΩ�L#t���nꄕ։AvqW���ɪ\~�G�������&o��ى_��Wx�+_V��s)X�"t�G�]�����iQ��uc͋E-�+K\��b8���A��	ާ���{�/�������L��ۋV�Z���֢��.r���.@{�<yL�wξ`��1�k��Xܛ�u�o���H�p��atu\ �s�Ε\����5�v(��:�v�ACq{.*�{䚤n�|�k���B!�R�l>�e�c�k�4�Jz-���o��oA��8>���<� **+A����i\�-���k�P�󣵵g#S1��q�[�h.^���
L�p�T3���3���a�G[9���>W*������;��.�굆X�{D�ڡa-Pa�7�
�`V�.^WT�c�y���
܋�-�{��k}��bP3̠R �n��$$Mʄ�ϧqbP$������gD���^�VBtA���� r���;��[�����m����ܦ(|W��&�oI��qk�@�4	J��X�b��n�����/_�bD�+WbF����bht��OCkg�&:���E���?�u�iIpo2�h[0�dl��G�����8q���I��ӧ;�(��N;�ɚ{�2)�K��6NVYua�'�8:X�0B!�B����mQ�n��c�4bw��'̱lc����5G��z��v��	�FGF$�����#���LNN�����kq�,�7��q*��11>��ǎa`���BA���\�e���O��`?�> ][B�#��w}�U��p�w���]�˧z��y	�XZ#,����X�L��)��Xf���~���H�C�{�02F�����@ii��`��L�������3�E�Ps`)��%IN�a�d�ӟ1Z~�u��/��/�_�
�;��CcC#�\{M�B��D���y���T¾��q{NE�ľ9�m�n�z^ @[������r���jl�č��sg���҂��)���q�L,_�\ri���111��p�+*f���)TTVi>�}���:��z}���Z�����C/و-D�z��i�.o�O|>���u7�ү'����{����A�.r�J���k����B!�B����YS�?��K��X�:���$��{���2�L>c�������̋{����8�w?���FB�#��:�IP[S���\��i�G�J�X��� �`ƌX�b���H紡��<s
m�1� �����	�w�Aow�w#U����5�\��ݪ+&���Xr��ԵC���|ߙ��M���c��p@��-�cK;���C������t��M9�pc�]܃A��#����� '�r���g�NV�Y�׾�5lٲ��� ��?�9���k�7^t��E�n���: l7h@6D��m���m
X�ؤ^7���b_��p�#!x畹����U�#G�_S��u�--�����K�`��E��������L�'X�=��Ll�]�5�F�k��u*�ccر�#���1�}�po��XIy!���v�$U($�0Ӻ0�I��f^���H( �B!���D�b��]�˰f��a)̱����V(�˥vqW�3"z�Hc�������_�"�����;�4�Bm}V^}!�14<��C��kkj�d�Rlhh�F�LM�|�9�;w��y���Ι3K�.EeU�8�a`x'[[1<2BHv8y��ZZA��3�<#�`�f���:�նd�X��XH�������+��~����aY�bwӽ�P�^Dt�Q5o>ƮtYrP\�����J=�bP9��t/��;�3�5k�{�9������4eee�6m�B�%��ɢ��,>���w�ug䦭Jg��{^�x	�� �F��H�~�/]���oɒx1��]]FEe%�	Xu�f�M���˗q��XŬ�5��vll�CCL�-�w-��ݗ��|�8�n��� �`��=�h>~2�J�D�'q\�~Z�8���A��zD�]�s������0��!��Abߋv��@����n19��n_�����1}�tL��������t3���v��.��1��T���+ǻ�d�F�.r�oE�n�M��K��S��>�om3�����,�@���Orw*-+��Nd�os���������GǤb�@|���?�-n�O�8)��������[�xN\cY���K�#�<�6�Ny[�VL0�ޮ~V	ۣ��p!��
���$UM�t���vB!�BQ��˟�1V�>-�1VT�l��́1�a{�c}��4�����CuM5�-\ B�}���p�d�V(t�.��w}Rʣ�ĥ��R-lpp�Y���1�|̚3%����.vb߱C��i!� j���s���W���<7D�N_��gǽ]Y7L)L�%ʦXAS�v���B;���i	�^��"cwO�Er��/'�R��eG��|����&��uqϕ�SɬG}���=
'���q�����+���9���.M{����Gy�Z`$������5W���wm7�֡�!�Z��T�i�]�N��c�����I+�9�6��
���V�]���4�DOw7��\��Z�V:���(��X�����]m�R�F�G"�_[�����1P?��lX���Zi��l ��K�q��qId..n ���&�����ݾ���*��+�G������}�s�Wr��Z��~����xי'��kkPSW����$��X�Yc����H��`�KǠz��T@����`����+�3}�F@�̊���M����F8�Ϟ?ב�&c��nth�sg�&��1k���>�{��Bߕ���/�;���DaA\c��8����ˆH�h&I�n�ׄ�2V������\�ɨPP9Ԡ~�*>_����` 13�X!�B!DI�H��K�Rc	w�ce�|�����/������4�8�-�wy%��v�m1i�s�p�� �PQY�6Vĵ�n���Y������S&9n}w��?�c����������TK�!��E�cU��,zr�ꄢ�%ȔN�b�h!�w˨e` r̷���m�ω�o&�/j�������_�W���n�ik�h�`�
C�Ҷ��Ν��߽y@4	3@7(��V<�������~w���3��[�}�%�n����[�Ш8Q�sω=7��z�B��]i���KU/L̯l��+g(n�
��AܺbF�.K���T�ܣb�`d�:2(;���KVes�����ꫯJ��'y�o����������+�����'��O@���N�f���"rk�o�?:<X�8+�L��+�{EE%*++��f�j^�S4��k�v���(�&3��+ȸMz����{yE�鄁�}�m��ݕ��'r�����G��6��:=rðj��(���W�Z����@�#�@� zzz�iddN!@e�_r�����pK��{����>�E���A��1�\���]����>k�D����uY;��ņ��w�l_�=:�a��5۷� ���K�.-�l�,e\t�v��dD��lr8��vA ��t�	�cI��>�w?:�;l���k,�z߭�y})�ͳg�v5�de�v>cڽ=6���$��*Ɂ!:iE��$��������vWL!�B!z����1V V7LU?�c	a{�����(F�{��wq��������<y*���+��/r��K)��-�N��>��&'DoKW������^�u�m�������{�H�Nolpe�Ű�+*���5�7{�T/��9v��%��E��!n_�t)�@�ubT��.SUU%�g͞���ӥ���y2�y�"�"�R_YU���d���f~B0�c��ݏK�p���qe�mE�ߊ�]���l��w�b���d�)�Z��k,�n�n}�[n���w����|5�J���ͱd���$Kq���$+j���1Ɗ�����`�>X�8X;�
�!G�����!���?���p�Q��r�HJ��r`�M7݄�~���oA���#G���������z�E���X'�Vb�������� *5n�Ia�c�{�";�s�վ�7u�Ŀ}���|�t�;�Pŉ���͑\�++*�s��	G��ztt��C����G� ��B�E�_r���	Q��|�+���ҿ�����$�q�t3��i6x�������]e�x7����oؤ��n���y�jl��z�N�8	�=6l؀/|��8+�[�[�:Ie��Ҿ�s`�wb��C��z�Ae�J*T�-A0L�vB!�B���@7/�����1V��$9���1�$nE33�ʤ�X5�z�W�)�l�,�##���|�{]sR̈z^��sҤdxh K�.�5�VH�A	)�	����w�=�������n!j�bD1�W���ɓ��7�O�c����Ckg��������f[�v���}�פ��e�ŝ��:���/IȮ���'O�eqa{L�n��5{�BL������{+/���"�dw �.�����dG�ȁ,:Y1iQG�����&�|YMV	��^�Un��|7q�۹s'._��->ڴӧ��M��lQ�h2�����+J�C�����[��Tp�Dl�ž�D��/�b��e�J)�5��
3������ʊJ���J�!�B�'}V��"���yrrb�X��A�?��>��3:6*=�,����P^8��ϕ��I���p]�c%�)v���X&M������@/�.v(D���a|b"i߄��kD���Έ������;�~��|<�3]�8��	�{������R��g3I���Ʉ��%����u�$����=��r���$F��t�I*B!�BIő�,	^�7�ҩJSd�/�c�����X�e�&�oN����!�7Z~�7JN����A�E_��ݱ��y!��0�j��@o_�2���^?���쪕(�N)�F�����X�(FF�1<4�9*�ΝB� ����	VuM�+�dX�_q�E�+D��}�҃��˸�y�4!$�׃��n�@_?��xꩧ�v�ڜ��-�n=0�g�?�V$�+m�Pg�gف]6Ē��)D��I1�`u�%<z	
܋�։�莊�S82h��"	��dU\�HV�fC)�2���7�l�s�̙x饗�_������_Gn&k��ڵ����I���R�l>֒`��\G���`s�Y���W9�g�:6Wb_��2g���H=*T�S�Z;�E��P�1S���`�[k��m�d����k�q�̮Լ��j�N
���H1#�\��n�����x��'�~�zǓT�*t�&���q�*[����uA3Ġ��_��K�w!�B!$�k��F�$cɓ�'��V����"�U=(�������،�v�؁�/�x����8R} �n����F��z��JS*D-D��b��Ƃ�3���e�ҹQ�ʅ)���d�%�#1���wq�'����K|UU��'&Y�xr*�y����Fϗ�u�q��(zGq��Kzo�w%��?��CW��x�b<��s�y�VC���V�ە�X!�)�~�Pֹ*G|���5���V�۽�E���)<��cÃI����{�{�Mwe��D�yA��Rw����7�)^7�͛7c��� ��?�9^��KX�d��ޒX7G�vg������x\+���%v�&"�����V�j���k��U������w�&X7[د9�ۋ�W�v[��l�uC��<R�g1L�f�x��z���U�vNp­��gI'a�����J��Jvo73̠<�`ii��� E�N!�B!$F�T=�Q��9V:S�`��/sw�c\�1Ɗ.J��9e���.�3f���/��������h>v�Ӫ�j�� �x�Oˮ�@���^�ԅ���B�8q�(Z�O�xq���o|uuu�����=.`���R�ci����J����X��@�ܣ��)��i�������i4�1p���INFn�v]�u�U@R�J�ٕx>��r��_�u�߿ccc �B�����_ŬY��L�Js)V6�S��6g=ָ�&��C��
X͋}aK�k�]�q��H�wq@�������e�x�V~W�`Wnk�7�k{rX~�G����	l۴�c� �C\����zWD����J$���̹��vaH��-���3�k\����@!�B!f�{Ac5`lx(!P�b)���^�1��ϸe����cӦMضm��8�t UUӰp�bB!�hi?ۆc�x�x w�}���Vn�e���bv�~/3�v�1��k��KY3���f����{
܋��<�d����+�U�F< �۳�������U������իW��_�2����{����G���x��WQ[[�i��͑�=lO�l_�k뀸=�"r���V�����>����M��h����T�:�ry���3��W�v��k;���?�ÃC ����ý�ޛ�$��I,{�ǧ�=�F��MN�IV��T:�Z��f�A���� �B!�b�󁙘���͚bY1�*)�E�U�Cc�_.��p��X��� �B��lہ��
̞;�B!2��.b��] �D�����+����!�S��S,e��h��t��F5De�P�ό� �۽	�E���*�5���]$O����:�g��R���v��L���~�����q��i���ׇ�|��x��PQQ����\ۓ�s)V6��-"7������������žV�e.ΚX8sa��X�������a��ߕ��6����V~�6����aa���k���#���Jw�7����kI�܈�3qoONRe$l��Q�$U
a�ֽ=���oX��n��B!�B��H.�Qc,�!V@�⮬�5�*)��W
�i�em�ʕ+���O�����A�����ܲ��̽��>�B!}����6�:�x��^z	�-r�F�d1�g�k�Ɏ����F~N�O�ޞ�n(���x���v�B�{��LVŇ����]ϑ�L�J�R%�����&��I����
N��h���Ւ#�[o�%�{�=:;.�g?�1�~���;#l��،u@��h��ľ��Y���m��0ڼ��l�V���	������^lA��[i�����ۍٷs:�;@��8����X�x1���J�<���0�k�U�Ĕ�}P��
��������~l�aF!�B!�lD}�+�)�9�d�{t~v��
]خ\�����1�ɓ'A����$�o��~�~TVU�B!����0�m�,]o�a�<��cyU#tG螬�1W+�^KN��XA���ں���L6���ޅw�JV�\܅�ƍ���=�^���&�R$�"�O��dUt�ۉ''�if�m�݆�~������MZϴ��?�',[���\۝���X-lߴ�7��{{�v��ۮ�F����&���kr�s"r'��v�wk��Q6��Vb�濫�!r�_�gl1rd��E��wY�v-���/�U*�I�D
�Iߍ��{�*e0Ġi�����fD!�B!���#�G���Ȑ�+��{�ߘ)V�+��9Z7L���XJ�,�C�	����䋉U&�4����*����9�>����>������B!�����}�c�c ޤ��o��&�������۔8m\�Y���a8�di�g�1V(�� ��
�I,Y5�#��.��d*Y�%����LV9��ufs�x-�U�w�Fww7�79y�8�&&q�'oW] �V�l>֎(�86�bes��D��������m��:m����(6����m�B��F�����Z��-�.,	��g��[���z!	N>��c'@��HN���ۨ����s:I�ny���$�R�0�JR�b�ȅA<����/�Z�	!�B!$S.c�ܗ�5�`�y���9Vd��+1�s�1��}�b~��4�~趉�NlS+��y���7��&��ضi�._B!�±}�bhpĻ<�����,�����ν=q��5���5ŊNA�Xto/\(p'�3Q��MV�M%�"��KViUJQ�V�+pqRˌ��9ud�d��ٳ��o���.�w�|�������?�c���X���D�v�f�i��L�+��ޮ�c�~W����uLD��_s��n�3�tm��`�����4�Ʊ��A�ͳ�>�����4I�F+�:�T�\�U&.V�TF.��K0�Mq;!�B!��a�cc,��{�f�_���{��`d�'��5C;�X����5�c��{����ě\��EYi��Z9^� �BH�#��?��W�@��ҥK��/���F�fQ��W�g�eT;jꅉ���a-��
܉D��*����bSP�̴�*�2Q�x��,�>�Kɪt��A�ne�C=��۷�����.���@MM-��.S�/:#`ͥX�^�~[-�+�����V�����LG~+�`�X������n��vm����$X7g�].?�b%��vs��m��=M �檫��W��U�$��I�l���[���J�����	�S	ܭ$��\��~|�B!�B!Y�+<��X��XA��(F{���BP��McA�WU椊�kƌ��7��w�yĻ���`���q�]wH�!�B
q���m�|Ļ�7��M��չ^t���&��R��bI�B�u0>�s|h���3"�
�x
�Ie����]�*7!|ɪHg�����i:��{�D�^�J���U���Ӊ#���t������Ž��	��� ����ǴiU���cr)^tB�k�]��{��&l6�}�ޜ
���/J5�]mÍb�z¬�݁�꜈܊�^g�#�{`WD�����4-�7�<]ۉ�K�]ػ}����;o��v�m���&��-7^g"A�c"A���R��HRI��{Ҁ�{�H7�7B!�B�;ڧLc��
c���Q����'p�d����K���{�̱���?�x����۱7�~K�\!�B����۳m.^��6�>�(�㎼��Z螸oӘc)�!��hv�g��=�R
��5�3��y��
�Im�J���6Q%'��	�H����d����OV%92@-p����J2���ϟ�W_}����@�Ϳ��_QVV��6nHZ朰9sq�mn�v�[�q��[��Tp�Dl.žf�d�N��ڦ8��wuFDn�����|Ws�����r�8ЏP�m��]�c���u.�6O?�4n��Fx)	��$�n�*�dօANRE]�e���I��PZ�Öv��!�B!�;t�g�.�1��n�o�ҭz��n�1�ۗ����ۇ�/�x�s�gQQY��7n!�B
������<��Y�p!^z�%ռ��«�_�O�ꆖj�s���=1i�i��ۂ��{{a@�;Q������:�{�2Y�OVE�4��Һ1@�Z�O�OV�M,�˂��Gy[�nŖ-[@�Ϳ��/Q�+���I�s)lvB�k�]Fq�Xu��ir_Ym���vY��|�iC�����pm�ݼM���X��p��|�� �"r�ǻ�8� G�Wa��}���:��;��=ر�c�:�x�U�V�^P�s:�dkv�sI��bBJ9A�LV��T3��UtJ���qo��%�B!��Mv�O�E��a��{�W3�����;i��+�l�o���x�����~�9<�s��I�����ցB!���}�z�������ַ��А�5�t˳UCL���̛b����X�b��a����D��� ����Ã�d�*Qe 4�&�CJ����U�ӑ�L��� �K$'�F�*%�$\7��L����W�C���������%%��\���gl����R�l/V�����\>�`�fŵ]3ۑ�J4X�Uf��ι�g.87�Wf�oi[0 ��y'\ۭ�Zܛ�3ږ�8������I���1jڏ�o���x�W\o����4I�+g{I��ܓE�	�3�*���b*+�cS;!�B!�8���#��qwq_��c�
����h�Pi�U��7�
��c�Q��*� \�E}�h��>(c��O�6����k�_B!�x����Ա �G���y�y[#�E�j�PO�.&=S��#{�����t�b:;E��B�w�ĩ��\��ڵBw=�A���/����dUII����ua���P	ܕI��]۩�p=��F��-�׿�u�����@������?Ǔ�|�פ����t��D���;�M�5�"rb_�X��]q=���?�"�,�9���J��n�9q���ݠ�s�A��{�M9"Bw*� �W��~�SSS �����-����$��$���'N*�ۍ�T"9��T	*Iܮ^0_@�aF��N!�B!��4�R9�+G�N���A?|¡=�F~����X%P>�4�����(���Wu1a{���HUK|��7%c�K�.�x�cK�?_}�ZB!Ļt_��s�gA�ς��+��լ��ܮګ!����(5���Za{jS,1�s(a�%Mi�Iu� �f������$up�����R%�dwI�KT��jGw���&��bw��aMG*w��y�L,��f��_���Ȱm�6o#��_���x�٧q�իuc�
s&��Ю�X�f��ka_e��ᤰ\�R�׬���j��:m��m
֭��M���C#������k{�D���\�S�n���~|��QV�۫B`ٲex饗T�
=I��<!\�bJ/nO���VJ9I%����k�������gB!�B��D��zMc�uÄ9��K9�s�K[/�k��$���6ƚ7o�d�����f~� n���Zk~�gB!����N���e�#��_�u̚5��̰�����L�Rdc��4#>��
c�c#3"��!]!A���`�/G��D�2Y%��+�Vqa{ܑAt8%�$UB�LV�"�'�d�{�d�]a����pQ��\�Z�-�y��8q��� �F��ӟ�+�=��+V����;&`�)��6�u������V��K��������oC��9�v�+p"���*�ǻ����o���$C����������� ������QWWWTI*�r�	*��[rp���bw�[{��������1YN!�B!�9�1֪es06xEe���i��^����!���	��XJS,�1��^�c�|�+���L�6m��}�; _��Zy�U �B�w8}�$�D����� �������_�fX֖�SlN�{:S�ĨωZa(6iGz6����6���V��*0�.�zX�b.F��S:2(��j7B�`<i%:�D�x-��:2��hE1R���9%����ƺ�b.\��^{����(J+ ĉ�g?�q\�n[D�+��v9&`5�}K^'�������)��+�ς�ּX�¶��n@��k8���`�ǻ�:���-���m����h�ُ�5Df����� ��3�<�[n��I*��4WG�n�y!�����`�A�}մj|p��vB!�B����,p9�K3��n菊��џ�I%nO�9I�Y�V�n��i�,�j������-;v/^�>�4I�,[��B�Μhơ�� �����曖�J���Ś]nv��{0�Y��!idg���Jc,i��K%rW�cB���5��@

܉!�z����r�SP:2�ĕ,f�
��Mv0�uc�%%���:�*ّA+p�]4�*iN�U��`%q��#����	��A��,r�`�U�����-�mp-ę+��t�Y�w�x�岀�8.�b_+�2km_; ���k��v9�]ͭ���n�̩k��88�������ׇ�� ���5k�}M5/���F��Zn���6Ġ�켠�'�0��I�v����{������@!�B!�@�K;��v�g�1���}��?� ˧�WL���W/E&�|��!
���Fbw�c�
����*�r�عs�⭷�¿�w��0طs�t\�XM'wB!$�ii>��{���G<<:s�̼���V���Q�c���P
���c��1�^�P;�s�h9Cq{!B�;1��?��W��ؕ.]G�N$���qd��yr�*1�`A+t7���Q�N5_���l���7��<x��� �G�|����K_yk��F7�PD�+�ѧD����E���C�{���W�u��p�v��3�[�+V6�x.E��(�7g�K�s�u���n��X'z1ؼ�u5}�W���͘���`����_��_cڴi�'����̓X�$�4�t�Jx�T.�@za�2IUS[���'at?H!�B!$�$cE�ϔ�C��=n��u����c��d�1��պ��>�ܹ���oA
����cb՚�A!������q��px�'p�]w���Jl��'��4�X�eP����c�ҍ��c�%�p8���@��w��m+pCyX��
7m'"'���x�*�Ŝ�J�z�DבA%r�Z�''��dU>&���,X��={6���oKO���G���;��g���O>���U-���R�k!Ζ��b�Y�w�x�eUpos��ͥ��l�>n{_g_�O�v��լ�����>�um��_e�d,Q��݃m�6cj��х��/��k���I*�$���~�Am�*�HN�sa�'��΅fE��c�B!�Br��+3Ē'�{:�n(��*S,�B�����tE�P������r~!���Ki�u��9�������I��ukA!�������c���R�PI.�~n���k녲9��ڡ�^�1�
&j�1c��|�)&z�&y~��E�<Mq{�B�;Iɥ� *V-�xO{\Ԯus׊ەw��Ȑpc�&��Wrr*���:����qd��i�l:6�����;��c�ᗿ�%Ha ���L}�Ql�x�����be�dEDn���^�������|��}mM�6g�ޜ>4����޶ۇе�|�ۂu
���s�2�o�SS�7�t�|�ɬ$����R#'����ҭ]��JNV�D�DSHG؞�ĠMRń�u�x�,�AB!�Bq�1V��K�n��
��_g�gq��5�J�F�!�S}��^W]C�Wa���Ϙ1���|�M��A
�c!9��n!��>��&R8���I����Ei��~��f�6�
��^����>�cik�w��β��� �	�$-�;JqG�/1�b�Ay�A����/��Tn�!�*��]ב�DUX���I��7�M��qdx�Wp���>}�p��_���w"w%9�Z�sB�nMDn �5)nwFp���v�ľf�d�q�b�����n����k>`�_0����k;1I�������X,$�O���|�;(//�]^Lnj�:Ae͉!�vl�b0*r���%��)�o���wB!�Bq#c,��]�n�0�
J#?�����F�P��k��O˳{뭷⩧��O~���A���q�n�B!�=ăg'�),��ylܸ�hͰ�u�dQ{�z�~�P�gu��ص]�*k���a e���}���B�w���� J,B���:I��jWԍAv0(�3�UQg����]�l��G֯MT�'�	�BsY�[__�o}�[x�7�.Z`��������ƛo��;#`ͥX�\�Q�Y���j=/`5�]��S$���Zi�~��6~���bs�Ј�{{�tm7�`��v�tu\����I׺���u/[�,��'+�NmK;�t�
�e��^�*�����$�ERJ���k�K�vB!�Bq�$c,�)�_�K��Q�ea���]k�%���
c,m�P�0(c�+��n��Ċ�/���d�u��Q�¡��q��s���@!���spOΜ<RXlذ�>�����/��-+��"we�PY/L�9$��
��k���:bd~ii)6��"�
�.�S|p��5T�9�+n�:2$����z��%�����h+w����\����zo��&��_�%�������o�ѱ1|�t�: ��爀�R,xs&�7�|���Ή}Ͷ������y��.m͆�=��u��+�����ݬ����Vb��o�>�϶�i�.隔��?>�����a!�I�t�R��k�JP�qbH��S1��ƠLRE&��4PiGQ �B!�7Ic�%��1�{@��T7�w�)�v�gu�Pk����'r`�#@;e���u9e�%�����o�����)N=���Il��ƴ�"B!�dq��o���i),jkk�Q����t�Z�0�1�y��u�䑟�\�U��ͱ�
a�4?0�����f�С���bl*��i�Q��j8�V�.�W��ew�h�Jv0��'%��ve�
��]�ɪ\
���v2�������СCػw/Ha��O`|l�>p�o-�D�+�ͥXY'>+"r��\��Nۣ�z�vžV�e>�����~�Nã��'���9�v�v�}��v��S�n�ph�>��dѢEҨG�>E�n�\�q�Jߵ=�HR�9190(RF�ve�JρA̯��g�P�N!�B!�����x�1a��4Ŋ����XZS,�޸n�4�sd����+��v������/����RX�4����>q�-�<!�B���.ݳu:Ν)<^�u�^�:oͰ��fo[	х�V����k��uG}����+놱��beU~�RP�NL�Q[��c�#�"w�$����/;�xMR9h(r��EJ^A+�R�28�Ȑ/ɨtɳ��r������y����;�n���y��O���-��gE�j�bs�4l�M��6��V�����8�؜>aAp����ᰅ��S���u��������o��\�aA\O�������.a֬Y'��rc�e��ȁ�8A��� '�B�2��/�HT���-��!	!�B!$? CUQ��b�+�+����퉺a��ݠf�CΡ�1��"y�mx��gq��alݺ��h?ۆ��n����#�BH�ײ;�lť�.��C���裏:V4�L���rum��K�~�5��3ƒ��Q��ͱ�������%�
������&�Z�0+0 i�4Ԡ$lW$��L�����rP��Ҿ�R1���{ul�����B��n��Δ����WU�������S�o���\پ�nuuuV�u�L~���5׮M�ʐ��t^�DӮݖ4�ר]`��+���뽒r�[��Z�|t��ȍƁ�}iV`e�fE�����FG1<4�.f�"l�t�PX����a�m����i�im���4:2*��=�=o����	���<r��:��M4�Jd��GO�ޘ����H��^�S�2+}~�n�/E�r�Tl��N�Z��u���`�+�b����z��0>:�����vڝa��M���D������]����9��k�l^gX��k,+�^to�����э�n�J߭�ع]��ҋܵ����%�롸�B!�B������z�������Jc��џCIuô�Xr]L!vO��X�XW����"g����hmmEW�Z�%�=�@n�[ۗn��gc�Bl��͸���#ksy��t��S汝��m��}ї��}�������&���}����u���nQ��;����oK���?55��[������y��k,e���k,+�~�x���9k�z����5C$��qm7�9�9V0f���W�����Sp�Br���������MRi�Ը2�_!|(jP)r7rP�����EC4f�+C��*+�n�,XIb=��طo��_�E����/���}Y�499�����>��]�����?��+*5K�_B�~��7�^�i'n�߲r�'�`�B]�ё����x��v���7���k��� z{z�l���Z`��TN�G������P��l���S�V��}���`�X�OXqm�zq��3on��n�l�Ѿ:q�(��vmR��m�h[��B�~��5�Ӟ��ŎNT�֠���DK��6���i��/�z����+þajr
]X�|���M[��]��9g������/]�m���J̞?� ��};v�|۹����5V��3� ���<��5���w���%���S��1�KR�3�q_HNVA����MV�0TTV��y(�B!�BH��%8=5������]���9��9�P��n(f)k~��X���&��9���K���s�J��~��q�����UUUp�Wrk�⻋I�?r��l}����ܼ˯Ziz
�{�q뻋<nW���P��k��藄I����]��pd��cc��OF�\��B�.�P�P���y���Hn��&&091��b>���vdx�"FI9{����-��ݾ�rs�b����)�73�7���=˿���3g�̉x=_j�Fˣ�Sl�A�P[7T��
�{0.n���H�4�slY����v��^,P�N,��W����h�#r�&��	�`l����];�`ԕAߍA�����G;^�s��s�@�溲!���|�M477��ѣ ��pr��?� O=�4jjd!�� �쵣ia{4�\���2k��7)̵)`�&��<.ulvž��F��]������n,�"�p�^���� ��+�;�Ě�m�A���m�9�sK�7Ļ?ކ��N�¤����***t��C���Z�`$hW��]�b�����T���0IE!�B!�ȡ�SX�|Ƅ1���]�k���~1O������亡Rخ�
i�Os/%yh#c,%�P��.�m�뮻��#��?���3n�&���_YY���)���NcMNM��ލiiFz���h�.\ 7���K�-��~�i���]�~1��˝QSW�i5��w�L�/a�Ⅾl_ț�.��;257���Z<P4k�W�`�q;<4���lK _��X�K�󸅙���+�ছn�k�s5B��DM��+]�PL����>k����55CQG�m���-��˜���U1�ۙHRiD�r�J��roW���C&;2$�1�ܣ�&�2h�UN%��-�E���jjj��|/��2FG�y�8���.|���{<��3�5{V�r�BIkbes��D�������Vž%ڇt���V���m2��"xgD��*��kǵ�(�����dlV���~�@a�;ǖ�~���+ ���&��e˖e%�TxI*��	q{����=�Z��J����B!��Q�^��5%=�{=IخqqOvr�Gk�:"�Ľ��nhd�%>�}X[�g�%)o�sQ�溲e�%�<'O�DSSH�!�r?��p�=wazC!�b�+=�R�pb|�0���[�r�g+��Z�\/���OV��ʚ���];�sP��rr�N��zv�L��͝�S�;P�N2bsG��E�Qr�J�ZύA9�V�.'���jG=7��]�.|Њ�ԮF�^wY����k���^�����0������ɧ���K�H�r+V�k�V�bߜ
�3�K��7�6.u���������pm7/X7�!��|g�0�������i������N2B�/l�`��/)\�x�	�{�YO6���l���H��3IR�LP����TCtU�` '�9� !�B!��;����a��˧c��4��5Ŋ������Fu�0QKT����ʆY����+z�\��X���*|��ߖ�����A
a���p˝w`�� �B�y�:.`���%CR��Q��~���9�fX�c��v(���^�P�KYC��S�c鹷����q���b�w�}c�Nh�B���K$��!	+��]��Ҋܕ�Ɏ�"w��+������1q����&����СCؾ};Ha21>�������_�UW�6�9���,��͋E-�}=/`5/Vv��<�Bd��F�Έȭ	�Э�߆�ݡ�Ftc-	��f�os�o���=z�{�c�G���.�AO�LfՁ�knV�T�T"A�.I�/xOva���Ӹ.���uU���p�CB!�B�'�X�����u:"wm�P�'L�*��N�rmP9����]4FQ7L�?�Xn	۵�W�Z�7�x����@
��T ;6��o���ZB!����L+���#]k��D�S��=���Vb�yz�v�	�z���=Q3L����Z0�Ҋ���~ljRg���$c�|.��ά�7�qq�KX%�%��q��,nOvd�{-�,����NTIsJ�;2�C���甯���s����R����?�'����q����/V�k��6)��"�Չ7ܺbSU����}�����.&�Ypm7�k"�|�� ��+�����Z����ݢ������B�SWW�����AmmmVSVב�X+m��3����+�Uz��PH� O!}Q{�vщnﮎ���B!�B��d��`½g�5Ø)����]��=^/L���X%I�v�~5��a>ce;�����/H�X�6m)L��o�n�����ցB!�?tD�Ha#�a�ﾜ��|.����Ê)6GY+Lc���#&�#?�������u�)�f,��e�ۋ
�I�L����?�HRe��.%���VF"w�9�SB�r��$�WFu�%���Ƞ]�f�w��믿���1��������Q�uϧ�cS�}���Xk"rb�|�ڊ͡��t���Z��I�$V6k,�\pn��r&��k�w��������e�:�7P��.gN6����ܷ���׽�W��zb*�r��JvbP:�+]B��v#���{{E�"t����B!�B�ğφ�9�059���c)E����h�P�9�1�@�.������9�����&���p��a��E��FGF��OH�!�B�k���p�������ǫ��j��M-�Ͱ���A�9V���ܕ5�T��t�XA��]���V�k���X����b˹ ����Ã��+V%�����=��23�`8��F_G;�h�N^e#�n���(3�'l1����������6t_����(*�˥yFb>G��a��w3�̱��^���J�v��	��	�ai[�b-}W�������[�׹��3��G��C{����S �ϓO>��~��y��2�l�!�I*�����Cl*++æv?8� !�B!�x��`���P5r���ݴ1VL�.�eq�c�D�Mm����Lb�~�h{b���|�;x�W088R���i���(n��(+/!�B"װSS���v\��	R�̜9S����:�uA��p+V;O]3��6�֥]׹=ͨ�qQ�A�P�=K��X��������^�t*�����\��{ّ!��J$�tE�vHI*��=�z�A�d��$�2��x-�\9}�4~�߀6�O6�'��<���t�[+���&"� ������w�/�5�&�u���Ní������[����r�x���,<a�m����{����w���� R�lܸ���ZV���в�^��&���ۃ
q�����
�������1t9B!�B!����|i�L�����6���}�Q��N�F"�T�X��f9�m�+۱�4�J��5k���������2/Y�\�Ѕ-����.�}~B!����0v|��|ȯ��b��e˖e���K3,+����R-��#��L�5ĠB�n\?L��{]�8�R�^�P�Nls�7��V.�ؕ.��=#w)a��ۃ
'�dq�*a%�MZ�eRՉ�آ8��`�Y��累�z�-���p��"�bg��������U��X-��M��mǰ]y+`5�]�tmOw��5�Z�}mW�l.�9y>
�a���U��w�߅��p�\ۣ��
�YD�>#�����G� )|�����i�\ML�C�l%��\���r�jjJ5��n:�?'�T�Y!�B!����f`U�7zߧuq5B!x7��^�pq��C��aJ�;27��D�^�X=��?�_�� ��@_?6��'�x�- �B���������s�<����h�{���Ųe�5n��n'��۱c�]����q'�7{��&q��-�Mb'��E��"�V�3��f4]���$H |A���_?��_�8$p�������E[k+H���_�:.��Ҵ��n�ͱɞ������fuC�`,���v�>��m���u�4�g34�Wx�X�/͕�U�Rܵ���Ƞ�T�X��Q��-��`p�V8�PY��;c��Rm�o߾X�r��v����w��Ԅ훷b��Q�>sf‴��m�}�2�[��X��,>V6ҩ�W~LV_B����#s�C���+2�po�`�}��������{ة9��^쌥���@����U6 �=V�Z�4���	SV�K���"���=E�����,�=�\;��t��B!�Bz.�;0w���W�}ƚa��^h������#���ڡi0�keU�ĤC���lƺ��;QQQ�6��nZ�[��;�0m�t�3�BH6q��!l\�!:C�&��w�y�ַ��[���`�a����OP���bi���������G��8PFs{�C�;q�ږN������D�J#H%�&�q��,�A��h�*%�A|�
�{�w8!�!6���Q2��7}�t�X��>�(�uY��{y���ŗ_��˗şH��ܢ6��{9�M������u�Z���������mwbnw�p�}ú;�y�������/,�Mv�Fs�&t����8�M��|�������&.���#Luw=�"U���^2�R�TS{<�!Uz{�wc���!c����vB!�B��~$�S��Tc{P��97e���f��S����y�u%��4����R��ѓj����x衇p뭷����w#L}��+wx�5o!��l`���ʃd�F�>���BW����o��V��J�JR7�q���Nmb{����F�{A���k�s���B�܉k�q�7�돖3g�b��ԟ������}�V����U�
�J��"�����.#�����g�g�������Z�:N?����


���Dn� �7}�t�}���6����]1�K�:1��l6�x_0����1��ذ�����o�I�X۽A�^wlފ�;v�d˗/WZ:����nû��P����<���Š��=77o+�:NތB!�B!��ƶN4�����xr���.��Zab�0�3���@ch3�{��`,�8k�XZ��	vw=��9a�<���(�TӬ@���46b��s��SB!�7�b���ء# �A~~>V�^��cǦ% ��6����x]PolO�e�On������n�ţ�t<�ڙ�Nhp'.�� ��:�C��D����hnO�ȠMqק1$3�KD��ஊVF�JY�"��e��]c�v��;�@YY6n���ޱ�+�p�>��*˜���ߣ6̾v����nS����gSj{d�3c�7&�L4���&r�72Xg�8�R��p��:�����B剓 ��ȑ#�r�J%�A�Fw'��c�w"����Bz{G���`B'����vB!�B�M�q�7��֦F]�P<�њa���њa(��J���܍uC�`,q���3��Z��'B~��_�d�fC]=λ����B!�7!n�����P_[�=�~��X�ti���UO�_&���2b��j����ϝ��B;�v�(�? ?$�>'�!���U������#�\{���nLb��U�D��`��McP�`%�	k�*�e63m�Ay"C&�QN��2����~����ѣGA����J<��_��[nI�86��0�z`����n>6�f_��d�M�fa������Æq�o.�lX�3��k55�{pӈt�N��n��K�/���g�$�hll��-�PWG�*�())Q������0ee=#����w�z��L�
�E�N�@��Tک�QR�9 �(RB!=����Ĥ��<�~Mc3�����e!��<�� ����Pm�����Is7�ۭ���]��)�f&�ȱ$�Rki�e~�e�QK��o��ػw/�{�=�젮�o��*ιp9��B!�7P_[���>A[kH�p��_���Z��uA���f�6�*�e��l%K��cu&7�'3�wv�����1��D�����;'���(�w1�Z��)w��n�b����Λ%2�1���99�Q�Fa͚5��������4�����w��EX~��'���XG�v��v_�|�S����6���ڃ����v;c�,�_��~�aYr���s\q;�q��&t��{=x�?ژR4 ���}�=�`��i�������*.T�E�pT��=$-�*�Z�23��$���0�� �BH�c՗.�]7/�|?�'���_�B�;!��@v�`�)��RsR�wY���n���)����F(3����w�6�ҭ�QMЭP+7B������#�(ɗ�4���ڰ���0k�\L�}!���̉��Q�g���F���3g��{�E^���������_���z!j�F��ՎϑyC0���Vh���â�c����v�w�:UM!�G�C���������X7����V�J0���ј���^�R���Cvƺ����c�/V��x�	���7�F]m-���ӊpiĺQԹ)U���{/��1�¡���1�lӱYءa=#L�����3�1��X�n�ph���װNc�w�����۰g�N�|S�Fz/_�җp�7����%�)N�����T:3�{"����G��r��	!���H���o\u�r���/��N!=�7�by�x����n��9�f��uj���,��=!K\�F�A��}�Xɶ7d�<��c����ǎ�Y������4��c��%��+!�ғ��:���Í8~�(Hv1x�`<��8p���@7�v���}�5���p,�P,m0V(V?L�eZ7��H0�����c]G!*4�OX{�׎*E[KK��`�`pO��I�*c���@%��2t-�Q?��I>�����2]�rc��믿^i;��?�$�ؾy+N?�>w����g�a��!�ސ�.=V�0�ߵ3ú�q^��~_a��6���������a����F��{��=1�3�=3��{_��"�����q�m��fn�4a��zFTS{�'$�T&�,���He�����ݿ(RB!=��?a���*_��b�����yI�y	!���Z;=�>�7�Gk��g��Ě���,�][3��@��H�0��n��il�n�k3�ټH�|���z��X]�d�*�Lc#ν�|��B�	4�i�o����Z�d"�}ժU�:uj�jz^m�ͱ��`�?#�2�	�?˂�B��ϝ���p�Q?4u�Lo'zhp'����cx���C(� Ms��U�D�@@op��4���(X���+�����l���]w݅cǎa��� �E�J<��_��ǔi��w�d��4�:4�:4����q���N��f���Dnq�w���o�ll:Sϥ۴�[g�/�����mX���[j�k��;�)B�>&L���+W����u�(S�����#R��ۥ"U�4��؞�ܮ�0x"��in'�Bz��~��/�e�_�|!�]�&�+��	!���ZE׍ꋶ�f��ݐ䮭ƌ��Rj��`(ftWk���������;@�c����ow=/��b��+�@YY�}�Y�좺�4^�e�s�29�BH&s��1l\����A�q�*B�.��b��~l�;ce����aX�B����`�`��,�=e��~����Dhp'���D7M����q��!�A+V��Uc{ "TE�E�$m�{��nfrW�*%�A+Z)�*eI��D��y!@Y5ډ����x��q����� �E[k����������/�T�{X5|���z������qfc��ߵ������{a��s\޼V���x���3�xKž2lٰ��QYJII	y��92m�t��)��H��,}!��S�J�0Oo�U��E*C���~���
!R%��B!$�)꫾t����+#/�I������1c��Xfwy�� rB9�za V3��U�j0VHW'hk����X�]��ڟ��X���wp��!���� م����[�9w��H�qB!�F���޶Cy����\~�����Z�ϫ ,��pg���]b�2��)�j=��eLm��
M����a(�Ζ�]׍Lo'���N<卣�8�_^L�2�2�&24���P��Z�*��b��`k9���4.^��Ȑ�t��lo���X�f��4515���G8q�8����������J�6lX�([���jl����t�n~\��)B}�`k�dr\��n�ܞ^ý�qfc{\j��qf��	Ǧ���8
'�!R�?��n:z�0Hv"�'z�!,X��w1�+q�;�ӟj�E*�$Y�Q�2m-hG��=/D�!�!��Ƨϙ�}�*d"�=�ƃ��x�E!=���A̘2-5'�>�5DmV��.�՚a@�HLqצ��b������h�{�D���X�XK������h2ǏǮ]�@���صu��U���KQPP B!$7bmX�>N?��̝;W9O��Km��DӻW��k��p,+u�x��������X�Q<tv�gݐȡ��xJ]k'�F�EA]������VB�2U9�e�XZC bp�ъU�R�J&X�ZF�*dP"COHg�7o��^<��� ����G��/��u7߈q�G��0�z`�M��5�f_��d����:�8�d����&����{;��a>m��fc���Ә���F�t�%�i�o�＇��z��E�/\}�����NaJ?��7�T	���ʘ�.�%�H���`�͠V��Η��e�!�����1C��)N�*kϠ����>EJ���M��ꕋ�)M�ҳX{� �W��]�U�{b�{��ܣY���|(v�,ȂX?������ ���[���ӠA����"���$�8q�^���8���<t!�?9]Y��Y�֖��d�СJ������Rt�.hwɞ��!�j6��k����ΤuC+�X����	3;�94��y�`�L��z]��\���\�J4�kS܍b��`�&2h[&&2º�{J���H6�u��ȑ#x��h��R�����������/����V/��}�=��jݬ�ɩ��֎�dޤ��7b�D���o����W&���_��ƍ�2��mX�w���8��nT�I�r����[oU�T�0��-tuwV�K��� TI�)Yz��0�D�Z{8�!���C�����Ϣ�8uJ�_����?!w���|�R|��L�&wqJ���O�;!���:�P4E��	]��5D}�{0�f���F�?�dŮ����o"W	(�1f��=���t{3f�P2W�ZE�.Kiij�;��^��ӧ�B�};wc���9�N
�f�L�<��Z�W����/~��<���&wY�P̧LoOQ7�.��b�Gu��q!,��^hp'iaC�@��Ztt}@i�۵FwU��&3��4����V�2&1Ėu���I���ԽD���2�2����w�m����/��H���{�D���p���g^<41��-�S�&M���}��i�������홅�7��D���{'۴�z��n:֖���X�oz�3֫�b�����O>ڀ#�d7���H`���8�M�N��۵g[��s��`\����IA��v���"!����ɭW+	�xm�~W�����2Mfr���$w��	!����� n�4��5�:��nh4��ꆁP�~��#m�0bt7��wH�z�{dU{�XZzc-��K/�ѣG�_�$;W�?ڈ�'��slkv�BHwikkæ�*]EHvs�]waٲe[t�.hoښ`<+fj��eu�����v�h��n��>��W�Y7$ɡ����C�A̛2Շ$i�C�hpWD*!V)�Z�J��`4��S�-U�
G?�ӑ�`w=?��V���Ã>�S�NaӦM �ˑC�������3�2}��I��^�#ce#�}-���k5ݗ�C-�����5��ȭ�����o}loHm�o�}s~zozq�M�=jNWc�{�q��Hv3z�h��?��|�2C�21�kE*�8��Vf-�Ȕ*�!�
V�����!��^�.���/��r����q�Ϟw�ܮ"L��<��뗚�&w1��y�&wB�!|P�s��E�����=Z�D��ω)����ƚ��XWR7�c4�{���6�3�կ~'O���������#����9矇!Æ�B�ʓ��������݈s��}�s�������6d�ˌ�aX&uCuj��?'��Z2s{��]�%y]e�����d��N��+�kF����-1�A�v01�!bj���S�U�p�ܵ-�P�2E��z?���J{�;���^Z[Z���	�/�%�]���|O��5����k��LVwlvnX�4f�C��pg�|�u��5la���s;�צ�-���arw��c���w�:���S�g/�m�̶�%%%x��G1a������D*c{A���(X�ZS�۵"�jt���!���ŤQ��䷮L9���_�8���ٱ<��k�V{�u�&�/_�P���N!=���!̟2A5KS7��Le&w��5���H0���Y��vHk���ab0V ��"�r�&�F�/fv�*�����Ǐcݺu �KKS3�]�&f̙��sg���!����=�wb����\|�Ÿ��L�9�0����2�^A�SQñ��C����˳4+h^743�ñ&�D9�$54����
�@�H��Z�Rڵ��JIm�ܓ�UZ�J[�5���T��Ƞ[;�(7��8?f�<�����;�����l��	�9�kn���=�.����X�H�f_���V�k�fe�c�3�g����؞��ng�s������;��=���l\����@�8�衇�hѢ�	PZ�����خ~j&3���0��
f	F�J�fP*Ti��(RB!=����ˊѧ� �����%%��k��k"��^w����	!�g�jE׍.U8���ܤ�X��a �Zu��U�;�u�x�0~���nOW�΍mtw?��Y\\�tݻ�s�N��E�}�ںU�*�d�y(.)!���MM���Q]YB�̙��~��kZ2����mĉ��5�N��C�����3VC4{XMn���S��uC�IRC�;I+�Ot�)��RsR���L[�)Q�{ fpW��D�J+X�S�]"CT����	&w��Tx!n���s��G��ի�/��T���s��k��EX|�����wFSk�v�f�LNmO=z�ޘ�3�p�d�f�k�72�`����Fg�o6֋��3�c����7(�~���~;���j����2���==Zc{�ܞ*}A+X�j�Amk�Dc�Q��ۃ�!���g/���SG����o���lG���o�*��^���~��?��w@!$�	v{ۇaL�AC��\������E��0��H����ƚ���VX��9Z7�c=+k�^�E���'�?�:�Њl���)�����xٹ9f4!�'=xX�v�{�5��F���{��^��`��񚠾fh��n���vh��nflW�C� v�C(L�!��$�y���(\���L��	V�x���&�!�X%H�Ȁ�K�D�G�S�exe`�2饗��ѣ��/~B���ۯ����e����A����O�0�ה�.���X��պ��� d�2�D�ý��N_�ߩ�ˡ9ߖ�^:�:��CG{����@����_��~��ʹ��_F�t���T�Jan�	Vj�A}�A}kA5�=e���k��H��u(B� !��sҿO�1"�}կ^A�Y��4��}Ҩ� ��3�q*��SFG��D��^����jpW놱���y�g�����b�BE��1������<K��D�ꊓ'OV��x�477�d7mmmX��;?y",9y���B�k��HII	֬Y�	&��������Y���u�XH^C4��uB㼾n�t6�
�������C�a�~�ۉux5A�NmK'ꇍGq}��Š*T��d&�@�����rbI�r�J+R�%2h���8Kd�� 姙�l��_�2�;���<����Y|��q��Y�1�X���{Cj���+����p������ՙaݹ	^��f7=��nnp�p/��g�홅h'�q�8�x��,[���{�r]�=��nu2c���l�����a�մ�&0����S{L�����D��!㱻��vB!�����w�y-m����}��;y$!��|�8V���Eꁚ��1�]\�����X7T��dݟ��B�k*OrWǨZ�{�XN�ᗙ�l����Ê+��SOQW%
�����J,^�C�!�b��Q/\�z5�>�l�k~^���-��BM1Z������e���a0�v(��l�vD���x퐰+w����N|�CA�2y8��N�����hnOl;Mtb�X%0�ݵ��
VP��Q�y"��Ft���"N"��>466��7ߴ�^^�??�Qʯ����_���w���/���;w��硸�HY��Ԅ��:�����[7��8���6���X�n�wf��t�II-����d�������[�^{C]�=s~�m�ؽ���vԛ�߳���T��ĉ{C}}�}Y;.{���D�������jٰn�D]*�nolhH�	;7BX;.����52�N9��X۽�x�g�����YGE�P�yK{{;�|^ڻ�曻>w���i�'.VS�vq�V�w?�U(?���$���>���χ_�y�������O��$~�$�L��-L���꒰������ۓ�jRۃ�-�UQq	^>�[��B�<�ob��S�Cs��!��P�B�б(�/ӥ��?�S�՚���5�Kꅪ�]`���ؖ4�=Ffc��=7�o��F?~�=�M�DA���]�&Ϙ����5B!Z:���vnݎ};w�<�����q�W�fnO����z�>�hjצ�'�ڵݝk��a01 ˬ���VN��vjz�4��x�D	���E(Y�A�ԮNc�U@Me�Ls�D!V���Q�h��D�`%�����*��vaa!V�Z���zlݺ��~�4����k�~��t���#8������a�СhinAcC�b�غ$�qc�~fӆz���|�E[��ܬ�M��O�e����mm�kO<9vh"���"�Q���v��ܺ����[��wb�M����l������ar>sƅ�s;{��{�޳u#��}%?~apW���3��kMv���Hji��õ%������;���?݈�w񹓗��Z�\�쵋���=�����w�Z���{ޭ�����M|Nn��9�?�8�����}v�X�"T�J�� KaH&TS۵U*QJL�F�c���dz;!��ۨoj�/��!�7Y8��'�@sm�i�gY�gm(����
h�?G��dwy�P�v�!�]yN+qfO0��y��q�m����/��2� ���������EO�?��뵧SG=v�0j*�0a�d��(�DHʉ#���n������D�o���߽��o��Wj"A��|�	�Ų����c�9>�PD�د߽�Ջ0��OzyO�����OIQQ�k��s�}�W�N��D�������������կ~Uw�\&�۽4�[݆�^h��YR7��e�Xj�gY���ܮ���aHq�3d^-���؇w��͝83l,
�*t"U�wm���堚��$��*B$�=�S�Z"�T*�����5k��������S�8�i�&��!T	����ɛ_�]��߽��[���Y��`�ĉ=v,����e~�:�|\dy]m-�M+e�Xm�ߵ3����_����������ʏK�5cƍ���:|���%��uu5vL��zj����/�W>뇍�r,\x�F�k>Z�2����7ld��m��-��Ò%}�����Ү��\"�Ю�w/>oR�!.��;0d�?mW;:�1x�Ю��/�����.���ڃ�[�)�^�
%~}��y������]|�t�������Į��"@���d���0���5"��X�����^�Ҷ���^2d6���N!��FN�4*��B�ۼq����S�3�ݟS���X��������o��ѥd5C�*\��n�R��\��]�Q�K�9�-����{�Euu5�}�]K��K���������kW�~�ڿ�϶O�`��0i�d��=h�����oȫS���e����j���(��p�|�o�]h��ί����]�ep�h~����&�����3�o>�D���طk�'�Cu��v��{�ﺡ_��<S�u�K.�w�u�'`��9����)|X�0��6�ai뇪��X;������A��Y�Pch�.���Û���e�xH�w�+o�IC�\_�`l�ލBUlL@�r0'�N"�*X�q�v0]BS:�.�H�|�'��ɓ'A��J���#K3fʹ��sS�u��s���c2٦U�sdp��ɍ�V��vƆ��c�پ,�ȅ��S��/���a��zeBw~�qq�Ѧ������{�1̛7/#��~������Gj\��='�&�P%K_�����4wM�BP�jдŠ$�]��=,9(RB!���:UB��Զt�a�X՗'��w�Fh�j�ܕZa4�],�u��j�9�5��녑e=�ޗ
7�)�Wy��X�۶mK�_�W���j&~���ӹ��������cJ(Va�?)ڂ����/~����������p ��������������}��w�����w�~���`,��멯���|���՞�[=?��6�1�~�����z�j�������L�3Ʊ���3l�ޞ�vhLmO��9����kK&w]�1�t܉�W�g�FL쪩]�~P"T��wE�Jh9h����^5�kJ����w~E���D\�R�%F����jf7��6m�br��{���B���[���E�(�ŗ^��b��Rn�����F94���=0���-�Ӝ�niG�&�ݹ�&8}_9����8[�e�F���oc�ݱ�>�奸�i����])�8}�}��.��ߦws"�v�H�
O	I�a��v�@%�Zs�����TA3�*:=�?g�)RB!���&���!��~�>�-�����>��$K;��5�Xj-Q��Y��Ko�LE�P���Y0�nK=��ne~���x��'���!Z��N+uC�C͘3˓dVB!�I::>��͔)S����[�n�'�����YV7ԇb�������X8�y��I-Q���2���3q ��wN6��2t�j*�,��'��Jd�?کN����U\�
�?��63����E����+�����f׶8PV��.�g͙�{ι)5�f_��d�M�fa;�ou�W&rٸ��M�ĥc���LHm�tL&vlη�Z�0��؞Y�"Ŧ�?Dc}�!�o��V�x�aV�D��R��A�J�ޮ����������JLK���'�!��^Ms�>B!���,�5�'��j���&�='����푀�x0V�T�'j�T硽v�h�ᰶ~hnrWɶZ�1c��SO��;�Du�w鬤g"��vE;@���\4�Bz7"�}�����6l�r�8r�Ȍ�����iq{?�uCՖ�։��u�X&�C�#�v(���t�vc����y��x�?��,����N2��+B�e�`47�%��R�c����]�Ȑ��.P�c�0�T�ct/���Pv�/��2�t�����?!2Z����__ā�r\t٧Ч��k�̾��_��fa��{��[v�;}����.h�ؚ9���;1�{eX���[:�.|7�	���wM�r�-��k_��o	M~�^���aӇ�{���P�Mk�	U]���B���h�̿{B!�7��ƛ�!�xKus'����ri �Hs7���X�I�w�#!�=Z/D�(�cuM#:�ZgT��Sk �ZK�1c���):�577�#�����k1���5.��	!�":>�ٱ{��dj;1E$�?���J�{&��Q����6����X74N���ꆲ0,i�0��0�7����*j��4���ლ���WI[P[��IdHl;�(V	T�K��������YKd�$�������,N�>����74�S��ڍ�r,���_�0�ɚ��d��]���3�[k��J����X��+���m���9�����	�������c�ؿu�u $W\qV�X�ܮ�|-~M�<�d�L��`4��MR�թ\��TRڃ&	Ʉ��`%�����DWB!������{B!���� n�<�u5�za�a�N���`,s���8�%�#�n��XV��=�\�Y�F��,��1"���;v����X�t	B!���&���W�����Ĝ��B<��#�?~F��3����J���Jr{b�3��9Yr{Bz��9�t�!��*�>���dG�C�=y<B���S��G�D��0%7�dSm�{\�
 2Dk.	@fr�᷁=���'��z�����������ގ�־���wⲫ���a�Ƹ��nѰ�Yj��͚���:6`\�Ny&�a�S�����u\�n�����a��voiin����p������$cٲeX�z�"Ve���Ix=���Pe�ª�=�<�]�b�3�b0
�[����1�3d^-�ٍB�Z�Y�"���U������V�0!�=����cm'�$)����	D��\�gc�{���/GUU~��S�%�����W�b�䉘�x��1�BH�D�@�����@SS1C�������K2�>���c�����>S��k�C����P����ܜ\�}BxB �)4�����!�4~Z�MM��$U�R1�*�R�܍b��^�\�Ҧ�k��[�N�W$r�}�ݨ����/�B�q��	����a�ًp��磠�@Y.�H��W�{�Z�x{f�$�u+cM���2��-����nB��ku~#�Cýt���uK�E�7U�ۏ���)���b�x��PZZ�"��x7��4�Am1�1�*�T��)z�*3�u	R�J�4�b�_P�7��"!��t��O!$=�h�}�x��V���k�j�0jn7���v��l냱������ֺ?���f�.����466◿�%Iơ�8u�$�,���&�BH��P�l��	�Z��ERr�w��n�vm�+2�Ψ�@2S{�$K��k���ڡ�n��c�C�L:?�@k�ɨ�bHq�IF!ğ������r"�~��ܞ�"w�M��T|��փ�yDl#*X�q��`*�)L�ݙ���W:�����o��d���'6�l�~\z��?Q&ZY3�:6���uh��gvjV�6�;����1܇-��oמ�ܡa��8��Non����>aܤ�&x�=��N�7����Xa֬Y���A�e�A=M��H�{��d����Θ@����a"T�.�����B!�dy�9 �B�����e����IjpO��D�9�wM`���] ��D녝b��Z/T-2�NЛC��!~����wp����3�[��֖l\��U`��g�o�~ ���45���n@剓 $������(�V�I׼�b�Z/t��Z�Ϋu���Iz�����ax���v�4���C$24���Z�*�U�����.��VF�*jt�<9ֈ�b-�!��f����X�fZZZ���T4�����#&N���.���ڀ��l?�M�VM�^��XwL��q�o.��/���kej���*�\`�W��,�xG{{;vmݎ�=��{&�?~<�|�I><#��~`��vui�.%S�*�@��"�v�P�
T��Z�W�hn'�B����|B!�Bc�U���iP�G��`n���a�v���?�L����Ѯ�j�PS7��]0Vo�+
�������܌���/ $�'O��_�Ysgc�Y3,�!��q�w�.�پS9w"�
��r����&|�gBm�����y}0Vb�g��]�ʦ��>��X)j�2s{^׵�ۧD�~����d$o�)��T{�R"�V�R���=�⮊U�&w񝠊LF�J����6��4u����Z2APJ�|߾}����������A��W���CX�d1�,]���x�c��X�\{fa�fe��v}>�c�1�;�?��p篵G����O�9�Oc�ݱ����`Yvlފ��6b��#G�駟VL� 8e¼9�B��؞L����#˂��`t�^�2
Vf�����|0�B�.�YR ��^��B�<��m�c�C����eqC��6F��.P��S%�=�^����j�^��熁]K����������T��֮]BR������T�/���a�� ���8z[6|��3g@�U���Z�s�=�ya&����ߞ��.��l|���[�Mo%�
��Fs����}�����X�]�F����%X�7/��`��`0&E����F�{�!0N���ӸȤMo��,'S�#�����z
=��m�B� N�6~���܅>u	�͘��W��S�u��Cs���ꉉܡ��޾`�U�S��������8����?7��l�߆u۽��T%�l؄��:bq����ӧOO�8�&��R%0Ȧ֓�5˂���Xr{�ւ&BU(ԁ���d�AB!$�`�;!�?Xw�7O��S�k�Zs�����e	��j��!�`�Ȑ�F�e1�|���?�0Z[[����+45���7�Q���^�Ҿ� ��g�e��8y�8�ç>�)<��(((�S��x�j��ݮ�qs{0I�дv(3�w��a�g�4������'����2t$Id�&1hS�uFw��=�� �M��b��*Nz������c1b{�1���C�@�U�.�^���`��	���K0h�`e9S����D�v�f�����X{&r�&zc�֏�����{�4�`��-8T~ �إ��T��3w�\WM�~Mn���Pe.N��������v!P�+��B����<;�hn'�B���B�	!����#��dP�r}����ż4�]ol��H��x=���YL�`,��]��;@3+�|�>}�f��\�6l !Vi�������S1{�<����B!�B�o�۹{��T΍�Ò%K��KJJ2�p�	����$��$ݞ��w}�P��������;L��E�x�H>��g�6<�'͆c�i�h�ԜH�)Z�"UL�
h�+��]�� ����U���"ȉJU.�쮁�O}w�;~�x%�S��9y�$������>�y�`�ҥ(*)���Ooj�4]ܡa=#L�����3�1��X{�{����eq��X��4�{�*N��z���L�Aqq1�x�	�w�y�o2APJ��;	�*��=>Ml/��خM`0�����?����'U�B!�ҿ��B�4��q�1<X&OpOR3T��j��Z7Tky�:!b�X�r�l���j�PS7��o0VO�8p��%j��w�!VZX��8~�(�.^�1�ǁB���@,�%��˜9s��O���Q���ym �6+�1�ǌ횺�ݮ�AC�0h��Y�vDk�ښ�:�`�ژ�N��w��|� W+FG[��؞��`�^�JLq_�JkrH�*�4���$���w��Ϙ1?���p�}��ĉ ��k�Ə�s�v,X���,A^A^��[4�{dl�l��e"�s��e��a	{&r���vƆ���!��{�Ą��Xb�{=v��}��MM �;��GŅ^h�$�X�ռ��@�.��+�F�T���"���Ik�L�jz�Y�����#�L�Ǎ�
��B!$[ط�B�_l>с��Ek���@,Y�P_3L��9��92�k��`,h�2�қ`,;5F�p�>O?��br///!v:�����C0w�BeJ!�]��N+����*�f͚���2$m��t���=^34>:�?���ܩ��������5�Ȳ�O�hn'�A�;�xZ::�?8cC�ʇ�,��htכ޵-�)��P���U@��`$`1u�A�e��	M�`TwSH���̙3�ar���0�O{{;>Z�>vmێ��/ǌY3��s[&r�f]�fa�fe�խ��0�;4�[ܗ=ý�qfcәz.ݦG7789&��~��.��f*O�ĶM�QW[B�K~~��V���.�,2e��ӻ�m��d	��vm�*X��0$�T�V�b�s�D����B�f��蝼4#��/��gF�A{kK�F$�j��j�P��	&w��'��f�Xq �eٝ`,;v?�n�رc�`�{ｗ&w�-���W�b̄q��p>����B�3�MD;�lS��	�.S�Nŏ~�#�9�3C��5?�ǥ5�k�>���±��:��%ʺ>��]��V����Gqi_��@. 
��;hp'=��:0y�8��>��nP���UZ�*'n�7��L��/�݅��S�7i�AU�Q�<�&�L�D���Ǹ���Q]]B�CcC#־�
�oނ�/�#F����p홅���7�{a��s\޼V��[��L������?��8u��aℼ�<<����k�
=�`2�{�nC�%s�>�!���O_P~N��`��BU߁���;B!�d'"��K�-Ŀ���B���]m�01T�܌�P7�>;>[��2�
�S%K������̞	u�t�Ǎ����TQQB��й�>�Iӧbּ9�/( !�{t��cώ]ؿkO�7EHw������3fL�0��a����%c��~���C(V�wy0����ʼ!K�-���<!co����^.���MMq�J���A�$wm�{N ��x��>��*m*�����tu{�pf�N�����?�r��0���׃��r��	����)ӧa���0p����c�3�ݑa�5��Dڞ�<��ƙ�������;iin��m�q����q�0�?���4�[�7۝&0��e��v%���ԞL�����ە���!����ۮ[�la�ޣ�`�!����߸B��-;�_XEqa>!�d/{���:e<�Շ�����f�7�'����fh��R܍Y1�ciɄ��߆�I�&)ݟE���#G@Hw�X��8\qg͛�IӦ*��B�#>?E�p疭hkm!N7/��:1�C{wM喙>'��	�R�V�>w�:���s9�'`_9���{hp'=��N`S�P��iR>4#�
9	�2�{d^/P���`�&���U����h1�ir�c�x�b%�A�hr'N)ۻ���c���X�|���{ީמ�ٙa���{G����Z6�{`7k˰nq��1Lv�	ݫ�����ػc�"��sB�"η��s�!�鎹=~�]\�R���L�jZ�i�n�T��&���"!�8A��ʧ�-tt}�|�'��7��}���_�	�~�Y�w����_��&�!������N\?�?Z�u�B5+Y���n�} ��]�����h���ac�Ygʔ)J��=�܃�Ǐ�����ֆ->F����1w�M��z"!�d�{�ء#ؾy�π������z
'N�V�/��������N��$5�d�Xj�0���I��]���X���
�8Hz����(�1u��Ք'��V�X%����8���9�J�v0�� �"w���I��t��V^�IB֒%K���+W����8A����Y��b΂y(--�-���t�|�d�S����N�
Lm�w#��X�����W����m��Q��}س}�bZ%�rss�b�
�r�-i���%@�"q�=�*uCb{A��`0�b0��U�*jr�J�����in'�b���\<�����O��W?�ɽ�Q�ؒr��#���_��t"n�����N�4�BH�'��ځ8��L$A0Z+�e���؀��YMs7� -P�S�!jk��`,��.��Q�JT�զ�g��]K�u�M����E�g�܉S�q�طs7fΙ�1ƁBH��'���ͨ��!n0b�<����M�=��翹=;C_?�����5Ci�g]8�y0VB�g5���i}����1�Iz����8^���#�T{*!�!���vP�̠m9�#��9�85���b�A���"�6�]��={�Ťt����ҥK��U�V����8E�mo��	��맜|�_��Iױ��,kbVv`nwj"��Z�]Im��/k�쌵g"w�n:֖a��X�7b���:S��Cm'�k�v���6�ban��������7ڻ{�^'0����*��bP+RE�������B������oƷ�<^�hH���܊o]�3�K:�W-��������]��Kp�˒�y��x��� !����Dc'��GIC��(7�Kñr��Xڟ�5C���`,�SM0V$K��J�{�:�v~�̙x��q�����
�8������w���D�n��Nc�'[Pu����0���'?��3,��2��矹]�q�E��$]�Շ��vyb0��n���b��>w��t
�W1L���I��#E�lh1:�ڢTb�A�@��7Ot7�1���@6U�ʌ�q�B�v�س�@FK^��.� ?��z�j&��'g�� [�.�.Y�9�梠Pot7{�[7;5+����Dn��k[4��7܇-����ü#s����-ý�qf��	��mX���]c��r��EsSqq���_��=3��[hr2/O`�$.$����`��)D��D�Ǳ�iڃL` ��}���W܌���Oi3A�tt�K|�g�c�3�FQ�y	A�����bǁ�8|���cz�㮛�'#��>�<:B� ��=�{8����FK��x��f���.ꆱ4�@@7�ĊeɃ�T�;ľ�Bc0V�t@�	�f����E&��gϞ��E�{uu5qa�lmnAmMf/����B�����ؼ��� !n2r�H��>k֬�4����n�.Q녩ñ��v�`,IH���Ϛp�����J��$���Nz$g�;�?8�:+�mL��y�@��"�H�;���@�ʀ�(�R�úm�m`�û�e˖)�=�M��UDz��＇�?܀y�b�����ݳ�v��iJm�gwf�wÄ.]�����n��L6�Jj�a��QzeX��=��;�8z�0��؍3�� �mĹ�+��/|�Ss�ߦt�捩��H*��v{	r�J���T�����.��&����vB!�����/��}�y���n�����U��o��Ƿ^�t܀�"<��-���ߢ�ݛs���"����I���N!�͋�}���"��lV/���1�����������Y���x�~���?�ɔz��ǔj������<� *+�2K����c�c�ј5B魈.����у�A�ۨ��~�ۓ�W�P�&�hl7Io7Ȓ�u�X��a�@,Ӯ�Qs{QI�t0I3�x�ǲ�T&L���Cq� Z%3�'$o;(0
V�w�f02,����{��ݎ��t[�{��ʰr�J��y�E����6l��>Q���-@aA<���,l\�Ԭlc�w&�L4�;�8�ܮ����.��9߳�v�64����P=r��v�Qn���M^^|�A�x㍮�ۍ�mJwk^���x
�F��el��.�$0���*������c9��B�C��u�͸������3x��MX>w�9ﬤ��N���~��_�ۗx�}�B��������BH[0���C1-|P��5��ljv�	Ħ9ڟj�F�{��]�cA�����fBݯ;��t��Ν���E0ֱc�@����N�ʹ����w���N<c��ъ�묳�J��݈�uA+�zc���.��Sw~6�
F:=�u�P4 +dRC4��,�ak��.�I�����h^��������Z#B�[�	V9:�*� V%��b�1�]��F�X*�X7.��{o2�kq[�:�s�ӟ�T��z�xA����f,<{fϟ�$�'`��n��끉<�؀a\��lӥ�s+���zps���7녹�+�<1���<�@Y9�l߅��f����/���W��n��W�(��{=���ęU�������Tg��P0h*Pi�j*�(,*�ߏ�	��^Zۃ�#(��EIQ���N�4�� _I�����?�u}��T'��~H�����7��>~����n�h[ڰꗯ(�8n R�����I���N!D��:�)�ǣ�����sN�4�d�H��1�]npW�\�`��~���y&w;�t7k�"��g�Q�܏9B�Fkt?k�L�;!��&��VU���	�x����s��i�|1�gB���v5��v}�c�C��Za(	��Χ�ʻ>Ob�g�4���0��}�KK�TY��*P��D�J+\A3/o;���݅9��.�H�q@k�Ӧ�G~O���3S�J��%{nѢE�`%�B�z�xE[k+>xo=>ް���ż�PRZ�Jj�U#�w&r���S�}u����wj���rhηe���ƄNs{z�>��+�w�0���/),,�#�<�����U����N��V���I�Z��?Sۍ	:s��H��;$U�����6�T��n���w��/�G& Һ���)ǉ�{�o�w�M�q�d-��)����z\~�4�:y�9��{nT�_�g�N�̧���������@QA�r��?�W.��vҜ��;v؀�chn'�b���N�2y�j+����Qc��!��}h���=G[/��]SY0V$K���&w-^��O��c	����L�%ޠ�G���sgc��� ���Bu�i�پS�����x�ĉ���'ONKMЈ�fu���0,Ӯ�����e'�]]�a5)�J-1U�gY��!���2v�'�A�;��T5�pr�Xj+3Mq7
TV�*y��ؼؗI*Cm�����t���y�#ar?u����v|�a���>c�Y��x!�W�������s{�|k�1ۗ����������n�Dnzs�l}�XK���7������!�|�~�߽�� �k����f�\y�=�ܞ��TI��p�Zv��Z�d)�;h"����N!$5w��_�Ζ
�n�-�oj�W��/<�K�Γ���܅n���v�d>�+N���7�+nH9v��H4�B1��%�h@�r���fh�^7�[�j��z�1Kot�&w7넩�%B���Q1������8v���2l(��>KIv'��L���
{v��	�S�*��&LH���o���y�f�7��S�e�X�k������
:���ϯ�㩿�����
6��SƢ���i"C���wS�;�r�$�AO<�A]7b��2\��=7w�ܘ`u��Q�%��o���c�X�d1��8Іa�y&�a�u��pj7kٰ.]����2gϠl�^�W�|F����s�W\��B������ԈT���!s�J+LY0�ǒ�%)����
B!���;ۻ�K������߽���<��OI����V܀����m ���]��c��Ǫ/]�����N!$)u-!0
Ãe)k�v��j���]��Y�*)��h0VB���jlW�[�N�/���4�O�8QIr�X���!^r��
��|G	Ě:k�Mԛ�!�/�w��cǱ{�Ԝ�!�@t��cǎMKM����0A��Y���!Z��v���h�0�P;4�ծύ��L|�w�kx�"׍폖3�1I�n0���`�vИ�)�iE*�pe��5�DЦ��7��H&�C�܌3���z��I�(߷_y�?�/���l����~�O��f��3֩�ܙaݖ�܃�\1�K��oB��=}�V��w�Q�b��$�_�~x���q�d���ܘ�S�O��0H�Z�E���ݮ�]��`La����ۧ"��3�B��_X�֎ ���������N�����4���ן֡��߿i�o���wᶟ�@s;!���l>�uS&�����f�c����������5Cm�PE1�#^/�w��MF�����3�Nh����0a�y��\��v�!^SW[���>���1e�tL�:��� ��t#jGR��gAH��9s���>f���xF�c>�}0���.Mo�P7L��Tj�A��v]r�!�=g�$l-��������	���������Pe�� �?��Z01�!�t�9�w5�!2&"�DZ*si7��axw��.�܅`�o�>�.�:�<DB��ys0c�,�(����v{���p���Im�n��e�:���n�po:�_�:��CM\�EKAB�������SO���v,JqSd��Ю�W�)��].Ti��*�H��TJr�=s�Q�R��b��P��B!�m~���PR�o��-L�:e�_on�|~�oo(S?L�"���vB!Vy�<�'BsC��f��J��n��ꂑ4wm�P<dI��pT�b1,.��7�H:���:"9T��V�^�m�x�$I���c��]�2s&M����BB�״���B���ݏ��V�N,X����1b����tڽ��S��I��G���#?%��!������ϥ���r�<Hf@�;�U�h�x���T�,�4[�}���P��� ��RD,$���S""��j����=��[�L�8?����裏b��ݰ���^�_�Ȑ����}��/����/Ӈ�݋��n�vqb����رe��<


�4Jm�mhmnQa�/����@юL�������K�HuHb�¤kwg�_��Ȗ�߻��MҒ͎������^�{���ֶk�B����ZT��oe��mZ��L���=?h�������[�345�Q.
��ٵn}]]�{�F�����������~~ר�t~���گJ�wQ7>|�r�5{�l���q�"ju_�R���ZIo�	VR�J1�����O`��O�hn'��"��_�"�q�y�����{WaK�q��G�܋
��k�I�>��N!�.����+�ci����X34v�R+LU34�
��X���`d�z�|zM��zQ'�Ώ=ZIr�ᇱa��.Z[Z�㓭صe;�N�ig�D��@!nS_[���p���rBH�Y�l{�14ȳ�^wֱ�]��!��k�� \��j�0E(�xN���R~��ۃ!��X��aA~>^?Q�u=E�d4��^Ǧc�v�xt���B2$���%�OhD������dE�RS�)�P��Qѩjt(_d���v7'�ūQ�F�駟VX�֭�T�W{{;�@��kէO455�����b�����W�����br�N����c���	f�ƆT�>��&ꖛ{O%&r;�p��;wc���}���t_�Ǌ�QO����Im�.��:�|.>�z�y��k5Mm�"��M��X7X���?���M1ۢ-�ݱU'O����O�R��0�O�:ٗ}��SG�c����i�o��={#�T�Y����������[+����ɼէ�
?_��������a�ԩ%J9]�+,�6e����zc���	T����`4��O����k$�B�����9~>�P~}"t�A�J@zk~�w��𭫗x�/��	!�t������)�?�1��5ø�]�hpW��S������jz��{_�g/�2d~���'���~�-Q��
�;��p*?�R��M�i|X��K�1p�`���k�+�P,A]M-���ǀ ��/�kk��RX�]�kp� ̎�MMhok�e��&���v��3���]����[�練�������x�
D�.�����~�
��-�X˗/W�唖�zV���:�fh�����O�w~քbj��S�������ۃ�������	�ma0�hp'�����i�`45�F��I�)� �A�BJLd0�S���F#�Ơ���v�����='�-p�c�ڵ ��{rߞ��cА��9kf̞�u��P����[2پ����Ec�sý��`q����f5��e"�e��3֡�^:�}úW&x�}�<v�w�E剓 �ofΜ���Ǎ�(e�?�z������v�Im�br׊R�H�.����w�e��`x�"�k�K���F1һ7| &����f�8��߯��8g�8e~�#hmwv�!�������m��y��U�{��տz��TaΤ����t]���w��{x�B!�{l?с�J0��x�Ϥf�c������;�k��iL'HHqWuUu���Yݟ��V�q���S�E�z�)���˰BQQ�����g0�x��_KK�/��;,ī�����S����~H�&MH08
��`��A�?�������%�}|�����o�L�J8ըqc|�����1b�(��tS���;aN�����<3���J�P5�;��~�Z�� �>� �k��ʕ+�s&/k�n����)��Wk�zc�$K��9U8V�`,%KIp77�kk�f����8;*hn'��W"��=�l�����Z������[�փ��t)�5��p¶R�n�ʭ}�5N�??����U�򗿀?�9]��＋M~�ig���ٳt) �M�f�p���������>ֱ1��ذ�����5,��?�7���nѶT$���݇��f�	,\�P�ap��ᾋR�Yǩ�ݙH�OmW1ڭ	TZc�^���/%���)��U������V�T�wq�����7�oI�F�?؍5�Y�cU��D.Y8O}�JL)h�>T�����n��靈����X0u4H��w�~B!$�y�<��'CSmUb��]c;��CM�;��c�t�h��R7�uYqTc{d^����v��v���5k�(]�_x����7Dw��mĎO�`���4}*B1���������v0����?�y�X�B�Q+Sk�F�7��KL�>'Io7�!&�
�܃��ꆚ�a���c&H�A�;�Եvb�(��<�|(���bL�����Fw��] �'��6�|�i�ܭ%2$#BV&�܅P%�-q��?���񝶶6l߼Uy1�ƌ��c%w�;5����%��7����Dn��ō�2��2����p/�	��v��'��Q���U.:	��-[���]���:~	\qaJ�,ǖwjR�%$/�甶�Am�AU�
�No�̫bUp�$�b�e��Ogn|f�L\0o�]�[�<�I|��%x�[WB�Q5s�0��W�;?��l�s�wB!�������b\1��m��ρ�4�d�CH����XO4ܣ(ݟ%i�q��B���0��Q'���Hk}������~�;�'B���W�<��S�`������!�tv�8?rL���3�$�����{��r���2�&�t}o��.ϒ���>�=Y�0e0��Ƃ����=duC�(*.��G���UC�o��Nz5;N1v�xt�ԋPI�)�p�D���-�F�2��(V))��id�jt�orO&�h�$�Jy�.�G�5x�]w)���}�Y�)���B}]v�؉�fb��4d����V�E�'�'�NM�Lm7�=Sۉ�3�gp�� �U���t�ȸꪫ�j�*%��M���8��(#n�TZaJ�b� P�����FD*5�!"P�-CJ�{|Y�ʤ�`�����r�n�%���י�U�u-�6fH���L	����уAHo��x5!�B���-��#0��@��s `�t����;�6��?��v�x�+쐰)Ф(�B��=K

m�(P6!�UF_(e�Zx�{�@�jl'�^v�x˒��邏�Nw��>Yϧ=t����$ǖN����~��.���.�r����z�\�Rc���,�ǨkkVHu�{FF�=�\��}����7"$��t���#??���M��((*!$��ڵE��K{k�t]B�]���wu�	'H�J�T���H�z���js���5������ĶөNm7��,�d���a|3X5�y��EĞ��NF=�Z�qt��q�zC��l�W�BZ���G�R��*훟^��xc�\����G�h��=�w�#���>UUU��[�p8@�]�7_}--��J�ݎ;`�v� '7W�o�Dn�ֹ��#Rzhc�o46V��ǆdX�8��qY} z�&ڰNc�9"ma��.���2m�ؚc�=�w�����fn���%�Sjc�B��S�������*c�,X�*Y�r���z������6�#������� �.�BC�NB!�$��nr����m�n���Ak��-��;?�F)�J�{���9��+6f�D�詧�*%��~��� ��U�W�R�k&Jan���ːckV�B{�2��-��͕��~��1�Z�:��j���v�H�۵�X�����r9�����⚤��	��4��B�;I	���Ay������-�He0���*�H%�*���5�GSp��������xΜ97n���Zlٲ�؍�M����ه������v�v��ﯲ%�Es{�l�&�P�F�0��s������P��sń�:��ƈ����eXٶ\*�����;"���:�,��`�[Zm!+ZsY�<��T�R{Au�'�����ss�6yA^ă����CNB!��	�BI4o��0�y�;ש뀊��1���������u�:�ۛ����,cy�%O��x�8�s<�cPYY�����5Cb;�T�o��
�k��8��@������X�b%ּ��bG���p�Wbƌ1�Zs��Hj�ʚ�|�.�U�X�Zb8�}�X:�C���ҭN�P����k��R�.{C�;I	z�����b���`e*PV�m`*���J���Ms����F�cl���]�]M����փ�_~96l�W;zBd�貖Vi)(,@�6۠a�f�W�������O�z�&���uǆdX�8.���s��	=&�T�gk7V,[.-b] ރr����w��K/�!��ւV��UȲz>�ߢ��L��k/(�	�In)�3��R�v���BO�H`�HE!$��ݴ'r�(KB!$q��<��/�@_o�B�АC���v~�� /ݣY�k�R������E��?ۥ��qӧO�m��&�׭cj.�B��b)(,���F�75 7/��䣷��m�280����ۉm����u�]�)S�Ĵ>hu\<j�њ�_/������ImW������|Fv���nnn�j�y#�/�e��aC�-`%��-.T�5����/@� X
�J)X��ƕ�MeP
Wfo��4w(�*��M�b]�	��EOd����cB�������e�]��K��;��݃%_-��¢"4o���n;���-]F���i��9>&x��qKm7k�1Li��v�0�=|�����#4oڰ�$eee�ꪫ���Zq�����]ml4��R��U��v��@��\N�}����J��A�sB!�G�G�X��Ԗ�B!$Q:��bk�f�y��B4����c��=�=�����I�}j�A���)�rh�/�@�Sit���]�Us�ո]w�,�j�--- Į�tw㻯���K�Eiyj��P[_��lB�ːÁ5�V��u6���J��	�+;�#���?a�ĉa����E����KknW��C�P,�ڡ?+0�%�`��X.��v��azF:>��!�0�;|%)Ň+�0{�D86��ܮ�` ZiR�I���u�X�V�T��<���4���(�����p�B��Β%K@H2нu+���KiWV��m&�y�IRjS�Ck�𘥶�-�38U��4���E)aj_�f��!��d�n�V���x���^j�����`)}A��`�^Л�>r�?��X�r*��}%�x��B�mX��wB!�$�[\���GY_��g�1#��%hQY3�z�6�][s�Q��)�B��f�X������<O?zsk�4i��\q�����A����"dG,�|��U���Ԁ��Zdd��C���ڕ��޶��C�t�@,�*//�g�/�u�X���vm�0�P,�`,�v������N�E̵&s"�v3�$��%)ǫ-i8��}[:B���o[���\y���c��B�ʠ��'�*�փj��ԂM���UTTছn���_����$��:���O>Cye&66�q�fz���10��*�=n��n��ذnql��|��z�ƎV���NFF��T7�k1�����-m��"}a�zr�����S���z�vi�SJ�{VN�\W��B!�.���!�B��b�f5�c��=�.h1(K��[3���:���ʘi�w����1�����B�[�|��u��7��k���B��;,�Ų$�KL��Am�DT���|���!4~Q7\Ѷ\
�FSB���3g���/GAA���V�%��.�c`n�	�r[�k���c��vhhn7Jpr�=��[��E��I��y����<X����J��nx�O����4�X�Oe�o�I"��X��V�9z���+紛x�1�X
V��ŒX%�>��3 $ِīu�勏?���'5���	E%Ŋq�G��Je6N�=��qFc�����c��n��ݛh�z����X�zM�d�0m�4)����4,q�l�h0����򺜾�m+,�A?�]���i/('0i1h R	��BW?E*B!�b�Z�	!�b^ku��*�u���C���5��!������2�u)����%5�x�+**�7܀;��=�I&���޶LZ233QY=�k�Q]W��Z���#o��׮ê�X�r�����d���y睇��,[��=&�㭝�_Ԛ��B���cik��`,o(��klw��U�v��aA�x<�B�I.xuKR���n|�W��ۥp]A*�p��U��,V	dQ)M��}:��JNv����j�{�D�h��q�O�`_NN�ϟ�	&`��;!Ɋ2ٽ���M�k���q�����c��nuRc�}�&���Fj��?{LL�LmNOw։�����ظ1ed�1g�\p����K2�O�*��#��/LI[P�����e
��8e�ܮm-�Kp7I`P�/hD*�s[�к�׺�B��'߷�p�ٙ���#�k6mIr�2p繇c�m�a'����7����@�G]e�GG'}�l��!���<��b��ǴF(п߬f�4��������r0t�?�!�z�@]���=�Z^(��D�����/DYY��>����Dh�"�G,��?��k�뤄wa~'���0���9�Ծb�/X��dE\��{�8��c�^��j{f�en���]��6��ە�XnˡXz���ڡ���:uk��.����C�+,�K#�{I6hp')˲�NT�L���V]1*����m�4����܁�7�1
C�R����^�M��2����l���O<uuu��k���B������E��s��P�0�#���jT�}�V��0�GhX�:�;����o�T	7����[<߮��X�j��l�`�$]�k�y���SNAzzzL�'�s�K���\������j��G��On�����U"��e��n�d�����	!�ؓ�Vlĉ���^r��1�p���^ŏ+6���ń'.�5�Mi�y��0��'��+A�AfF:���8�gۃ�Y�ُ8�ƿ�bF>B�����K_"V#���v~V��KrW�jס������v{��k�ꚡ�h��U'�w�Phg��~:���q��ף��_>"ɋ�庇�ݮ���	���mvN!�����DJ;;=�ф�^s饗b�̙Q���K�Q=�c��+���._��bOm7KnW�إ��r����v����>Q;��sNI6hp')ͧ��8��C�jJ�zPF_��jS^�
aK��.��
V����Oq��*2���.�����*U�NBT4+y{���X�`���J������B_~��i����rm�D���kF[7����n5���o�	>$úű����n�\����p8ذf6�[�5+Wa� ��Fd�ꗿ���K�~� PE{\,����v�X5�M\P%2�ۇu�)��]���t��+���:K��2<�*>Q�p�B�	�^� �4����C�~�4���l.�۹v%+3g��6��3Es;!$)X�Չ��ZT-�s����4c����.���P3Ԇcy����n�S�w�ۃciI�:a(��QO<�����Ϣf�b�
���q����"(*)���jL��W&B��֮-�/�lڰ��6jkkq��bʔ)q�Z��N�v-�ڡ:�s?�uCM(V���q0�6K�jk��±��� �k�م�$'4�����a�T��΍~Qʤ��@u_��� h[z��i��e��PR�;�b�[ό�ڡ��nr�Q��<y2.\����
_�5m�٭[����>����QZV�ꉵ���AyU�d�Wb��n4������>Xk��,�M�a}�����ذ�׮�:7u���LHUU.��2L�:5*�پx���=&������v� ���D*���/Py�+e��^��P�kn�?'/o�.y<L�!�b��o���n��ogs�?�ً�4�B��o�:1�i"�|u7+FwM0X�л#���B@��?'��]�Ь�w��W3\�d	M�X~���())AgG�dx/���2�z����v��[�FJm'd���{H�6�|v�ZKs�q�P���P,m�мn�2�҆b�B����N�"B ��5��6��I��+U��$�E+�0�"��}���`B����h=x*}���Ms��X%����C3�kG�ūP��<����jjj�$��n�	���:�dTӱi��|����kJiy��Q3�cǍ�1Fj"w�1�p��a=s{��{���0��jl2���#	R"�}kg�n�
BR��w�]�D;�x
Tј#��h�M��ւ�@�1�����{o���T�P5f�i|�[��A'!�B�I�ȅ��<�ڌd�o.�+7nAuy1!$YX$��&U��cm�Z�aѰf���ѕ�U�۳;����L�J�Q'�em1�8����>�pz���n�[o�BF#BOl�o���Za��T��B��RVY���dG�΋���"k���~O�hgƌ�?>
�^4�g�:b��|.��]��9�P,m0�����t�nn����j�B��$^Bl���W=��9k%����*x��r"��\���5�q�}�u��X�ǟ���=R�)�BT(iV�H����J<�� $�G>���O?Gn^���0���UU(X|46��`հ��<4ý�qF��&ڰ>ڌ�=���q�zlX�}���}��� $U�5k.�袸Tf�!J�s����MaP-r�A��ւ��԰"}����R
Q��T��6�7�}#��B�>7�y���H�oq�[�bnx�m�t�)�\�B��yyYfO(B_owj�r�P�ߚ�D��Y�v�_p���9��Dc\��D��0�766⡇u�:!J�����SZ��7+;�+QQU��	�_�ZIN��X֬Cff&zuDBF3���8��q�YgI��v�Z����q�z��X?4�2�
��w~��c���f5�`����b�cYL\.�$4�⥽˅�	Q5���]Z���vT�����e��*��8�4�!XY9o��ą��~�;)��[nA__I%���}����,�WV����U(-/Hm��z�1�plH�u�c#5��=��� �1�c�Ftl؈�k֡����2�5��3ΐ�F֎��9kn����ܮMafn7N`��/�]N_p��a��E{A�6��V��	!�}��7N>x���>�a%�uv#�8�\����؋�~X�_�T�]"��d�1�����W�������.0���=�jñ���r�g!^�[����#���پX�q�Itk�Bk�7o���q뭷bpp������U�WH����PJu/KU�.DlJOw�T?ܸ�!
/!�@nn��u���^�*�C}��h���S�������"Ky_��XN���kvW�ӫ�۳�2�r1��$?4��`�!�Ѐ�ͭH3Ɠ�` V�&'2��Fw��.��`8�g�����'��ڂ�M�b]�q����c"�C�>��={�l�����C[�H��t`����"�Uƣ���W^(X5|Gj"7����#2�GjΏ�	=&x;!>�uut�c�&tlڄM�7b�����Ÿ��q�A|��.������v�X��Z�{k]�
L`P����)�0\�����k��R�S%��dg̘��S���C!	f�]�p�)�:�1��'$�9!z\��[җ "}��َq�!{�B���n��3��e�&w����f���3���LMHr=�J�gar��e�/�j���lΜ9����j�k׮!��0�eyK��-�A�V��ld�XcKǁ�D��Z+u}&$թ����W^��w�=�B�}ў#Q�v�h��҆b����͂�ԡX�ڡ�.h��4����{�EF4�����9qDs:V��z	*b�S��%b��KRʖ��o�R"�ț���b ���c���.���eeߔ)Sp��wK-?��CB<�+�-���b��.�,az[Z��#5���jV7�8���!�{��a=���@Wg'6m��Q���7�	ѥ��W]uv�qǄ
Tf��������J�*����@�m1����HYp9-e�*��v������ ������=��w��ڎ�&`��d�wG�Bj+Jp��DzC�k؍��~��vb�s���O~�x���ੋ�^��t>;p���Ď�� �$/?lt���%=��:`�:a`��5C�����<4A��?����h��徽����w���Z,^���2���Lx���Eiy���-+��!�Dh�;:�)B�F��M�08���(�k��p�e�I&��Z�:.Z�vm��(K�*�����`,U=�gl^;42��eKa3~Z9BF��$D��G5U��s��T��R�J�������+�7Y(E*]�J�S)�x�e�z4��X	V��UUU��o�=��򗿀Ȗ�-�������,��t��Ri;N������î�bal��{�a�1��s�HU�ҹ]�G����� !$83f̐��E{d��can����ZjĩP�����~mr{0S��1���Moţ7V�9l��{B!�_Z��;	�/}��:�����/:S�ƃ�6�Y#�G�� 7��^�����؅�]�!�=�p���Nt��>Y�ġM��l�\'ԯ%��k���>��B����]{�x���2N�z�vκ�:�y睸�;��/��At�Uv�/��E��]$���,��} �9�]��E���M��N��c��y睇��<�55�v�k{ј#u�P���n���2�V%�����b9��|�Js;]��N�B�yey6�.BOw�D�Ȣ�^��g�˻\���ъU�M��f3�{��	��OolNN�9����㦛nB__!�8X�r������zM�e��U<��8����=ѩ�FccaBOVc��=�-]]����eC�0kBB#=='�t�͛�����Tf�%^��ܮ0�+D+���<�!P�2Kn7j/(��>arW,���eO��øC!$:4M(�3W����|�[�?�T����1���&r�ɿ���	A�}�t5n��� �BF;���qԤ	��X�>���fx��ݟ[�9����><����5�"\�{2���!�FͰ��@JF�f�m$��� Ӄ	�"�f�vm����e�}���R]���XZ�R�1��L����������)���#:��J�%���.��9s���h��b�Ϯu�`�ve��j(�Y0�6�ݿ�
bb7^�˪��R~��>hp'Ā'�A�8�S8 ���P�KS�������,UG���
c�,P���9!�����E��hr��>�v�a����5�\���vB�#^�6�� -J���%A�d�X��YJJP4�Y��vӖ��~wk�vC[�ű�2�'��]�����{�G��:r۳e+�n���(PTT��.���կ�A�*P���]~U0�kZ���0lA�
������ �2c"ڻ� �2�ر�/�p
�\��o��9�r2�ĥs��@��6�C�:�w����x�6IلBH�y�5�3q,��v�
--�k�i�z�<�}A�?k���Z��/�������j&�h���_��ט8q"���:�]��s���i�Fi������,E%|vv6��D���oDOw7�:;%#��)2���𨨨��W^�}��Ǵ��ݶK0sD�����ܮJm�1��c�c���=�C�3��v��XP2/��LF'��&Ą�=.��[�F,W��C� �X�6���Ղ�b.e"����6-M6��s�E+y�d�����'oO�:w�}�dr���/A����^iY�J�ʼ��P�
E�C

QP\(����&x�8Sۭ�C�{�v�Hi
==�[af�����7�������&\u�U�i��l%P��øP��򺮹ݻmM��7��t�,P)�����r��	!d43��/�x*���)���鹪���Km)���~J
rq��g��2����t�BI���7�a���dٴ@���^��$w�~�����q�F.����R�����ќ��|��gt>y{��ƽ��+��,YBHh]U$v�EIfV��I���zaq1

@�|%��[��Xb]d�I���~�	�»t��W���.�^(cen�GQ������B���:�X.ej�y�0�۳�v�����|Nq3���Nhp'$?lt���%=�*Jm`N����|��/Zi�ӛ_Nd��vЛ� ��!~�E-Zɷ�`r6� ��������]w݅�z�=�X\L����[��X��_�
�'h!7/y#�"�!g��]n��������L��}}�"��==ҿ����[f̘��/��������a������]O�ro-^{As�rqh��J밨�!�$#"�z�M�y�
�Uc����w����Z��$��o��a_Z�q�>�Qz�#��Y?�e��A�=��7x���BI5�����
�3�=�X�j��f��_3LS��60r��8&�V"b	�����h���U3��)�w�y'���?�7� !$r�iO��.���-d�����/�-��f��ė���vw�{d������&��E-�9s�����/�M%��>;��ܮ�'Z��ܝ��v�N��J�зx��c�����Jt�3��^hp'���t�Цzu.W�K�~#|��P�o��`�fl���7�+��������Oo�H%>�s�����oFg'Ӫ���P6��[��S�}
û0���`�V��fdf�9�Dvn�s�G��s���TJmY088���~i]�O��}���^���vB�A���֩����N;YYY�5���/��v�5���]��`��n����&��c�{�b"V���s��[��-!�{�v���sמ���c-#���{űx{qn}�}|��*Da����_�}v�έ}�����G߃�NƤ��].}h!��Te�f'J��c�`+���*k��BE�PB�ˋ�-Yc�e������J������'R��=�mr�Ƹx�(����p�u�a�w��@�>��Atl˦�}�Y�RmP,��y��37/ϳ^�/ൺ11F�Ɖ�܉[����W
����ꮄ���7�v���裏�y�d��vh�q��9xoC0�{;Ak�=+��5À`,�SSC�	Ͳ�%�^�Q�U[�@�h�wB,�j�s���ױF��e*�Vz�)��g+!N�$2$���q�h�Yfs��+��3g����_=����]B����,X�OCMZ�H{��͑��"R<K�d*��ʔZ ���v�ȭxM��&�1H�H�AE��.}�Y�*#��Q���!鹉u�����W�ş}A�:!I��s�E��?�y��P�&�x���B�B�@e�^Pafwi��J�IW��i/�_T���sC�r!���b}��/x�⣱�v�����k���w�F��؊����}'����A�Fާ�F>�de�?��{��F>�T�b���J����.�6v���.���翣��B!$��z�J���`\�Z/�����a���W@�PO���&�a���4���]�#i!����-Z9o4��OolFF�Ν���f��r�JB⇨�uun�=�����˗j��6(��R�07٢F��#m���ъР�җ� ,����R��>)(�uEB�ŤI�p饗bʔ)��&���1��8��]Q?�N8���~0�q�g=�z�P,����,����~F��!1���8���]�+-Z�'V�o4�}kҢ7�v[W�&�`s�aV�D��~��q�}�a��x�@I�8#�p�8cFa���"BF�3��#�+�ۥU!�9�oҪ͉��[!�mq��c�f8��RA���a�}��%�\������Nњ'�sDz�`�vY�����[k�����ւ���ZAʡ�^PY�Z_�A'_�	!d4�~s���	\u�/qƬ=�JflS[.-�d�5���6����p�AR����;���Vl!�B���\�=i"�V�X�3��y����ϊ�fݟ�Z��5�[q��8F���4��]�����n�/�j������}�������3��}B��t{{z�%77�g�#=#C��yB������Δñ���R ���c�Z�t��M��Y^<N��%���+�-��"K�';Ep�'KQ����)��}}} �$��bƌR0Vyy��ꁱؗps�X��
��v��v��v��}�5[����%�7�:��T�X�bz�D��b�剐��˝�WV���b��l����Y���X%�T~�*����.��&�{4�	�[XX��.��'O�-������ �!�yj�x}���!��!��D��9�#	���3Ϊ�= ���*P��u�yr�YCff>���~�T�2�y���7����p�y��� vd�����m����@I uX�ُ �B���[ܘ�4}�k��Bx����a�qP����0�~��uQ#T���55C�^(��&w�]�F���ت�*�z�x���q���K�!$y�%�b�A�_����7_}mx�X�V��B�����78�䓥����26��A�sDfnG@�PU7T�CKn���S�=uC]�u:?�M��K�DBR�		�'�ֆ�?nHj�$�JJ�JO�ҊW��Ei���ʠw3��d�O���.Hf���|�̣7V,�g�Fcc#�������B!$���R���P�LV��l����:�j��X���خ'L9t�)���?�j�jK��<!�؛~���A���#���u�o~��.�6w����B!d�#L�/�e����г�S�O*�i��Z�j��z�z|�=�Lir�Ɗ����_h���
e��"����O�v�m�믿�֭!��s��,B�����_,u~���ݶS]1����ncs�\7��jð̌�RJ����21��u}XF�?�KJ�b+�$��o<!a��_�T`��U��R�R
VZ�J�R���&bbmr�:.Z�������X�G�)�"���;��{�-B����G���L⹋o����f$�Km��=m���{��}�'��ً��,('�T�������߼�;���Ĺ���0_o�N��]\7̟?_��\"�졌����9��#1�%/��*��]��*��v=�J���sn�mď��@!dt�j�q����1�p�Ȓ>&1א2Α����~w=�!��B!$�^YU�Y������ӌ�?k���ݟ�8wh,و0���
�Fݟ������q�d���x���?�	�/���Bh�@�;��n�Ν����5��G�!$�T�����g��$�D�މ������V�s�=q�e�a����b_2����XúF�p�>��u�y�Ex}U>��mIjA�;!a�b��ٵh�2�DO�� ^��E*�`�qh��.&�h���>A�c��eeeR���/���o����P�ݎ7�:nn.#b�lǘ��.>�����@B�/~/�sO��]����l6u$(A����|NN��X�H�ss�5�/-,�������A��&+�]�6{�8�쳥ߕh	R�k�}�6��/ȷ����ݥ����Q�-u*��2XҀ/���N!��k؍[������?������C������M�ZB!���㝍c1}���<��ݟ�5C�Ρ\I�ޤ)��v��Z;4���a�7��k� Zckjj�`�<��cx��'uCIm�M��5���D�_6��g���;M��"e��e�y"�ŹU�N��]��\��¯����x�s�?�x�v�i�Aj�0��2֎�A+���06�{������j��QZ��0,E�g�w;;;�m�^G����$
�	���68�[݈��6�E����)S�*M9��1}�J�� �b���"�w���<�#�����o�w�}B!����*���X�Ad�n�6����4������t�,�]�;t*������[)PBH*��+1��p���9�!'+>�m��>���x��/0�JL B!��d��o_eUbJ�*_��\/��Ú�����Q��J����^3�+�`�͛�����rV�^�;V��!���Y*Q�O�sO��Δ�?{�7)봉 �=�k~"��E8S��'��NxG������,��uuu��������P�&�>he����$�]�خ���h��\N]��Q�P^���1i�z`<6�&.X��DB�;!���!��P���eҶO�J�Or74���	������`&w�خ]��`lA4��k����;����~�BIM�u�hK|����v�
Tf�b9.�v3c�O�2I`0La�Kn&��%�t�oI\�B!�g���mϼ��}��LE��q1=ߏ����-A�@b
}�B!���.
*jQ���ݟ5چ�n(��69��O^�����m^�W�0��+����ӦMCss3n��V���{���BI=���̙3q����"f��P�M�:��9�)������:>�t}�����!���X�ވe����.4��Y����1�Ѯ��dCS���4���U�@%t
WJ�� �g�B�D�H,�vAA�ϟ�]v�w�y'z{{A!���A$!�|��8��ӣ�V0�c�/�v+���6��jH#L��e�J�ܮIa([�Z�A!�:���?!�BI.D�������k����oB�'�!�w���c���5C9�R�x����.HthV4�=�h;a�)���g��]w�B!��&���8��3q�	'HI�^;��h�ۣ��Y��vq(C��u��M��J��IjC�;!Q��7�4O@_�i[����1��ݕU`���خ$��_q�L�;
Vf��h_$c��%�<�l����z|�� �B��gҤI��K�/�E"@i�)^y���=����͠˰��X��vEC~Q1^Y���!�B!���瓕C��� w�2i;�[/T�e�A�P���ݻ���]`^3t{M�z�����ܵ��ء��X+�fdd`�ܹ�~��4����BI�5���^�w�1ej��#��ve�0h0VaX���55D�XJ��2��	����(��t�T��΍>�J�ʠ$�h�_3V���W�h=�ݎ�`ξPK(�h�Z=Vޮ�����#����.L!�2����g�ƹ瞋�c��M�
��d�onW�/�	T	^�J�ܞ���7׏ŀS�EVBH��ï��WaM�V؁�vn�!{oB!�B���_mØ=i"��}z�Y��s�A�PQ*���]M���ĺ���F�S�L��wߍ�n����*!�2���G}4�9��Z3{,����nX;t���ܕ���H/��E-�"����(�r��m98��=]��}�P%��=����j;`��q��Qb���+тU4�	�Ġ�����Yg��=��7�|3�.]
B!��*++q���c�̙���h��#�ˮ��	T���0-s���hjWTF��R�ҊTY#ׅl.CW?E*B"e��K"��U��O���>���6!�̙>�=����\� �B!��^Z
�\�~����^(�{���}�xMVZ���[�&w��X3�fPVqq1�����X�`:;;A!���GEE�T;<蠃bZ;Lֺb�s�5C��a4����v���ٚ�ݡ��.��-�����wB���0�r{�q��{�_����	+��W,Q�\�B�`�� �b���B�'�y�n��nx������駟��!���L�>]�&N�U�v;Y*�}�2�k����M�VZ��4"UzF�����NB"gI������㯧�(��>']�7|��
$����=m&�8P�zp�}��B!�2zx�5s�ƣ�s��ܮ0����X(T`T3L�������]��5C�c�r�a�a��ɸ�����G��B!$y�6m�ϟ������
C96�u�X�ۥE���v����uC��^���\PZ��Z��OH2C�;!1`�	�km1fV���G�/�+T)�X����*�ocf�G�S������c�:��c�mk�*,,���G��^��[�r�JB!$���˓:�s�1��Ȱ� ���3��}�JqJ�O+LE��ndl�jlצ/�jd���q�`Ֆ!B���O�+���K
r�ܵ'��;^�+�Ǖ>&:�`�v��c�������7�kA!�B=S�Km����R�vuxJ&5Cy[�n�ً4hǇ���j���c�ӊ���|�7����a��X�������^����B!�$/999�7o�Ν;*j�v�#�����I�0Ts������
Z7T���v��_R�۲��9��wBb��A7��4�Ǻ�P�LK�dT7�"�,�!-��[�*^�����V�w�����m���.���kLf �B���w�]t���#�Bݎձv��ܮL_���]ܺBk)��t��SjK�C�&��	��L�Y��x`��{0���U��8�������`8��vB!�BF7���++�pX�}[��w�ݍ�v�Pt��j���]6��ռf(�21����a,��233� ��~�M7��o�!�B���v�MJm�v�mm[;L��b��v���$��d�}��ڡCSK,(��F>/8��#D�Đ��a|�^���y�,�7Y��w;�E�V���pe�� ��#������X+ǆ;��]VV�k����n��6ttt�B!�E��;�8)}A�0�E���X;�S����|��~k�H���FwS�J�4�b�M����j��	�%�L�"Q����BmE	������q����/���w�3Cs;!�B!��������م����0�#-GM����]��#�� �k���j���~{<��x���裏J�!�B쏨��8��3�^;�C�0�������bn׆c�kn���i�s���ݡ4�k�?���5Et��Ę����6�;�Y!�aIh��>㻩@�<"z�L�i�Ie0�L�
g_�Ɔ3W�m�|���i��p��7��?!�B��;�/�S�L���=�m;Tf�B�<�06�{����V��C���v�oh�`f�֦��,N��4��,H�����/�K
��{^��]�X�矾�8L�)3Cs;!�B!�E������\����4�wS]%`��j���&w1Ә &w�z��#��ŲF���8�!�G�4���B!ľ�/����ԩS��Vʱv٧W/�ܮ�!Z7�;+���`,Q;����[�Ǣ�As;!F��NHh�4���ZԻ���a/V�H�0��&�����oe"�L�`�}���2�A�]SS�;�o����N��B!6!++KJm?�3���7*�P�&B��M_���e�{l��C�"�6�AޖƔ4��e4�O��]����c���SP_5KWm��g�*����ڇ9W>�!�B!$u��v�+��T�Hj�!!j�����Տh�1ɺ��13�ۥfm�z�k����v��<���<��s��E!�� R��Ν����7(((`�0����~��e���ˊ��}H�خ���&�k�۳���QW9�\ �C�;!q�N�V7����s��:-- W!�bUzz��T$�`ev>�}��g�H�3220k�,L�<Y2���� �BH��y������첋�Z��H沫xejn"R�-A*�K�خ4�MmW
U^�*��o�R�"$��Ի#�n̟;�p��;�IK���ڇ�hn'IBq~n��,�+ʕ���߉z�B!��TCt�:c�f���Y�ñ�V�UIT־$s�%����)w~�l��n�brW>�x��Ý�h����\r	���~��X�t)!��x����?�{ｷ�m�z$s٩vhnn��:?���±�en7Km׮�I�%�㱮�	B�94�G�\=��k1�w�Ȗ��n0�g��j�{@���T��+�9ceV���e��Xm�����nÿ��/)�}Æ �BH������ܨ
J�n���x�W���ւZ����n&R��۝f� �J���P�7�d���	I$���=����/��}�O��v~�#��(/��Lm� mO�҈Ң<\p�+ �����z��uk���z9���bD�f'�+jј�L�$�:���:nD���]�UuC�P����a���ѬZ�?Z��k���4�|���$}�B!�G���t�I8����l;Y��f���v��a@�P'+Z�v���]el�C�4�Cq�?f�i��Ųͼ�#�
4�g>]������1�K�V��so�T�(	V�ڧ|N�������x�t�A�2e
,X ����@!���"�E���?;찃nA�.T4粋@e����nfl7��(�7�;u�z�vS��'T9�UV��[x�F���ɝ�v�l��f���2�����~sHj1fL�&��uM�3]x��)eI˚�=�¼l��Ǣbl!Č�7!}|��$-A �$a�
���$מ|5Ñ���
�Rv~V��S�5�h�#�&:�;}�t)���~ !�B�ǎ;�(�EQ`W�z$�ڥ���on�3��r����C&�v�C����%.�[�&�in'�*4�� >]���'6���u�M�k���n�{��d���9�y"�7s+���WUU�n�A���N��B!1"??��vN8�)�!��T���(P	��:�-�۵b��0���
�ܮ�^p�6��/.���;!L�'.?逸���v����$���љ�B+��U�c�%�b��@l�0�?}�q82A��Yx��ˤjB���vc�P�l����C���m�������Ё5C��D'�T�Z1�Gc[��z�!<���200 B!������c��g�a�����XϺ�|�cjn�t{V�����B���v��}(Hr����jk���1��n�梟b
�$�ڝ���&�nmS�K�ұ��D��L5����cx�5�<VE�p�鍵��$��b9���%����ƫ���:�B!���~����Css���h�b5֚@%�7���h�ܮ5���*M��+4s�R�����6��/.B��X��G�m<M�4��ddBY�*K@R����j{�����_/?G\�8z Į�+��?�?�^��X���q;oq~���8�m!$�Y7�1�0ah���bR+�خ�y����T�B�Ь�>�=�v^^~���Jz�m�݆o���B�.�=W��ϟ?;�3k�qاgnW�hn7����B�"2��u|����]X�� }��4��@�mwbFCе,`_D�n(4����z��4��x�O�%3�zY�J3^b�Oz�a��zl4�e��|����kp�Aa��駟@!���)--řg��#�<R��_"ŨH�cul<�P[��Q����>��us�J����ʪ�<��ؚx��in'��4g�$KZ�������~1�p̔��x��_c�Oah争�RR��g�>'��>��򘟯j\���ɍU ��p�z���(�o�/���ڵHV���]><X��^��\3�[Z{��v�	��?�q)ͽ���B����"��HnO�����d1��5��p,X�ۍ��ۅ�]�v�1�7b1�턄�$����p`c#�ٛ�n"R���Y����S,	VдT$3�Ee"C�+�cO�(��`���>�:u*�y�<������!�B�#�ifϞ-��+++��(�Ĭ���MZ�[[�d��А3ts�7�!�l<�o����d@��ǌIì�m�s���y?����$�nC�{��'��!{o���L�1��܀��������HH���i|Q^6�~���.�Z�X1u���c0����1'!D�竇�gu���I�[g͌�t�Nc��f�u���F(F&��5�P�srr$}sƌR����B	��*�S��ߡ�����C;�
C��ݳ�nh���Z0�lj���1��܊y7�7`���6  ��IDATJ��		�	�o�9q`c�yY��Mn���/���(���p�*X)�aUL��(e��v��Ǔ���SO=ӦMÝwމ�>��B	ΤI�$q��?���E&�����*n%N�
?}A��hrWR.���%s{i^l�
�RB�}X�܇�B	dJ�x��dmG7���ǘ?w��9�'�}�f��Ի $^���p�uO�ֳ���BK�df�K�g�#.y�u�������������X���޴�?�6!Dar߻�c�D��a:֊�*��Rw�����5C��i��%�fI�/�5�h_�)677�;��;�#�W�ZB!�X���g�q;�0_�h�
��v��rl4���E�kP7ԫj��c��C2��[o�pHeno�'4�4�b�js�WM�pt�nr���{Py�B�
K��)yd�B� �*.ES�J���HD-����&,X� �����ΰa�	!�=���p�	'��OFnnn�bS���`|�T�
7}!���#VI��+�@e��n`n/(����p��N!d ޶wj�I]D��c����b�q8f6m��#�}B��[_-����õ���3�X>��;7ཻ���}��]���A�:18�OR��;����d!#ã�]�(?Y#ۓ�����8?'�ǿ�eN�����!���j'~>�[[U�[�*�����_��������҇W3��q=Z5?���Hk�b������>������E!�c���q�QGa޼y())a�0
cC�*���Fv��ݻn�������B����wy]��Z؈OV��NH���N��X�:�Y�pl
4��IKzFt�[!PI�[�8k:�P^$�Ņ*�]$�h�B'n_"�|�|����Mʊ	>��V���>��C��^{�{��k��&]�B!�����q�9�H_���9�%@E2W,�+S�
��J�����skfpw5��cn��J�КIs;!��QC]�X�e��.'n��wp���t�u�,����� $^l����z	o/n�mgj�5+#}�����$�����<��	!���݉iuM��V�ܭ���[���ļV��SZ���x��Q���=ܹ�n;�r�h�q��a��������o�?��[_&�BR��N;I��=���w�vL$�ўst����c9M�������_҈���?!рwBl�k-Ø%%�/�8c1B+Z��+!TɷR�;4��(�<I�O���k�m��/�W^^����Gq.\�����BH*SSS��O?=얂V��i;Vǆ;�����v=�ʸ�ఁ�]ahw�'0	UJA*0��/���vB!A�p�tdg�_��-/I���/w�4r}��h�r�sk�噎K9���~#�ɀc���$ux����ﶵx����c}%����e����k1!$�_�Č�F���w�5!M}0�y٭^q�ӽM���\�>Ǻf+#{4k�����5��SC�u�]�$���z
�<�z{{A!������v�Ν����QW+�n'�̮��3����R�͍����4aX.}s��~�W3T������D�WTIA^ku��m^�C+R�tS|���`�� '2x��y�!b[\�$��K*��VE-�c�L��{��-�c�=FъBHʑ�����>Z2��*bT4戗y=���!Pi�ĭQ[���a�J_�
����t�핒��9B!IDiQ�8�@��d�t�Ʈ^\��[���왇�"&��(s�o~���KBCnv&��㑰W<�O<��g �CۚNr�#���Cp܁Sa7��l���<ZVw�B����.L�oDږ6�1�X�z�[9�ʷ�-����� i��U3�EM�i�B#=�Sp��/�^}�UB!�Jzz::� �u�Y���N��a����)f�C�����v�`��n�N�+h(����Q҄win'$���N�M�g�0f6�����4�P+�?=���`��Ifٖ�ޡJb��>+���1�����f��/�9�h5{�l�ﾒ���g��.�!����~�퇳�>�m���mw�)���"PYI_0n-8���-]��А~{� s�V���/�Z��r��&�b'2������b�mk�:�r\θ�Y��؅)M�q܁�5�ۍ�N< �}�#Vo��:����~�g9n��,��d&�!I���9�}�͑�.BH$��܅i�M�71���z>m��������w�C2�ۨfI]/Qi�Ѫ)Z����W\q<�@<���X�d	!��TA�N�<Y��瞾��c̶�9�N۱:��<�ui`8��vhP7�3�w}4��&vC��Y(�^ ��V��-n�4�uhp'����m66 �����d-�|ӗo�+�j�J9��p�Lc𥹏,�ANfHK��1e"�Z�R>�h�R���!y��1eee�?>9�,X� _~�e�/HB!�Iss3�͛�3f��9db!FEc;
RᎵ$PE��hpv���AD*3s�Y{���	x�%��vBIB�L���]p�϶���4���- ����}�sI���de��?����z<��XҲ�=�E�z)�7����/���U�_���j�P�#L�:#�7n�,��B��ʺ�\3T��#15�h�c]#�G�����>�}����s��G��͛A!��fJKK�n&�s233cR���^;T��=�r�PYC��ܽ�C�]���X�Z�+�vh�e��Y��]؄�2JH,�����V���؈�nu*���^m��R�2�<�-����9���4�4i[�#0�A����(M�z�&�h��c!Z	v�a�w�}X�h��^�]��B�h 77W�N<�Di}4�Q�n��Xk���/��4��i/�W:/��������eG<GQ~�s-�ƂRϟKJ�t�&�����f��NGq~N��->�<��q�����~BH��d���n���e����!�A�
���V��W<�B�N�\�j��ܢf<��>5C���QS4#:@w�q�9s��������B!����̚5���oQYYV�ʘdގ�X�$�-_�PZ�=!����F&wW`�˿m�ܮ��,��Z؀�V��NH�����$��v�dr��n�nsI�ֻW7���V�U���P%3xE+��HwW]̈T �/���}E�dH^G�J�G����x�	<��3���!�������?��v����&N�s�]�H��*P	�#������ghw�TA*=�ʻ�SV����BI���q᱿��غ�o~��؅��M�A�|��J���5��C�|�����9t/�t�n(/ɏ��C.������ŏ��KB�%��vb���/��
xA2�u��B�;@�	�3������4w��X#���h�>�7F� }��K�/^̀B!��)S�ଳ��ԩS��x���1G��
���@� s�b1Jm�^7�1����������m�U�#����NHL����$A�ܧ�5!ߛ� V)D#��s�VhVn�v�/R��*�1I!RAn;�Hpcx�G���i��M,E�pE�P�H��>�p��S\\�s�=�gϖ�^y��"�BIv�m7)uA�
���l�]ŭh
TJ��5��/L	�H)X�)�P�Jb��`(R9�SZ�in'���g��.�Ӹ���AIAnHǮٴg��<z �.\��h�.��Ղxx�#�ɘ�HQ���w��BF��rb��zT,Ð�O�kfD�o|uBU����@s�R��#5�H�|��&´NQo�N;�x ���*z�!�^��BH2��Ѐ3�8t���h����u��.�B��*�jr�P�~hT7ԫw}���v|V��j�rJ��~(n�n�f5`�j��	�54��D��}j�P���i=(��b�Y��R�
8�/V�}ij}������E+9�Ay>Y�2�����F[�B(�U]]���Jv�ax�G�t�h����X�8NN�Z+�D۫D!R�E��D�ȟ��s��>�?�g���.H��^�[<�D��'���D���}����.ĩN8�P�����1v5��{l$U4��"���]���/([��ܲ:��Bs;!ɀxI:��=���
t��し?�Ʈ^ؙ}v��#��$��>�޿��w� �E$;��ۅ d4�����=��+A0r8����#A�!�W�\��.�1��L�/$��@k���U�T$����C�Z[3��ӭ�i�~�0���h��beZ�U�v[�9c�<��x��'���B!$(,,����O<���q3��sL*��A±t��w���p,�Sܧ���'Z���4���n�0�f5b�Z��	�4��d|�r��6����w�_o��֭	Vj�J��{.$�b�����a0mME�4��D�`�|���B���m��3��1����.���R:�ʕ+�bJ���M�D ��x��盨�gee%�܂D�����D�_�����^��s��߼x�~��|s<1��x<���RI��3g���X�SV�$Z�J�\���*�G�֤��/(�*�"���@edr�(��[@In�7'��o���w�}Y��̎%9���_a��ɐ_R�0�����r)H�Ѻ��7n�[��ɍU ����u�7�kA!�����C�j@�s����EY7���U��݊���f���*g�X3�GGҫ��i�Q3�R�-AXVj�� xꩧ����L�-���+jW�$�痃�䰚x��?{�3?�D���'����Z<w��E<���{A�~����u;���ӭ�wF�T��?�C9'�t���,����G�/s$c�P��Hh�����6�{n����Pp�{��ݻ.X�Ո��NHܠ���$D��w߄	C�U�ҍbݳjlt�]D�/VYi=��If�"8Q� ;D+�,\)��^��+J�A�Jt��1Vƈ��������^���7oF$����d"H��X�|ip�/�evM��^~�I�}"����a*~�@	����>��g/��"=H�,//��8eeL�ŧXoG��`���=4�J-N	ûn��N{AS��������ڒ��:;7�W���yٸ��_a��-�������p�/&���L����)�u��}�#����2|x�� �B!��uC��G��ro��[U+T�b���
��|G�w����Y�P�'��=�v1:>5C�eY}<��a���Ə��.��f����ߏ�?�8j�����v]K��e����)�$U�"�Yև��g�= �ά�w�&K#�F9L� !� Eƀ ��c��:,go���y��ߵ�������%$`�D"#,��Q�a$MN=�߼��vWUߪ�U]�]=s��ݷ�	i��3���|����y�ݞ�����y�3���gϐ���>������_,������Ax|:sƲw�tΘG�b1�#4y�#��nޡ�34�cY���;>�y�v�v~ΟG[im@�����; 
ou20u.5%v$+y�A�"�X�Tҝ�m��9)R�����u�,�m��73�w)Zeb�xNX���)̦� (AJg	�-[F�\r	��������^   cٺp�m�QSS�˕8�3'j�V.�e��!P�50��w��v�H�s�&4ӳ���C"  ���K\��'��|Lrc�u�vSTش��:{���     ��~� ��ϡ��v	�C`	�'�&Gf��ͻ?'���=y����A����y]x�a�`����Us.\(v�~���?��?hÆ   ��w�!��}��������w�;�xoi����^}C�b��w�����v>JJK��,z� �� ��9|  m����I�����ɭP� ������1yS!�'+�Pb�z0-TY�i�j�AtO#�*"�؊0w�����k����ٮq�4i}��n����>tO��   @��}�٢u�N��D~�E]�
��_�*mp�T�w}�*njl�cj�h_07/�ĩ�p�lo7T|���fzak�v�   0����I�vPT��o����_�B     �0hm��������V脡��%���td'���I��ŗg���I{�|}����u6��WO0�׺��5����Yg�E��v=�������v��E   @.ijj��~����}H�d��5��^�]��:����ڵ�����w|v�+v|��>�+��׻���vx� ��(p6�Q���tZ�>�7ni$+rnb0�d$�96��P%5�D�}�A	�ԸݭM�i�J^'W"T.�������|={�l��W�B�^{���x�	q�   	�9�S�8�x��y����Zwl,�߃Z�j]V�r��4�+�TT�D�T5��!P  �-��������"�    Phl;����t�����c��(n'�&��ٲ'��a%y� <C�.�#���ǌZaP�aО`<�0甕����_OW\q=���b�{�   &t��7Ӳe˨��"0_0�9Q�ú��;�� ��o���<CS1������v|������}
��w@�@��Q���!�M���ۨ��;%X%��av��!Zɛ�&��@��"��L
W��Ny���=����+�����R���wz����sM�st�͟?�����n��F��/~A�>��B�   �s���-��B�^z��g��8�gM�_;�˵@e�䶂CC���N������-%ʹ~v�  �{^۰���Koo#     Px���g�&�ES�Po��.A6���)�n��M����̕����9:�Q�UUU	�pɒ%��ϰ���   � ?~<�p����|�&L��w��n�{�����af!�|��o��cs{�;4z��r�ʚZzz�D:܋�O �	� �t���d����1V)�Jf7�&�*�,����0r��̐le0�K�DU�7!B�*2l=(E+qXW��������.�慠)]��N��~���v�Z��L���
   ~�3g��_s�5TZZ�wqJgN�Z�s��vkc;#�(�@��w�*0�jD�ri_�in磤��6΢�n  ������{;�o F�     �{��؞	t���j?dnq���v^��1lϐ�BR�M�!?����F�#�u�=�:�aÏ}�ct�W����/���   ������.]*v|�2e�oP5�+��Ϛ(z������z����_�{�v��q�o8��n	���]��k�O�G��Rw�  � ��#�CB��|V1u9l�SJ�J>U50XĪ���!-z��B���Zd3C�փ2�n�I�*�<�>�G)X?�lD"���l_�~|~��w��{ٍ�|�������{�9��OJ6l���   @&�u�������@5nܸ��t��:��c���N���!���d�}H��])R�)���Jz�s*���ւ   ���Z�yE���!��7ѥ�M     ���HЃ;�i���>|`���4�[��v�aJ)@��f^�������x�f��J����/H�/�{��v���ɓ鮻�%&����C��	   ��7����3g�1?���XT��^��*�
���C��v�b,�ops{��zzh[5�ǐy 
 ��(CV�j��R�j۟��V�
2���Sc�g��'�V����I�����dн(��`k�OZ�J�v���֚0��q����O/��"��g?�u��!�   ��1{�l�馛��k�����@�(�X!X������}����a7���ڕ������z�P=�F�  @nx�͍t�9Ǚƾ}�s�o��u��t��TY^�{o�j�@# ��8oQ3͙RGQb�C�f�V �0���RA�4O�����&w2��Dꂬ�3�w�Щ�]��m(V5�g�ce���Rϗ��u����0�����вe�D��w�����    '�/������[o���F1���w�Cw��z�hl���5�����lo��<�V���PT[ � �0
J��M�tM��n�m
��T%�Pe|�jeQ�L�r��$�M����:螺�H��i�A���U���pu�Ma�v�x���y���:��9�C�/���~�󟋠;   �_#�ΝK7�|�خ��l�Y��5�
Pn������@e#N�TZ��#�P,��j^�k_0	S���	u������?D   @���V�c��c���������HQ孍������+7PmU9m�w�n�?��vw0�9�q*M�PM;��-{Qԩ_E���{�W6l�� H>����'ŷcye�s�p �X|�sΦ2�z�,�;�CY�e���X�q7�0l'��ar�������E�]��q�b7�c9{�E�|�a>��r�!z��ͺ��&���{EPq���j�*4�  Ȁ��%K��-��B---b,߾`PsF�wh�����s�oh��5�C'��T��볭wh�۳�p{�,Z�ZL�� D���]�ZJ�7�۶'GD*�p�jb�he0�V	�h%稄��he�g44(�����71�д�w(���Vˏ]�ȁ�����f������;�<Z�f�򗿤�k�  ��	�o��F�=m.��\�S~�D��^P<3���sq�8�"LǍ�v{��lO70��TN��,P�Ll���WR�  �c�b�ﮠ{Z+��쥨���ʹ����մ�`;�	�n��t���.����{�8���7���u��S�`-��>@_��TWS!ƞ|�}��?�W�Г��b���3	  �:�Y������H�m��~��K�Р�94�{����ӵ�G�;4x�F���Xv���K�Я��տ+������P�j�������u�]G��կ��#   ��B.��b���F1��`�ε�~��wh�[�錾��;��u�۝��<ϩ��*Z��|��&Z�Z Qw F9��]��Ltds�&�(S�R�V��ɌS�h�67����i�J�I����U
s#CR�J�ܓcىPQ��%Z鼷�:�1>�>�l�����/ӏ�c��nC  �ZX��馛�ꫯ[�#خ�J�=�kxy�tNjw�┎@e�[��*_[*Ī��3iek)�  �7�KО�N*$�z�F?��L_���Th������T���������ڻ�(J�������7�]���诮]L���c�;���6   �Yݚ�����l�}CRܭ�!ix�:�?z�1�^�lpWy�EER�J�9cY_g�	F�S�:ǯ���8o�<�������鷿�-�X���  0����GߛP�=@��F�Wh}���˱����ή�z�X����/�-�R��|�&z�;VUp`����9���{���@f+CJp"��A�2��^Z����ײ����V�sqV�J�L���32��GΊ�وJ~B���^�/�k�9'�1>�:�,:��3E����^z�   �>�s��hٲeB�*---�`{Ps��:}&^�
��"N��)՘]��N�J��kn-�jl7�/�7��/ �    �b��zR��Ҭ�	4i|U���6NQ�7M�D`lû �  j��2Dg�n�����34�ۍ�!Q�6d|n
�+<Ñ+����*�X���<��3$ˎ�F���'�+O��5��	r��؜9s�_�"]������GA�  � ����[n_�(��~׍f��)Ԟ<���y����\|Cǀ�����%�����fzc�  �� �^���6SmA��Dj���<%@����S[�O+�w��aE\sD��&�p��z�~��ԫ"u3C�!� '?"QP�R�B�1t��O�=����裏&o   4�9���N�k����;�<�<*�v�X���A\#8��x�'���s7qJG�rk^H���*׭!w�n��fz�5F      ���go8�>q�  ��Wv��MtL�.�����к�gH��a"Q�k�g#�/,J��l��EZ��]���#�u�=h0bcc#}��_��n��~��ϰ���   �.jkki�ҥ�kƌbl4��:s��Z_;y��\��7�;?���*��Z�e���ȣ]���7䣤����E��BN	����; c���ґ�YtZ�~���5܍7qJ�:�$yc�z0}SSb�ҍd�~FJ�ۇojR�U����|�%�+y�ea��γ}m}��~�����ur=v�	'����Z�z5-_��zzz  @a������t�u��駟�2�������?A^+_��\�v
�[��T�J����ۍ"U`�B�b�U4��m�     0�Yz�B��_@   �y�@���f�i5���������#�x�5�=C�|�ݟ3�C�Gv}&C؝�B�%ړ�s��)f�����
cl֬Y�/|�>�я��;��$   �͔)S��o�����&MJ��`��u��;T�3�C�o�j�R���-�X�;>;�+*+�厩���! � � �1v����xZ;uwq��Ū��e��ܭaw�ΐ�TXE�l�g���� ��a��r�|�555�=��C7�|3=��Ct�����Ç	  @�)//�+������Z:��c�X6����B�G]�J�s�W����~�(NY����S����]C��mmW�Uee��nl6���      �v�m�J�v�U�qf��.���?���~�'���  @�Iz�S��iG���=p�34�cI_(��=��S�}���g����g��!:
�aT=�l�e;���@w�y��~�a��ر�   ���"�~�UWQUUUV�`�cA�mޡS�=y^�7t�݊���3��*�P{�gEȽ�v<=�"�E��Bw � G���Ȯ	t��R�:r�F�J���xe�S*�N)��T٭��f�V�I���i�A��nYEFK���������#X�R�]5�?�����b�
q�۷�   D�	&Q�n�:L.��|��s!Fe{k�]>f
T��q�0e��D)�9c�]%R%�)s��1�n'P�D*Ŗ�����*z�H��D�     ��NmU9���7PUE���/���y��   $a���i��q�uhr��7$����3���3�2����C�Zʱ�~�zh�&v�a.C����jkkEȝw}��'���w�y�   D��`�����˨��,R�v�X>��w(����*�����C��5}Cۀ�C1��� �Ll���WR_,N ��w �(��qz`K-m�I�m;m�t���|������	?;��,\��˸��5�.���f�$R�yUD��E�ǠE�\�XaΉ�X]]�q�t뭷�3�<C<� ���   �̜9S�Y��;��`�j,jV>-��faJ-R)�)�ւ:"�N�BR�ro_�����G��:zb�x��G#"      c���+�y�$�y�~�����   31�������Ӷ��3t
�KR���g�����Aw;�aw�_h��#��W?/�к��z�`��A�_��rQJ��������^˘   ���ŋ�ݞ�;�<*r�Z\H�v��F�wh*Ĳx�N��V����w}6��ߐ�Y�BU���;�p{U�lZ�ZBC�� ��@��1�P�H|�PK#ڪ����2%L�+kK�5�lq7^S��.�S����T�LR�"�6���D+�"��5�uL%2�r���%K�Х�^*�U�V��;ߠ  ���~:-]��.��@��-Dq�Ϛ0-'a*y^j��UN�v>�l�[
�k_��ZP!R�L�NnG�C�      ܶ��t��6�<H�ߏ   5�>�ZJW�k��6�gHd���8���-��7���z�V���g�hqWy���#�a���l�??����(�ڭa;�8����$�ׯ��+W�O<A}}}   ?TUU��_N�\s�hng����sN>����5���;T��nޡN1V,������n�n�a,6H����r��� � �M	:sv��n?��'��S�!�Zc��(X���N��aڂP�ߥY��7m����KA�Ma�ڝB�ټ��5��p%[�n��~�V�^M�ʘ   ���8����)��"����]��`�Μ\�Q��n�c�t�)�XR����3�4��{j_P�T|��~-oM�^      ����4��n��u^�@�>����7@   �y�5A��i���-40���<Ì��P<��X$�d!�9�.w�6����BU���3�B*�>Z<� �������ԧ>%B���oh���   7L�:U�q�u������X!�Uc��+��V{�f1n�u���q��^��?���]�q��;��ή�za
4(dp ^��c�4����;ykcp
��JK���%
��Ķ��vO�SE�-M��H�F^#H�)**�T��xcc#}�3���o�]��W�X!B�� @0444�UW]%�S��2w������U�Xe+LY���T"�5؞l_��T��*q�Q�2�T�D��k���VT   
�����Ʃ"l��{;	  �7�JK�??-U�s�����Oһ��   =����6S3�Hz��pWd|�η��l���ܭޡq��/d�*���'�n���D"rO�n{�WO.J�v?~�)S��[o�o���z�)���M���B  ���?\č��!VTT��Us�ձ���wh���<{�n��V1��o�۳�oh�K�JiSb6��}�  �� ��ҡ�t��6����Z�"�p���Y�R53$��m?(�*�-�t�!L�VA	LaP��r%<e�����n��f�馛��_��{LX,�  �n=��E�a
S^�FQ�ҙ�����I�J��)��v���8e����8e��l�)�p��H�Uk|.�y;��   
�������A�3&�����3��/   }n[r
-l��:��76�O�:  ���}�tx�L:}����I{~�9N�k�Y��靟e���oh�Sa��P�ݓX�B3~<à<E?��Y��:Q�2��lִ9t��믋b��~!  ��q���/�=�z�b�P}B�1x�f�P����!�Zۭ���?h����U�5��p=��D��� �  {;���މtUcu����lE+"�5f��i�A;�*%TY[��J���>��I�6ZR�
S�
S����uY�\�x�8>��O��O?M+W��;v   g&L�@K�,�q�'Ƽ�Mv�Q��$`}�0e0���m��*�����!�ւv�v-����^j�B�;n  P8����ޒ
�3��i˞C�z�  �GC]��=m�t��"��  @���Ct�w2]>������Nޡ�7�ls�b��w(���Gq<.�T9��7Lb���~<�|�ؽ�w���-�q>N;�4q�ٳ��x�	Z�j�B  ���3�Ȼ=�s�v�uQ����LQu�����C�b,�p{zh�2,7�06|���L�L��UM��C  � Ƞ?�����ʖ94pp��V���`e�KLAw���20f�*-V%��Fa+��z�D+�s�\�6�w���Κ5���/��n��z饗D�}͚5�&  @�c�9Fl!�����Z1�Ka���(�S:s������Eu�=S�r�V�)Ԯ�gn-��������^[WO���~��  j*�9S2Ư9�8�  @��	�����C=  �?]qz`s]�2�znOjM���k1i�0����[܍c�~!#�B5~<�0<E�9^��(����O�N��v�������W^y~!  8PZZJg�u���.���21�����Q��|y�V��8�W�e��y;�0�p{U�,Z�ZJC	��; @၀; @I"QD�[�>��B�G�؋O��͏b,� �s�`e�~�M�������)�ȩ�A"����:S!���&�bQ>�'��ݮ��l�{��ضm=�����Sww7 �X�ۮyA��~��b,�n<�"V��)?k�U�0e��[
f�U6��q��������F06"R��)�Hen�BԠ]�}D�z@Tq   
���U����$   ��������J   �g(QD�Z�.in�����mX]q������r#���\�%���B��;���.?^��:�zN��t�]cܸqt�E�c����/|�G���   �ĉE)MMMbl,���c�
�g{m��a�g�P�w��s�o��}�ۥ��RbR��'�^ &� yjs�N��Ds����xK���<4�,u��x�$�`E���lg�؉V2�.Ī�J-T�E���E�ms�2'�u~�������s�ҧ?�i���?N�>�,=��S��/���  0��υ��~饗
a���.5n7_w|4�X�d����B�,C���P�U����Z۝�\[��T�*R���,tQ=*   ���	������4i|��   w��XC   �����贙-4�k�3��z9�^a���K��n��_h���8l��{~.�5+|.�к1�9Qs���������|���Nz�'D1�믿.tO  k��R.���~�������?/׈�X���(x��1c1V����ש��v�B,�%���Ụ��	 0:A� �ʺ=1:2q}�z���P*��pã����JK3�d����`'Z��܇�;v/2������z�7�:�S�!���B��������E���;v���{z��h˖-�  �Δ)S�K.��8��!4y����KQ+�k8	S��N[
�(�P�s��lav�m���#���)o�77�   (d�j*m�-�;�֬�J   �cp�{�8�>  ��vRӤ���r/����>����>�C���'hW�%}C�?(��I0��d%���3$�5��������;������A�׽\�����.]*���Vv���~G{��!  ����3fВ%K��.?�#���g;�+�P5^a���F�ޡͮ�:�X:�X;>��~�r�gKН�9��o:m:�p; �� Zl;����lvuڟb��˛���2׹���d�����*PYǄXemf��������@U�U�!�0�|�ڽ�QAW:�gϦ;n��vZ�~������A  P���Wn[��+�.�ն�xԃ�(	XN�HR���{5'aJ�C�vBU��v��{EU��5�v�G�  @�3������Ʃ�    �ȳ�P�ګ���tPg����d������N~�[����Tv7�c�1�1r؝�,Y
Y���vS�m�ٮ�2Gw�Ϻl�7��:�����'>�	Z�f��
��y���#  -p���Σ�.���>�l�'2��f�>�~b.�����C9�����<�ۭ;@�c����S{k�p/�C F;� ���ӊ��te�l��,8��W� ��Y�<�I
T雰�p%�(5�N�b�0ejrigP7��U��]���u6k���y�\�97�q~<��q�]wѓO>)ī��zK�4 @���c,��/�X�-ps����t-��|�X����z�S�=}^ue��n��`��ĩt�=f��ۥX�p���J�l����!   FU�e��o�N      �z����j����znW������]����m��r,�]�=�/�mr7{�d)ʒב�e/4���{{}P����'G����z�~�a���,�� @�a��k��ɩq���/��;�C�B,Sk��7t�[��:����3i��R��k4 c� ����V��9���{������F�op4*���&*砻Q�RWv�r,�����vc3C�HeE%Z!b=G���՘����������Z�v������O�S�  �7����/��-Z$Ƃ
�5�`�j,J��k�Y��R"���$Ly����H��Ӑf�=%N)ĪXl�J��ҊM�qC�  0z()��1�㛧      ��P��V�]��L��[\u);���?4z��6�d�=��j�z�ZM�#�w+<5m�ks�cQ��|�^�r�>��'���_/�6�b,�<� i��شi�D�����Ɲք5�O���B��\#�:x��J���]�����w�
����l��=ao]3=ފR, �� |��5M�K'U�����͏!��'�nlp7
W���t�]�Π��Aw��3�U�v��@%���Gy��U�ʇ ��P��`�G���~��1��9s&�|�ʹl�2z�����_֖-[ ^ �F}}=�s�9"�~�g��B�Ϛl�%/׈�X��)�9VAʩyAi~��M�����TZ��ǘ!��=�n���5|�}Z[�<z�u����   �H���na�gM�ڪr���'      
�g�т�f:�tw�+C�r	�Km*���BØ�U����|B����0�r#hJ�S{����a���<���˧7�e��k�^�x��c��=��Co��&=��s���SGG�B @d��a�=ĳ�>[|-e��5��`|Pa����Q���X�R,��c���J?�l\��g��[	 0�@� ��-�c��g2]1��:H��(��q����Z%%z!w;�J�7~F�ʮ�A#O5�J��9�\�k���ݵ��裏���.��~�iq:t�t�{��Ӹ=f.�luuu�Ķq��Q��?s��(���F���|�ٳx¿�|mߙ��;������������O�o�*_a�׃/İ{P��䣝H�y���v��v�@5����@e��.���*Z�;�6�@  `t��7`{�����>��{�]     ��x�@��UM����Sw���F%�C�;?'�ڗ[�]b�	�x�~���&�>���\�e�Kyi�%��.���������;�T�=�����g��uz>��nz��W�g����z������ �.���"����̻�3Q��S�Z���;��z�r<��w(��Cc��T�e��<��3<C�)��'�s&ҁnx� �Ep dEw��\EW�̢����7G�J��~�C63��gW�b�*��t7�U���
T4r6�6w�5^��W>ǂ��͸�5���x���O�^~�ez���u��aG��^�����G��?����
l���@���5&_���������H}S�/��{�s,,����Z�?���Yg�E^xa�$����)*�|�q
���;4/$��n�v�p���=����IS�U�5���   @�t�8o��OO��H��j     �z�j[-]�\C�������n1V���*Ŋ��ܝB��]�����5׵��B�ϊ�ڝ�#$E��|�����P{�A� ���]�iMUU�(�������z͚5�7d�T�竜)�A�~�3�?�|�3���U����Οk�j1Vex|�N8A4�_|�Ţ��ɧ8�<�\��������X�;>�l<CyTO�In.��8�R �*� �fh�&���bZ<��&�lARS+C�x���7X�6w'���8���t�D���e���Tm�f�ʊ�+��8�m=ʂT>��l�u������#_�җh�ڵB�⦆ݻw  x���8��y%ۦ�s���0��X.,�%�e�T^[۝�)�p{����оP9y��T<|_�q   ��:�r��)�w������	     �B#'Z�ZD�47S���~�g��j<�*�A�r,�������^�v���3����:?c~�������:��p�>�!q�ݻ��{�9Q����;����)���D����a���;��r*��LA��ۛ��;��?{��>����$dS{CC���a�<�B��TF��?��;{�<G`��ҥX�ޡ�g����5���0�A� k����sia�^���$������p|���$b��4�����I��4��a'X���w�-�XP��(����
N�B��@�t�E(�-�]w�Eo���hk���@;w�$  ����^����nk��&hQ�������cVa�(X�ϻ4/$���*�慴Penmw�L��������k[���9� !  dä�U5��W�8��:�W�AX���Y�J      "��<D�4����"L��z��9nis����_�|m��|n*�2�m��G9�o�=L0j��h��O�N˖-������W_aw���3 �0�P��'�L�w��O�:U���#��&����B�{�}���&c�`��R���+<C�+����f�IooŎ�  � ����)�BKf�Pס�����A������,Z�O�f�3�-�w'�*����@2�>��n
���X�*3��t��1��~��;��~�ɟ�惷%\�n���ք� ����?O,^�8���P��5a�[A[Q��E(�,C�r:T[;;�S:�vlE�240TU��+�� * @�|��K����V>�v�?�=������8���dO[���8���v�*����t�gD���     �"���5���ɇ���H�+4iZ���ӥX��{�d�Wt����N^a��,��������_��l�u����9�^y��8|������A�= ]xw��;�Ǻ�:1�0��(�Uc�����=T���P�4�b���w����G��I������� �w @�t��i��
������l��,��U�=����.�IQ*y#�����Nb�Q�2�U�Fw�6�4a�V:׉�Xs��?.Z�H��smٲE�����khk `�_W�9���Ρ��N:)��'���ӹB��Y��u���A�.���J�R�S���N��T�v?���=C��<��:��b�  �����64\VZB?��5�PWC?Z�
勪�2��/^�nw����ᯩ��'�{w/u�7yB5��篥��%ű�	     (L�uѪ��tes���4k]
�0ᢁ��ܭ-�	�Prw
��С͝F��$��}�{�s�c�����xPk��'M�DW]u�8:;;EН��_y�:x�r- `l�;=s����N����Z1���������Y�K����\���s�c�����z��:�v�p��7Lۇ���Xv>��nϩs�AW?��D4��  Hp ���7�i�&:�t7��o�4�����%螾Y��G��C�NbU�1�>����^T�׋�h�� �5��sMMM���멽�]���x��h�޽� ETUU	1�SN���ٳS���ӝ��S�
K�ʅ�%q�\�t��	T���t�=)B9�Ucn߳Ml��C  A��@;]������V�X[�q������/��S�D�8���o��~�w���cf��yfm+}��W����::oQ]{�q���H_��<����#      
�X�hUk1-��L�z�S����_h�o)K�F��3wv
���B��Z���Q���6w�o�v�r�����_�ܰƃ^c=?~�x������Z�[o�Eo��(�z���0�������;<��Sš�ӳ����ڽ�G)خ˕�h�/�2<D]�0p��l�Z����Q<|_v���^iE)  � ���FM��#m�&v�f'�*�6W���������GnO���*�`e���n���hejN�Ƃ��x>��b^x�8>���Ѻu����_ֻ�+�� 
)H�y�"�Ώ�snk��/�*j"V���U���ۍ�Jv���bU��M������������;�Z� � ������k��;s�N�����]E����N�H�����2��v��o��os�1����|�N�?���Or���ϡ����H      2k��h��9t��6���P��R�~n��sFx+tO$��ݟ�~�])�|�� c}-�B�6w/^�D��F�-~aP^��<�Z�(��O}�S�m�6Z�v-���˴f���(�������>��o��3Π���>��:�+�p4�ݳ��S��m�g�`{Bx��p��wK���`���V�UYSK�v������ jp �N[O��o��+Z�i�m[��ʦ�����xOV#��F,}Cg���Tb��R��8�-f����읂��T��_�)(�*�k�\���������M-b���'?I������녀�s�N�z @~�mO:�$:�䓅0�`��@)��$X����`���5Ԯ�|T�ܩqA
SI�*�nn��SB���o-�
��s5�]U�яp;  \tB�W����>���u����4&���h�j�9O�m��!�>����O|�z�[�SYi��<�~��k��/�7m�{�      (dvw���:������2���XV��i�紦��W����X	C9����F��X�%B��0}�j���zr�`�B�^<�(��Aڭ���y~lllǵ�^K���"��ꫯ�cϞ=�
(��3��,wz�R,޽�x�i�۵�<��UO��D�0{����+���+4�=�T���z�LZ����� �A� ��"z���3����v0�M�6��6���4�`�lv����N!��V'��]�2�V�`D+�X����B��r-D��g�vڴit�e�����Ɔ?����/P{{; r��F9��cE���N���]�q���s٬3��x�D�0�)��$R)����TV�ʮy!S�J�S1�s�F�*����� PRI}#-oM��  p�����%��G���Y�5�#߼��������|��v4���Rey�����6�6�������]�8����~�՛�/��:C��      ¦?��K���f*��F���T���چ�-~aiJKK��l�:����Z��C�(}� ݥ���F)���ot��;������z��Z�^r�%��y���b7h>x7莎���o���Zb���X�w�)������F=خ˥w�
���ܼC�p��w��	:��v�_��B����! �� 9�]��{�lZ\�F]���6C��I�rmf�d;��Xelg�[�����G�ж �㪱 �\	Oa	Wٌ�Fu��Z����ؘnl�y뭷��7��wny��G��0�1Gu���?�xѴ0a��0)��A�R~��R��27jaw��$�D*�}�O��^�����TR���n-�$T95��ظ�2�V�H�[	  r��[�C�G�i�Ǿ}����ц��}��$�Χ�����n̏V�Bg;�.;��y�gM��߽����rq�      @����!j��H�*�QoOOJ��BU1�S�=c��%��~�gy���·�$+	?&�K���Q��	����͸���u��y~�?�8���z�����;"��~!7��+ w��0K����X�>��w�P�jf��J���;T�ٝ�C�b���;4������>bEe��J�A 聀;  ����v�ч�k�����U���VN�����[R�R�3X�4ދ�ܭ�u� Lb'V�q
�) u��ׇ5���ds��Z��������O�tg!K�{zz ��w�_[,X@'�x"-\��-ZDS�L1�ѹNX�s%Xy�VX�V�D�`���WW���0
U:���im��V�*B9�/8�c�T3����SC�{n �����I���}�r��o����� �_����]�� =�������q��-�7~�     0�t(F��hɬ�lۧU��S��\#}��a�����0����������?�ҬD�����w�=Ho�mn��:�ֹlϏ7Nj����[������+�П��g����{B� m9��E;;�b�z�TWW�:�?�v>��aB�Q�[ǒ��o����om7z��z�N;>�Q[?��QA](| x w @^JЪ���-4sh�h��ݭ���X��i3�3E+�6wsC�J��υ`���he�E+�^��^ǂ�r�>�qݏ'�s^��9o��m��{�8���>v�����oБ#G �	��ܮ��v�N9�jhhH�"Ю3'���ӹ(S^�FU�"�[
�*�p�}k{�,L�B��ւvq�V�y����&Z�iH܋ @��	���ہ����w��|��W�;ν���i۾���O�E      �:��|S]��L��[3�Es�
嘲��R����7�osOͱ��y�c��w	?U�?&d@^��q\5� {���B������4i]v�e�`<H6lHy�z����_: @
��͛��a�0<�(��a��a]#*c:ޡ|t��!v;���ώ��P{Vޡ�3��"�_��&Z�ʾ!�C �7p �7v�h[�L�`Jui������Ūx�/v���������U���t�J�݋��p����习��̩��?9��?8­�7n�w�}W�X;v쀈��'����������4G�Z�:U�*
!�(�S��,N97/�m+����.NŅ�}����A��
VUц�i�n+��{�� �0�R���77�Ǿ�[��A����?XM?���2�7��rj��F���� ��~   ����-C�2��U���n۠�]���X´t<���p��۷��s'�P�ڶ�����K���9�����1��~��;��:�����B��X�4ݹ �=C.� ��?hg�����C<�3����\'�9�����c<�>���;��B��s��=�y�	G�P�3b�,~�7�P����#��;|�o*�ߊ�v �?p ��C�|k-i��ءm��vyC6�XVVf+V%_������ܓ�U�A�*6�uC�P��h�$S���$Z���B��>��1��s^�5���\�D9r�޽{E�}ӦMb�µk׊�w���h����	nV�����:��ϟ/�k�q�������~<�"�~�]�j+R��m���F�Jݼ`mn7�T:�
�]k��
N�N��^N��  Q$
!w�ہ�����o�@_\v��qe%�󿽉.��Oh��C@.��'/��xǁ(p畧��s    ��M�b�����h�@=vfcY�2�`��?LXK�F|Ä�3T�b�}Cݐ;?:��<|��i$=D�G��̧����|��s����9��Yg�%���W���rA�cmݺ>!3�3f�@;{��%.Z�����Lst�����?��'�͘��wȸ�����q��[۝��=x��b,CȽf�tzt[�"� �� �H�H�c�q:~j3�+�E�}��m�f�k[�ʦ����`���n��vB�HXnr����c2+�/�t ^���8�����^G~�>}�t����c�"�Y,d�����5�+��*477�;�*��p�B����(���DA��&a��ܨ�Svw7�ʋ@�l��1�P�Y�r��乢�"��B���|�  D�|��n�|�7���&�ҳ:��ÿ��e����)��# ��o��p<��f������:z(_p���n������m��8   
��X�Vn,�s����m4�~��k�p*�2y��R����&=���Z}ô?ȸ����������%c�G!�����5t��e���ds͠��ͱ���q7h^��X��G�m�z��E�B���s!�1�C'�|2͝;Wڛ��R���<��e;'�P���\����Gu���g�ޡ����;��ͭ��v�����<D�w8�G�S'��8 @6 � ������i�dv/u�kl��)�*���]���(XI!J�s�tD+��&Ib��|�ڽL~E'/�����:�y�9~�q8���������l�B�7o�;v��u�����!f��!E(�X��@;?�P{]]]�\�k5o�V���̍�8e��bT�Y�2ۍ��@�C�k�K�Bu�xz����mC� P8�#�p;��G|��WS��z:�i��\����7��_�_�Y�����H��k���;^y���3���Aˆ���c� ޽�w_MW�c� �y��z�    P���=F�&̡3�SW��b���_��&d)�˧�܍���oh�
U��/t��9y��1ae"�3A�~^����E��нNkt��g��|6s����,�:�����`���;���*�BY���� D��������(�S����z��s���X5�0W>�j<�P>�O�v�v7��/��=��l��ޡN{�kk{�Dz�`�9� � "Gg������M�Tܱ����f��rÖ�ق��<1"Z鵹;ݽ�ܭm�#��X%1��j�V���:�s^�g3'�y��բ�	��m�6����w�߾}�8@Pȿ�3g���|p��[ZZ���B9�˵���*w���
��G��a��0%���mE*�Pe��┍0elc��<��\D�8 ��C�ܗ�#4i|�ɓol�ۿ�p;�FOߠ���'��N��q�A�sNh�o}�
��& �e(���|�A��.�>w�DZ����-_���mړ������~�77�Y��Α��w"x   �v�Ѫ��ty�x8�ͶKu8�-d�]���cx�����KPU�e�j��l8�X�i/1��{>`X���|�lר�yY���9v�sهY�h�8$��c�ΝbWhnzokk�� �5'NeX��3�+r��w)0�7�;/�/��Q�úF�>cvޡ������;�ʰ��v����C�_��;7y.�ܔ���p @p � �,On��I���� �tv�������F��N�2�2�#���9�n݂�)��[����d��3E*+A�VA�97�q����9?烜���e.�d;���0�mooA�]�v��w��k~�o|� ��f͚�
��s>i��ɦ��|��j^�
V�
�{/�`���^�����N�]'�Ώ�!s[�J�r���i+A�0ŏ|��V�H��  2����?�ӎ��{Ć?g�����ϩ�w��;Bw~����[����>�O��v��~� ���{C]5=�n��{9=��5�iڤZ���?L���A�   ���D��o9N��B�b;D���b,���Z�&ݓ~���ݝB�����ih-];�%&�j3��{e;��sA��fN6�x�]ٌ-aM��A.ǒ!�7m�D}}}@�������T���#��C~��GM�h���	�Y���_3��# ��lwkm7���7�v�ͥ�Z�ћ�  n � �4��h{�$��i��ṑ�N��7��F���Ħ�At7
TR���
W��+����t�=
A���1�e��9����|�s��e;�_�Oǟ|���0���!�����~!l�s~<p� ��c�{2a��3g͞=[ls��]��?01i�$-�@�}������y<��v�/q�I�򶥠�0�(PY�t��s[�ʰ�`m�4zrW%�C� 0:xo�q U�_���u߳����u]L�7綾��J d�NȽ���~�w�����Q��'�
�c9f�n�9y���ہ�	���_���̫�ӏ}�   ���m��IM�ζ���T�a�3LX=ô�!v��{�7��C��;@�#�j#���lƃ^�v��Z��A�Q��2���б�!�����#�����^ܳ5ܼ>o�<��i�ܹ�G��bMM�i�W1b�sƊ�`�jL��T�Ct;����3?�",{�Щ���)j۵���S�]Ut�7F  � "��P�l-��ͣ����'�u��
U���V�DR����A�d;����V��*^Y,w�trnX�A�	z���{���y��~�s�ٺ}!���:tHY|߷o�ٳG��y��#�^x����z!2qco������)S���ܶ�'��u]PAu/����Y���uM�E,�cA�S<]G����m+(��:�l������������n   �%��E:�e:]q��y����O]A|���� v ٣r/-)����4�~<}��?�1,>����on��U�sn*�Ǖ�U���(���  ��C=qZ���>��B�[i�����y�����d)�!����Y�R�b�&w�r�0{�D�;@����1*�`T��0��x�~����ӵTs�ί�����:JF8��^ {���޽;�C4��yx���o�7�?� ������`%�0����<�0���?�u>������!:b%��Ot��Y]�e�f�㳝whjl7z����Vx� �pA� P0��;H�6�MC�spW�H5�f�����-M�j���Πr�G��SU~��޷!�v,�a��Fu��Z?�u���<��~�ۭ)++��S�����z���t��Ajkk��9��Y���w�t��wd�iڴi��ֹ���;��Չ����?W��g��a͏J�=��A��Z�]>�����)��(J�ۇ�x�V�A	T�p{M�$z��x�s�    ��Ɍ�h��zq4N�D��^#<���Φ�4c����������ڄ������G�;'Аyqq]z�QTVZb;�w-��^��  ���S�c4kB#�9�u��,�Rx�v>��3Lq�!=�d)����n~��3T�����=ƨݳ�n6�OX�>o7Gw^�>�j>{M�����:���> {���ݻW��G.�b���=A~��w8��>"��`��"�y������y�0����+��Ϛ\��^�flO>�Ɯ�B'�P'��KU�%w}6z�N�v���� r	� ���/F���:kv5적�e�}�g�{��!�����1)J%���`�ngP�18�ݕBU©��y�5��m��k�^�ϵ������l��5�n����<����Ǐ���f�:�����]Z|�@<������9"��2$��d�L�Ϛ[�u��,6qX]���o�ǡu��5�x�l?����R�ҙ3������`��u��	Tn"U�@������H��J����8e#T�aG���bӐ0�    <k+iѼ��q*5�����@G�j���2�׼纳�S��0X����W�D`l���Կ<0|�8d��ΜsB�nnG�   ��l��ʎ	����۶�6�;5��=C���g�tO��N~�Sݭ�@�[2�a����{�l�u>��΅q^wN6����o��Ǫ����w��A��d����â��[4�Ỻ��	�߭��V��9�.K���ȏf�9����:�|a�/�@���\����G��h'���96>�f�]5��;��<�f��Ss;��E�i�fx� �܁�; � yi� M��AM��C��*KC�j�A��3� 9�B�jB{��-�n��B��qB&�Aw�k����ky=�e���~���ӽ���:��]�~ܸqB a��	���? ��w�X�������uww�G����k�:��|c����9��0:�` �F|��cT�F~]YY)>��dh]պn�~A~�a�Z��B�}�V�
�g
PjQJ>�Sv�J�rn^H
S*��CFN┛X�!NY������j�M��CB�}    @���b��=Wӵ���Ǖ�Љ-�)Nh�No��5�[p��g���x�r�n���n   ��}J"A��&��f:�b?�vw�c<C�b,'��tO�~�ݟ����/t���'�w������Y��u��չ��g3G5/��v��ָ�eo������'�eX���k.������9��x/�h��g͞����G���ȏ�{��<�����񱅱&�"��hy�N�vU������7Tc�J���T!w��m[ە��A����?�N�M�	�!  � � (X��i��J����J;��@���T��M��*^��dh-ns���:�U�@�
���)e;���݃���x�k���|6s���4�n������u�ð�,�� ��F��xX������/������M����O/�S��y�K�����y�?^kC:��s����5, �Z~�ya�7^���Q���WH�U���(۽�.X*'q�*R����[:	S��*q��|h(F�&ϥ՛�?Ʊ   |[�ݿ�2�p{�����;.�~�D��-�rG�    *�;�-��芦��{`��˩���3t�GJ0JD)���w6��N>�*�Ϊ��P��ݑbш՘�����l��s/k�:��|�s���^��~׸�ӽ�g:Y���8 /��dA?�k~Ώ|�\~d����c흃���a�{�Mx޺^���s��s\Iϐ��9B��X�Cz�\�%K�x�]���	
��
�Gr^ء�B��St
���vav��خ
�����_���Yz���X���1��<�Vo.���  @�A� P�<�%F�&̥3�PW�!�wK3�]��Ѹ��%i��*Z���V�*�vϾ�!-RY�a݃���������a�Q��:�i���u:�u���VX���d#@�AX�\�o.��|�)��t.�aS�q�`�v�✟��P�N�1���ܮl�c\y�(�K�6"�   ���	մ���PY�8��N�H[�"0��w��v`d�������T���c?  ��Ѫ�Et��y4�v%���EXr�D_���_(���tC�� �vhh���C!V����~�{ϵ_����=�����\'�yNs�Yc���5t��H���~�?���,̒�w���G>�H���",�\"˲�9�3ң���#9Yv�A~>x�_��~�k��a�ٽ�j�C��a{�z�v�o�s���D/�X1�o����������(m�u�� �� �Q���!Z�QC7M����6���h�r�n;h/Z�W���Z�6�w#|���N�=�k��o.��9�v}���z=��~�;����~��|�sE��l�YH�U���ۜ��=�v��W��M�2�q�l���L�J'�.�C��z�Lzb�8�@�   �B�ނ��q�0��W��v`徧�   `�=��Z>�.��O�v9�����_8����<Y����ٮ�]wh~��;�ɡ+M�Aw/ss�hw���z�A�����<�s��;�q[�{/��sm;d��s#z��Q���X�^��B��z}~���?̗��9�n|�!���zkn���Y��n��M��zb{9u � �/� F�D�~s�fMh�3'�Sב6s3�%��7oeeeC�i�*!�hemrWW��(P��|lCn�]g��k��o��}�nN�Ts���Y��^�^��{E�\�[A�W�Av���t��C�ʧ���j����.�Sn���v�慌-]�����l.�m�Z�    >�w��{�>v������c�\��n   �W:�㴢��Θ5���v���Tm�C�P�z^<Ä��=�3T7�K�Q��8�Hw>(mOct�/rnX�A�	{��|6s��S��3�m��:������~�R�+a}��\7J>b<��j�:��`��[L���j��3[�ݛ�UM�w�;>������ho�\z�!  " � u�l����j:�q�uo���&��Q�hu/f�J�ɽ���n|���]�!����	'���0ƣp���l�d3�i��|�5٬ӹ���e�^����r)\fם�*Z��l�j�nw�2B�6�v��v�(e	�Ũ�~�nk1����
   䚿���hׁv:�e:�n�N?��k �!��������i��ρ#]�W�� �B�    �yeg�*˦Ӓ�C�{p{�Gh|���.)����EX����T��̇�3����aw�9��\d����	Y+MN��=7��ר�yY���9���;�n��:��^���A�g�ȇ��{��N>������=_H�a��&}>��1؞��p清٭ޡ:Ю*Ʋ�=�ۍ��n;>?������ �� �Q��[c4�f6�;��:���*cC|D���Mv�R�J(E���;?�5��s�{��=)^�2�G;��>�n��\�=��a���F���@D�=���7�^"?�G�E��ȅ��{��F>E+V��úFX�v��}۝�!��l�n�i_�[VV��{S�Ϣya� D��2��������c��/��o�F�O���+� �Nl����?|�     �L�`�V��I�[��x/���f��������_(�C�h�'ˮ�7Xl��EYf��vW=�|C"��{&�Aw>g�����ָ��习�g3'�yNs�滭qZ��V�:~��{:a�>��f�>�h�s��c��\����j�����{k{�?��5�C���iO���7  Z��  ��5D˻�����г�L��!��屙�D4�g
V��uI|$��ʐzW�38
V���vB�݃��xPkt��g��|�s���^��nk�Y��ϵ�y��N�F�������&XEM��f��`��5�n=�_���ڮlO=7���ۇ��� U�ϥG�� Z� yd��)��_���*ʨP�?w.��O�Ow�!�w��        D�������tYc���n,�Rce��ʂ,�����]����ZK���aAw�\����x���r��Z��A�Q�j���uNk�\��5�z���+?4���{�0��ss1�a���6�*��mm��S�e-Ʋ��9�ھ���� �	� �1��7TϢ��Pg�>��A���k����^j���A�*IXR��kfP�3�V�\܅'U&�=���e�'~�=�k�\'�k��r���{�N6��:��f��z/���ڣ�0E�|	Wa�VA�Kt�fm��|ە��,����TZ���g���,���}�[��h���  ��ʳ�-�p���E-���>I�|�!z�        ���H���8���K�ͽ����!����Y�Xb�g���k�	3=ôo(�B�2,�mН�a�L��ۍ�������g�%�Y��:N��v���u:ku���Zپ�X"�?�l�1(1����^+W�b �v�q���^)V\x�q�p��_��Z<C���մmp��!r �肀; `�p�;N�7U�y��4�{���������f'�J�?�+u�]������&X����aw
/�n7D ^�:�^��9/k��׽F6��u���:��^����^�eX>*"ZP���x]����X�r���į��v�P�Qx��T[	*ũ�{��vǐ��qA!P�{����zs�bq�� Ѡ���F���w3��ï�������!       }��ѻ�tyc�zns�
u��Lb���$]�e�:�3L���v��_�]�u� ���h��K�z�n�}�l<� ��:�
�=
�\��پG�Av/��C���^���3�>�ڽ��z�X�?O��q��v�R,�r����x̰�3�C @�A� 0����!�X9�.�5H=v��*v763ȃ�(�6��X%�b�kc��]�=�Ҡ����0{F��p�K�=��nܫ��GPMU���a�SA	S^ĉ0Ũ��γ%��G6�-4�j�	V��t�l�	��*;a�*Nŕ�v��v[q�F���0���D�Z��   Z������Ӥ�U4�/U���:c�\��7K��       ���K�6��Σ���Qow��+4���w�]��c�6�!�۔c�����g�{�]!���;e�s� ���:����e{^wN6����o�Fw��z/���=@�N����/�@���B���v�]�7��ΥXv�v��K:�a�?T��Z|Ī�Z���@��; � �$�{�rc	�4}5�ޞ��f�J��n|���`If轘�܋�����@e|W�e��[�=��������ݸW�����`������09��QD����$,!�,0&���:\��e�1��p}1~��t16� ,�BB�&�
	�6�<;;3;������]�U�=�=��<�U����ݙ�>���mC{�Tq����S��+�4� �$�!�%�̨k,�h���v�Z���^��.3���/(��v��JmW	T�k���v|f_��qS�"���f�'��/F7�ԝ����o|�m��c�A!�B!�3��<~����;֠8u K��Z�,���^����X���:_FY/�%e���F�F�;GU\)�B]/n�1�qI�������5�o�Nܵ��f��e~3��c�������v0����f�X���d�g��G�0�4��8{&��{�\��CBHgA�;!dE���~����vL"w�``���T�ҋUA�{:dr�Y�p:�:��,�=���5�W�"�AP��*\�i�=�fN����㌉3N5V6^7G5�d��:Q�L��Dҟs���E��`պ��ϯʟ����{N�خ�D&��P��-x�)_Q���n N9�������8s��j��BړO�� ��S��������΍��q�'F������_�'�� !�B!�t�"p��"6�]�������i�(	�2�f2�]�3�w�齱��I��$�����V���϶��c��/�c:W7�f��k���F��c&��V����n2�]j���f�	e�4���Ac�>��ZS��}>%�]�%�X��G&��;gFpxw�҉��NY����mc�q��4f�Ψ�ڑъU^�{Ɠ��ن0��`"V��M��u��sx�!�'\�m�=�tN�}���#��X��y��6kخ��sڝV�ZI<'���Zi|��*�9I	SBc�����]%L٤.�M�E��]"N9cu�v��� ��p��"|ew���A!��'�~ ��ǿz?>��W��'oю����~�Ÿ��u���*��\&�Bl�����ç�y�����k^�}=~����U95��>t��D!]��s��!<c�*�^:���Ey0VM�Z�e&�t5+S�vk���B](�������jT�BY{+눦�M��yQ�u�G]�v=�X�x��\��&�D]ӆ�6�7�f|Nq׌��(ɱI�[�����L�6�a�z�O�����vQ]�|U�����QR۳==X߁��:�v��	!��R���B�Ƴ.ê���U����D���g�s3�T��p�VoA(>ĦvS�;R�4wS���7�pՌ���ү[?�:��َU���3�k�F���>g����%�Z�$Z��tc�!h��`9q�s�3�#,T��)qJfrڋ�R��$/8�v���~`)�!���053�_�����%xٳ.3���{:��e���Oczn�B�3<Ћ[�������+�?åx�{n�<�'ֺOܺ���g��lZ�
����@!�3��`�}�p��<.�:�Ɗft��ce�C���&��L�T7��B�|5�XFwu V���ͪ��J2�j��q�����ج���V�>�z^�k���۩��R�n��z��nin��u�X�ݞU�C[c{AQ?Z�	w���	�	!�����،7/	E+��@� �5����U�av�&��7��z�mA�2�����o��bV�;�NQ�+*-���*[�i9RLװY/���@+���ψ:��(�q�(XE]���v�0�0�{�f���-�>A��Id�6�����}xl�����yBi>K������ޣg�~�ќg_�_y�����I�>r�B���?�Gs�CO6��{�Kq���:뽏c����J
=!�����b	�}<�K���%}'17;�B�����Za�������3鴴f(JxW�
EFw��V�Z���֕�������؊Za��	[��['�I<�i��g�f��m�'Q4�jS��/���}���ZTG,�$al��ݭB��EiZ��~hR7��XC�8�[����3!�����B��/TD�+7����1��]h��%�"����^7�ׅ�tM�R�V^c�hB����]dr�}BCu�@kJ���B�l�8k���g�jl��9�sMְ]+��q�򱵻8���׮��J����^��w�2��)��=���$�|[

��u$qJ��༎XۉO�w��e� ��N�����[����f�o����5���'p��y#���������$C�?2\�͘�_�_�[xp�QҎ\�k#����+J������G��p�__{�x�SwT�3�_�[�ɡS ��P/��]�ŵO����P?N,͢�x����<��!���<z2����q�I�`i�X��.�cej;?�ꆞݟӁDw�Za��.��ꄲ�Za�SW�5�Wi���^��(곙�?꘸�����k���I=�ShU-2�s��_N3��85����Z?��mRs;�glW݅��ޠ,�k]Qu�u�R��:ar+�����3!�����B<p,��ӫq�4J����(�Fw��r��	T�d�h%JbPA�JezwE�PbC���	W&�����(P%adoq�V0�)Z-F��Yݡ��rW�)ZQ��k�	S�6��]fn�S�Rja�����-�S����<Vo���8��vBYN>�����s���#�}���#��_�w�ӝ��/��q^�����^�K�m���;�ǻ?t�Y$"���;7�s�y=�{*�/.������
��ןǱ33�v.޼���_�+/�To���]x�-�$g�������w�?u�Va���<�S�gnw���V^/���>��B�\�E���El^��M���ٓ�zB�X���탱j;=W±j��tc��t:S�:uÒ�(6��0�;���vqHVR��f��ev��3&�8��(�esL皬e���Y�$����^��6c;����CQ��=G1������R�v(���2�ڄb�r9�N�÷N��n&�B��	!D�+Z�l�s7�p���Ƌ������
ƂU�^��^��i��u��n&Zɶ#T��+S@�
&4�W^�s��[)^�ε�Or�l��zQ�U�1���o�NԵ���f���Z�ώ��r�VI	[� Xٴ���ʟ!a�&q!hn׉RraJ����D���v���T�v�Y5�������P��%��*���=x�;?�y�k�qrT;>�I�O��\r�:�����|��veۺq����I�~��w�'�~�����g���.ϼ|;���^�_z��v��W\���66<�_�ux���H�3�׃���ո��m�����������ٲv�?�7��6B�|O�q�� ��t1��8�/�IC�t�X^c��v�A!]������j�06�7�%e����4�CP+����^�.��$k��#��X�x��\�5l֋�~7��zc��[QG\�b�1�T?tk��ks���6�#z�5��4�Cݎ�E���m���8ݷw�uj�Ԛ	!��b��|�}<�K��ē�`���P�*8i��v�A���v�Ӂ4w��=�ۊ�6����.<"Wbӻ;O'8-gC�s��o�N�q����9����M։�f���T���-�p�ѪU�vݘVVI�	�Q�k� 垅�v�E)���.Om��.Ȅ)�8���ٞ,�l�m�
�ϖ���n<��D%%���z-��u��'Yy�����ƅ&��#�tJї!�DO6#l���w���1z����7����W�˷����Ư���R��N�E�=�����w~�B�������$nڱũXZ
�b	v���EuB�>�螮��ݟӵ���^<µC��=���I�0��@Tt�hM�^�lC{�Zb��Q�Q�wl�9�y�kخu�($Y�l�e�S+��Q�$eV7���N�6�]������v���X��a����vO����܊/���B��	!ĒGN��hjϽhٹ�X\\�T2���hUOe���}�L���c�V1���/�������/��fn���k�g;V5^5G7�d���k&��v��WR�k� e;>I��J�T?c�"���njn���4��S�����;���;�z�:Ѓ��o� ��n�1���|����YO�a4��/����z��=�ĩss �BV����s���Re�V��<\�]�����Ç��n��y�D�8	B!�A��������u�9}�������2��Q0�~UIt���+��42io������U�CY���ae-T+����ܠS�qj����1����	uu�(�E�<��6kE]7�hJ�Ѭ�90�'Y4�I5BU_�����ިz��5C��uĠ�=�`,��a��S��}dr�ur�v3���r���B"P*�pϾ�6���K�?}H��P7�[�V��Zz{��^3��ū���o V��V��(��c|�E,��=(^uj�m�16�Dc���g3_�F���z^7ӌ�A�5�m�o�e2�S+���L�
�	�="�J��nl7���2S�ij�t;A�0���02��yfw���!���[����_��o|���k��\�k#���7�����!��R����#�|��?����~�>�G��h����w|0����7]�?닐I���;��|��q���#���!�t�g
�m�Wm܅��0;��f�Z��ce�i�3��au�g]�Pot7��j���ݩ�ðD&wO���6�����Ю����7g��X����t�mױ]ׄv�Z��fR�n���v|��u��P?tk���`��gh�T���!6s�ga�Г�^Lj�g��}pdGrk�=Nb;k������s�|��vN��U��03uFlt���]Ѫ��P۽}��N�Bp+B_�{����Xw�_�	Xq������+���C��W��:&�$Ǜ�3�o���zI<�i����s�md��*C�ɘv��)���ڤ����8��R�X��*a�4yAgn����ف�𕽎с���iʿk���_��#��_}>���v��uc��{_�W���x��iB!�NoO��x�;�c��������ct
�����/�o��2�h~�_�y5���7�>p!�t����j<�����Vw�ݣ��{��i��d�p�P���EuBU��^3T�
h3Ǽ^���v�c��j|7�k�N�5�~v�ӌ�3Κ�TGl�����=�z��0Kan��
��v������r�3��w{��:�k1y>��<��!��Dhp'���s6��SCx��1L,��¢��.2�{�L���@��$�;/�3&_�J���"C�N�Bɟ�Jw�
Yu��T���iN�{����3&�8�X�xݜ8�Lֈ�^�g�t���R�J��n:n%V��=���@�����f�S!c���]+T�Rڝ1����ԉm��~ W`�!�t:��>�9z���:6ܯ�qr_��o�k��_�Оc �B�����[^���%�o���o���½������;/��'�7��j����{�B��B�T�zrp��qs��C�l����X�za:�������&F�p@�,KV?@#�]P/t��Z��T/����K���u�f�u��(u�8u�n�ju-4��E]c���PC�:7������m�b�j���y;>7�v(Ih��<Wo�=�{q�N_!d�B�;!�$D�����ѓY����P:w��� 2����#Ni��Gu���6���kpw�+q��_��
`�v���J�R�VH�&5x�j|���,P�R�JZ��*�A��K������%Z�����v��=�2����>w����+J�
Tbc{8q�&�����Z�	�8ևS{��N!��7ڋ�����xu%�U��� >�'�����G���� �B���l�����MO�X:��Ǐ���/�S����s�߾�Ȥ������N��/���@!�{9s�������ɝ�j�<�O��E&wQ8�*KT/,�ϕ��t�����[4��YP/��~X�!.s�0�z���g[�z��:a3j���;�+I�[mog��Z�Y��u�V���?	û��n��^4��°LM��@�(�v���X��G���,+���I<<;��vB�� �����0�B	w�.a�+����ų��"U&S9g<��x�3�{��G���+)�{��v抅�F���]eh�ۅ�D�B�>���;w9��Q�u�G]G�Vܱ&s���͏�V��mh�a��ĳ$?��ku�hWpҍi�`e���Kk�S6N�r�('��D���*H�)�HezxS�[	��\.�щI<p~�w;�v��	!��w�,^t�?���r<����}�Ļ^������g@!�t�����x9n��	�1������),,u���N��գ��.ߎ�/݆o?r �B���g
�cWoZ������ka��>���f������F�{�V743��v�.Z�e��RJR/���F�$��~լ�8���c2O5�f���xF'ӊ�c�hE-�Sk�]Q?�=}����=j��ol��G����5�����ކ��w�s�gBq���B�Ĺ�">�;���;p��,f�G��Ne����e�����3��(d���sc+Bw�´O�*
�)�x�No��D�RP��Լ�R�W��̵헍1W�R��:G5�t��ZQ׍B;�ϣ���!�ڝ(Z-�`����~��T"s{]�
�SPS��TC��T%�0��.��m`0�=�8�D"U��ў��s�#L��N!�ι���O>������M/�F;~��0>����uo�B!�»�p3���'J�S���S8~v���~�۸l�z��Y�)ǽ�Ƨ��N!+�����`z7^���#����vۚ��ѽ�F!�c�����eY~�{��,�}�xh]mPD�^��Wͪ&mx�;�d�j��\�5l׊�R%ɯU�k��jh׍i����X`��α�F�
�>c�[O�R;���~�w2&/¿�-"_����M!̀wBi2����Wo��2'1w�|������t����zPbt�$4�[����긆ѽ0��ī��p�%O�{I��,�������(╮�*۔�V�2��ۮc���NHkX.�-����n;����ɘV	V"�{4�W�i��SAs{�^'D�M������h�T�ąb��n+N��$i�nOo/��[��}��S!d%�/��y�?ށ���{���d���;6N`��!���!��l���9o����}��-���x�;1>2 3��B!+�|�koý�p��"rg��Fa��1�v�c��F�U���Z�LwOůF�V��k��M0�m���(�Q��'�u�n��|ӵ�X��iv�1���6�یo'�{�L�?������ZX?Ԙۣ�c�R����n�2c{QQCtk��`,Y�й/��X�	w����"!�����BZ�}Gr�~j�ܶ�G�����j[f���*��=]��F�t�yX���Waӻ(�A$T��#�w\I��P���jv�6���Q�����5]'�I>��h�����6�����_�����e�vq�^���Ku�)���7��D)o_P�%/�D*�[���u(���8��~�B��|�'F��W>K;vx��wB!+�o�`/��G�mL�-�o>{/����@!��]*⋻�#��0{������R��Za�0+����]�tZ�%��hlv��/F��^��Kv�@{ۖ��n�gL�q��Q�����ͷY'���,�Y�]j���en��b��[Y?�ĊR7�����}��'ê�-�۵��ڡ3ndb�sv�/Կ��B���N!-�TJ����]���
�U�!��]�*�
W��z��ճ7��*<�fw�V�A��3���UB��ZD+�`����yY��~]��[�J׿�U3����1���k���I=��i���ĳ���ܢUR�V;�ڽ�2��J��\��E����]����N�!>U���2c�I
���^_�]�z3�u�'vS�"�Re~1g4��� �BV����~�#w~oճ0ĤvB!����^\�v'�<p��S(z�5à���p4�t��^pj�Հ,��銮��
�y�T�p,�к@,i��фe�Bxj���)I��m��Or��8��(�ustsM盬g][��l���|���m�v3���4�~轎U?���jMj�~S�8KV;t昄byw{V�
��à�]XC�axt��V�+{���B�C�;!�,sK�J:�X�V<ws�gU^�z������D�L�$_Oi(��kUE��V���oBC
�t�`��+b��U�6�@)�����&�T�cf�X��~�x�Jן�@�t�B3tsT�L暮e���Zi$�5ie���$+�q�Ni��*W>*<���.�l����H6��*I�ab���.��y�L��}S�ط��!������.U�)�����R��?!��Ng��"�}�_v!�������(��m�K�1a���s=��S3decc5v��xj�ձ��u�X&�wY�[#,���B�{_�U�FX��k���4��g�4��̍2?�:6k��F/�c:W7�t�(��褠��y&��V��U�_��iW?\�ꉡ1�uCy�P����j����Xn1�ecn7�r���!Ln�W:�����ބ�hp'��e��B�۝��n��O�g�b�#RE��9����h��oE�Mh(8�����P��"VY���L�$43�'mv�2�t�8���c2O5�f���xF7�
1+�gD]c9L�-�`e*J�*A*hh���P:a*(R�D)�����S۽T����ctb��M�ѽN:/�)B!�z�w�
�m_/��*���2>��A!���`v~	�B�	�Й�<c�zL.���B=Kdv���[� �]U��Za����Ou�c�±��Bw��Ю������Ix/٦����n�/c:��u�f�Mkw6�I�WjPV3>�kv[(�ɘV�ڽ׉�k��u��9�ebp��ښ�m������4�_�W�+�vH!Q���Bڀc3|v&�ͫv��0w�2�=�1��ݽ�����y�"LW��p�	�ݽ�U�DwU{5L��aP�j$�7�W�%6�&5z0����c3N4�f]��U�L暬a�V�g$��?F�;I~��L_���J1�dL�M� �d�.yAdjW����5�&N�S��V�R�������V��}��=B!�KO6���W�K�I�8�Z������}B!�{��+!�;
�7��ѽ'��ݖB��,..�j���,whC�{#�V3�
����ݠ3��kvO�����p�p��i�P�elx70��k������7g��X�x��<���kخ��ڝV�%�1�f�r�e�QL��Zb�@�(�X*C��nX�����s{�f�����n�U��Ln��SX�Q�]C!$
4�BHqx:_>��5�W�������*����4��E,�V�+Sߎ0lv�OtW	XJs���
V��╍��;V$^U�,�@e*:%�����k��g�f�n��f<ힾ`;�U�v�1I��E����.PA/N��(}ꂙ0��m#�M\T6�	����^qjpx����N���B�d����m/�O_�K:��vB!�{�U��B�=�B	w�-a�w#��������=�0��k�L��Za�Z�s�a��.�Z����ٽ��:}ڀ,Ϙ�x�+�7�;$evO�?��q��I�Wͳ��[#�zI<k���ץյ�f��P,ﵸ~Ni�^�������bi���X��[p��fN��C!��	!��}�P>�����������>�L�G.V�CbU��6����t(��/Z�����u�v�X���̠.�/X�E�� ։U+ĩVSq����⬳�fv�q�����W��\��R�I&�TP�2M\���(#a�.H�)�(�^�Sn�+:��^c{� �$������_^�K�chn'�B��|�wB!�[*������V<gS�g�w����J��*�]�Up�f�J��thY��,ѽh]/��9z��F(���>f�f��S�Mj�ɼ��۬��3��V��#+ʼn��^��~hS;����Xn��&KW/�1���׳r�y��v;Fw�$������Bژ����Fq��Il�I��L#�0�{��A�J.V5��΋wg�\��
P�T���%Kso�W:s��_���	V��aa��A�j�Ѹ���������7Y'κ6����Y4�s[�j9L�E�*J���qE���)[�{0�]lj
S��V����8��J0�䅠0U(���ߏ�ѭ�}����	!��y�n�/�|����vB!�����!���L���)lَ��-b���J U�&�0��±d5Co{�����T�Y�P��Ov�6��4Yh���kVI��^��_˶'���qꋪ�Q׋󌨴����?�V�m�tf(V�OߵI��=�j�qꇪڡ��4���É�ạ���&˙;�z�=ч�;����B��wB� �}(W�sWoZ����1;=-��I�"�J���	Wn:C8��MhHi��Tw[�J�ր�f� ����$*�)iq���6�DY7�g��!t%��8k,w���R��Ȧv�E)�X�JYP%.xSt�viZ���^�T*qJ(X�b�����o ��-���"���!����ů��:i?��B�ʀ	�B���L���b��.<m�fN����u@�]��j�DwQ�Pov�����B_}���)y�!�.��m��b�_߷	�J2�*�8�X�xٜ8�L�ۮg��I=H3?��Ċ2�SB��5�h�C��)&]?��E�<�M�f5Dub{�;>;s�'7�N��n�	!����N!�}G�c�z�jlϜ���s�4�um;B�m��>�nr��W��y�������TwSs{���L��aqJ���k��J����Q�����7Y'�I=�[i���U3��c�ѥ,4�����Ȧv4)��Qڂ���T$�= J��)m�T�j��p���iJ �bƛ_t-���gJ�in�l~꒭+z��r��?B!f,,�A!�4�}g����v���Dw�.вCU3,k�<��y���^ب����UcP�'���uB�k�:�{wl�.X[�cE�6��+��g�n~����mB;�e-w]3����n;���?=��{+S{m����t����^�%��k����}5Ī�ݴf%�bl_��?;�}{��{4�BH����B:���}��0�]}S�9w�BOU�*��v|��4w��cvW�=�n:C]��$4�5)��?��4��F�
�W�������L���֬�i/�*��׼�t2�ɚI=��h����s�-}�fl���{[S{Q�T�R���L�!J'L�M�6�TE�����il'��W��T�ɛ�/���y�s.�+���y�������σ/�=��O��� ~|��z�O@r��BH�9|�P>�ؼj�>��4�g�XYA0��fX�/hk��`,�ٽQ/�	E�B띠�/T�N��ژ݃aX���k�����Ǌ3�t��ZQִa�M孠[�l�%Y4�|(����#��S?���Mj�E;>G	�
cy�����ؾ�1��?3BH����B:���� Fp�q��¬ct�d�[J��u�����Mh���S�i�v��*lz�W֢UL�����,�ݡ�w�ؤǫ���׭e���Y�$�u��^3��6��&0$���^�)�����J�����lA��]������.L��s�@�F����E�4�B���=�/��X��I70>2����yx��n!.�_��닰k�d���w��%>5Bځ�S���cgf0��Դ��d3 �BZ���|��ݯ�\ąSG�N��B��]op�c��I0�,�]�t�/z�Phv�^���(�����V��p�8�t�mױY3�����&����U�3t-�ދ�[ej��AX��D�nϚ��vE0�kl�ޙA���B��	!��g��T�(��*�]w]��3C{�Y�L��^��Fw��]gt�%ZE0��Xa�_�
��t4S�R�Mj��<���kجw�n�BVψ��r�Vq��{��]�� � ��(%J[�Q��R=e!dl�R:a�(��+F)�)�	!����W��?��e��=����[p�3Ǧ5�p��eR�K��3��e��n�j������7��rL�&��7������~�F��A|�?��󝸰�k�s�{Y�#��Z�F�6�ڎk'��Fwg��[�=fwS�{�Z��N���mw�v�]��R3��vh���:8�U��V�	��M暮u�$��h�ע��XQ�td(Vm�I�7&����n����kl����#�B�L��v{.T�;�z#���P]#��.�5�_�i�{�p��)�=�D��#T��EB���^7�=�fFw��]gtOJ��	Wrӻ^�RWĒ��+��g��Q׋�~�a�oW�,ɏ���U�dbT��&��)�Y$L!,P�B��R���onۃm&��+JI���8�����kq����B"s͓��÷�
�=�V��I7�fl�wR������7r�{��I��ן����عq�=�G��h�3��4!�����t�jtێ�O,`���ݟ� -��]ft��ܫ5�zm�`Z/T�dk�&�l���fA}��s4xO�*C{��k���%�c2O5�f�5�zN�Ҫ�rbE���X�{��]gf��Uw�N����i��e�=ۆb9׾�����88�	�9ُ�4�BH[@�;!�t!���>�I��q��fOEڛ����>m(Z5�_R���.Ou/
�դ���e��^;�J�t���U�oU��w[K4.���9q�η]/��QiW3�	�����n��M� 7e�'FI����v��]�� Ml�l%hcp�R���U�8�I�y(W��i�!��˶�ǿ��5�����N��S�x��)BH'����'�!���>W(=X3��m(�p�0��4wQ8VV��n�tu�碸^�	�Y�-?�M�nOY'�uBQ}��0��k��Ú_+�p,��&kDY/�sH�_�Vb��Y�P��g�P,�k�I�eFwۺ��~�6��Ų�r��'7�;�{pl��Ec;!��4�BH��ӹ�ы�c;+[.�9Ry���U������L �Amp�EFw�x%��fv{�*������9��%�9���cM�ę��e�(k7�٭`9Ŷ$��*#��$��{��=x��`.F�V�w#S���]kj�Ra�z�12�?��
t��w�)
քB��k�$>�?�����4��n��o�:�s ���	�BڅSs|q70ҷ7lR3G���X�Jñ,w�6��
���ڢ��]it��5C�w�6C���Vخ�X��6kجw�n����$�oE-��k��dvQ�����6�G���ljl�
����d��l=�[��i�;�۹�3!��4�B�
��А���필�⹪p��nC(Hq���%��kG!�nW�9[6��īD��oM��gub��oKoxwƸ�q�)���sT�L�۬eͤ��-4��mu���<��*�)x��'�IX��ݳV���%��L*�ąVۃ�T�ޙ;�z���NZ;�X�B�m�8>�'��ի���4��n��؃��u?!��ѓ���BH{1�X�����ܰ%�U��1��n0�%�����Xz��xG�X&�`[��_3t��n��
�}���5���g2�d۵��oK+L��V�l�@��s���.Kiw�6f��M}Poj��뇲 ����8�C���?Џ��|� 0��vBighp'�����0Է�ڒBj�(B��.�l�A�*$RL﮹=,`�ܛkvwϦ���3*��-���]8J!dU׷���ʠ�o��͚I?�]i�����Zad7����6�%Oi	Qq�)[c�wKA�%�B�$Ol	T6┱0%Mj�
S�ԁɍ��>��@!�$������^W9�p~O����E|ꞇ@������i�&�b��H!��#Ky��}dRk�S[2X�S�;?�L&[Im/xM�
���t:��!��U0���.�#���}ú2˨Vب��;3K5�t��Zq׎B��ϣ���#���6��Ƌk�Qj��P�����y�P�'6����v��(6��LﶡXEo2��v�0��142�ٵ��@��HS;!�t4�B�
dn��;v�Л]��l͠g��/�V�+�P��sD���-hxw�&�6����H<��*�>~�{H�*�S�e�jbCt���?xWH��0�����5]'�I<o%ь�I��/�'Q[�v�lml�_t
�ۘ�U�vS��q��:S{lc�H�*�����̃BI���A��ǯ�$�����B!^F�@!��3����{:�8�ܰ�����(d{�fv��=_3�g"ݥfw�`,U�0z@��͘P��5�W)j��tw�{g�c���ͷY'���zv+Y�z�rbE�ۑ�Xh�
��q�Q�������2��$�+���`��WM�8&q�\��f(!�t4�B�
�Ih�ko���mO۸���c��I��[����Q����I:C���¦wo:�_�R�uVbIn_������W���V��qL�9&�Tsmְ]3��t:���xN�5�kf���ڃg[�*�������5���{]�
T­���R�c���(�zW��X8Y��A!����	�0<�9�/��;_w#��e���1����vB!�����Svl !��)<p,�0��n�O����'�L��@�����`,}8����R��lk����q��=�����a��c���7Y'κI?�[h��w�V�bk��1I�����Q���ݞm���FvuP�M�0N0V�X���:<va̡���	!�ӡ��BH�MH
���>b��.\9���3G��吕l;4��W�6_2�"��'ZU��)�\�����(����`�m
ux���F��P]����bD\Aj%
PqI�k���(fvQ�J���k�ܳNhR������]-N����%�(��n+L9���$��qW%q��vB�^tݓ�O��
t���V��	!�+:�?���^S��zA!�t��!`��N\3�G~�(�&wY�6+X7��c�$uÔ~hS��C�b�Ѩf(��g��=�i]�O�±L��曮eݤ��δ�6���X&s��Նv�b��.�/F�ǩ°T�X���1�;=[�5D��{��F���>���s �ҹ��N!�Ǿ����h�6<cK
��cXXXP�ӆ�h%Mo�T)���#V�,u������ ﶇΆ����+dU�*q*���%Jp���-`y�)[A����4[�j�p%����P�v�%IV�L41��ۓ2������K>!��KZ(9�Yj�h���@0�;�6&6����س����@!�DO6�w��ft����3��B��u�n��.���ĺ�a��/� B!��9|�P>R�݂�7�'qan��ӳ. +b0V�:F0��f���k�q�����u��|g�ذ�]M�.hj�O"K5�t�n�(�%���H;b�η�#�k��6+C{m�V�b9��&5�j-�����I�j�1�����&|�H��P�B�thp'�"��b	w�.!�Z���҃���9w6dtO7S��4��vW��W�_̒	W�k���!�p�4��g��G�

Yr�Jnz�!(�J��#J%)�,�Y�]�$?;V&@U�۪��4BTm��=Ч�T�]֧�䂔{�
P��D�*�*]b�N�*Z�T}����&�{$���NZ;�)B�D^�`�1tnr;��B���'�)�����!_(���G�x���#��t���%B!���Rw�2�5�r�zl�;���'�v��6fw�v�n/ˬfh��N(4�W/��@����\�W8Vu��Ȋ�n�u��bU���ۣ�U�X��ø�X��p�Q7�٣��,7����l�
��cx�N�'��9*_�!�t4�BQR(�p�A�D8������C�1{�DE�		V5�Ig��m7h-\	D�T$�{X�
�''\i��:�{@�r�t�"ӻ_����-U�C*Ԟ�0���b2O�f~^�I""��Dl
�Uۍ�����>�H%��������.3��)�/(L	)ߘ�Z^*�@%�T&�|>�щI�(M�s(w�JEB�\.Z?�n�5��Js;!���=�6N��%7\*�[���ʹL��x޵OԎ���kB!�E��>��#y܇Al�؅+'1�HE��x��@,�]�ͮ��R�z���ݮf���~]���u5�(�X���	v5�v	�2}F҈>�N�?._ V�O��`}Ѥ���хb�ꋒ�$C�d�2C�I0�p�g���_[l�m���*��;�f~pn?9�ݞ	!�����B�1��!`��N<}CٹX�_���t��]gxo�W�����6��d��^,`9D1�[ޫ7���M��P��$Tɍ��5S����L��щi�%|EKè�i�'2���M���kk
~�)x61�R:a*(H	��KQ��$fv�*$Li�|�g����p���0E!��w9��������4�B!�8��o���U4�?��n0�����o����q�}�`�5!�ҩ�;�/�ڎ�6Q:���v�B�.жuC]0V��(Ʋ����8�w�}�&tv�Hk��;<}�p,����F(C��$��&k%�~3hW3{�?�$�����p{�Ϥ�(5�{��bk�"c{5C�ݻ˳��=�3���^������ݞ�ñ$��j�{}�}�ݞ�s4�3��BV4�B���\��v�#\�+7f���OW�U��$��L�:�*hzO����]���䞄�]kx�VB!�}�h'8��(43�˷5ԭ�Ώb����� ծ�R+��5������r�{���׆��(���ꐛ���T8��+N�)�6�:qJij7L_p�9I?ëVa&;�of�P�"��n��؃�����]����Ӡ��B��1���_|�����'K�u���5?}��-?�5|9�%�燾
B!�p�_��7��j�6�TJ�env����B^3��=s�5C�"Z���������%�7��&�d�f��	�
���K��D6�{�k���X�`,�:���.1�;s���D�j��ݞ�q��<���BV4�B�Lc;�~lىk�*)�d�u�J(b	�+YJ�R�&4H��A�k|O����M�a1�!	�*$by�)Q�J��Yhl[l	Z2�Vc���6�W�Q�Gp�A|j&I[*���/#�t}F�g��Z��
Q2q*	C{�^$FE5�{�R@�
'��|��ȸncn%.�)�(�����þ�a�Y�F��!�t;������!�z:O�Z��q��!�b�cr��?�>����g�I�q�hr��\����a"�|����?B!��������Uy����l6[��j���mS�Cm)O���V�Ɗ��Jw��ܻ����>�ñ<�m�p,d�>��]_wl���8G'��b`�����k�a�����{mSOl^(BuC��]\K���D�����S7��h��*C���.�!gL>_���A��F�w��9�D�bB�J��*��Bڒc3|q��l�u[2X�������f�v�p��.2��S�S�kٖ�jӻ_��9؈X�kibC�F�2�E/�������;#��ޤ�O�hl��O:T��X��]�/�E��Jl�]��'�垛'N���p{��.�����L�R��m�*�@U�D┛�>84���GҘ�˴vBYi?K�8!�����x��?�����O���o��z��/�d�C=��������!��88W()�d6K녢�a�-X3�_7�c����p0V�P���R�{� �{�3���r�Di���F�>	^�n��xm�L�䠬f�@u_�����^�7m�~\�5EUm�=C�̃��;=��%͎϶YZS�4+���1��L��E,�v�BBY���N!$Qr����1)�`��	<u|KSǰ��'3��	vF�t`{BW̒W)��]$b��+�	���n{:{�A��v-Jx]����M8͡*8�����G�7C�5��x;C�h�8󛏍9]=_��L4���^_!���{�2��LM��k[C�J�
����!C{@��T޴���]gl׉UAQJjj�;��\���q�Q����vB!�BY)8&�7��3���{9�w�������4���8z��`���9���?����BV�z���q\1�C~�H�^(�ZV'�ޛ���v�n���B_�Ц^h_+���	�7�6�����z^�Ɍ�*�L�Y�ݩaH�x�J�r�����Ƅ�����͌���tufv������C�t�Cq0V�nhalW��U�DmZ���2����3�4&6��s���!��L!��B�ƞӹ�Aov3�٘�ƞY̜9^IiH��+���+`iīHF���� �\KhxoM��Lī$�J�;�bV��v��F@ਜ਼�K�Q��1�D��2'l���,���.�W{UQ�g�ƈ�ebS�^y]�Wؽ׆fv]�I���]��`bh�R�T��v���I[���j|�hg�0��B!�BV2�|o��O�C��7_��UC����_��O�BY��;�/)�n�������?7��ct��fw�u"�X���XI�ܓ4�k�)�p,�4Kb|��냺ڠ�o��wN���l����cb0���~=q=0�@,��=0�& +JQW+���	�2������K%�UIhl�����k���v��a�����<:>����~���3�B	C�;!����T~r�A��H?֏��ի�Ν���d2Y��}���uaʻ-������n*b9$ep׉Y��ꍱ�]�X�{�7���<�T,2����S�D�Jm�H`=��1V6��05��j�6�*1�='ip�nl��BT�2�{��8�v]�H��R�4��f3���G���#Lk'�B!���1�����������\�t3_��Q�z�C �BV:�KEܵ׹�Ήո|"����X\X��b���@]]P[7ݽF���XqC���Z�c	�M±t�º�����6hRT���z�x��-�h�g$]�F�0,�q��P=Ѡ^(�K����u3C���X��v_���v�nϽ}��ۈG���N���\B�C�;!���r|���g����tmO]���c��s>����=p֙�e�+:�E���=lx��M�+�������,�����{��%}J1�+V��6�������X�3Ë��ϗ����<{q�[�)<_7^g^�iE�ڽi����4�!��]��P��瀹]jl7��+��$�di�θщI�(��;�
ȝv�nL[ �B!��<犝8��?Z�{>yQ�����۴I�́S����7B!�Ϟ���B&�Wn����Y̞=�\.�4��5�[�C�B�N�㻿�'���[���e���u�޸>hXԙ����Ў�|
�Aͩ)FC����m°��e���������D�qk��5����A#�8˭�k�>C���]�ebl�����58Q���;�|�X?$���wB!��#'��#���\�9�u�)�?{&�� ��gK��䨋X�{J%b,�x�>��w0���c��2!+�}�-�iڼ��pl��Peon����U�iV��e�AqI�f|_k3�tF��9I��q��Sz��+PM�r#�IR�L�2��Fv�UOiS�C�H��}��G�9�E)B!�B!z�$���J�|���&��x��?��� �B��B)����q�1>��l �g0;=m����n�h�0��(�=x��
�ꄭHvW���x���*�{���*k�A�g�iM�δn:����x�?.��A�`a�@��u̍���i_�v�@,�0dj�E�DO�дVh\O���C��XX��<���}�ѝ�CB!v��N!d�Y(����~������W�$L_8�s��@��3��|	2�{�6��	�2�{c�_��wHB��1�{���4��{�i�XFm�>����k|�%�vEfN��4����6���BT���>��mL�"A�onOX��U�v���'����3ۏ�����)B!�B!v8&�_�����w�Ͼb��������� �B�S�Eܵ׹Ǯ��x�x��cX\X0�jB�P�%2��j��ڢU�0Z-���NhZ��_���>�z����f�h75�{��R��x�:m�]V}V�������^(�������c��~B3��.�%}R{�ڡ��.2�g2iLl�޹~<pĭ@!�D�wB!mž�|�pD���5���W���u��(�]`z�	X"C�Ѷ�³�ɽ��nfh��٣XqD*��]3&t]m�ߋڂ�y�8o{P3�2n�	
?Q���L�CO�hh��MƘ�EcTb��.6�{�%�(U=�)�e-T�"S�̮��&���|�����0��p�S�W��vB!�B!�XX��������ϼ|;:����wp�� �B���3��B_v��1����={�R�Ig��P,U���쮫z�}ie�P`v��e��t8V�s�ڠ��%m�z�uH���g��]�I�`���	������%;����E3����b�ñԻ=G�!
��5Co�X,T��kq"?��<�������!!�����N!�mqūLj#._����,LG.�'5$`r���Hh���f���=$b�c�X|Xܒ�Y�8۴��f���Mfz�{��k��Dka*e=�:JA8Z%<Iƕ$}Z㺤-��`"@��L�D3�W?S!J6޿e�����F��%7��(YH�Ҙ��BV��qc��#%�NAQ�B!�BH�8&�_z����^����-_=~�4>u�C �BH|�%|㠣Gb��"\�1���fΞ���LC�du����Ʋ�	Znld%���Y٦�Z�a�j�"��M�b����z�st�D��i]QSS��ez��%����P,��]���~���]bv^5�����#��^�	!�$O�*��BV�����@��Vov3�٘ņ��p�x�[:m`vX*K�������^,^5�MM�^�ɤ/h���9�����鬒�#�v�O �Ȅ-�8� �K�z�|eo�`�#듭ob^�]�R����1���Yڂ+DU�eb��ܮ�:0�P%2�������R8���:��B!��9{~�f06��k���s�!�4������A!���b	�T��A���5�W�)̝���
�I�2�{û�v(�JL��Z�����p��k��5CemPV+Ԙ�C�:��F(��ψZS����(�X���<�qB�Lj�&uBU_��<Klb7���&�X6;=��&5D�`,Q�0��chx���w5�?�������"!��fA�{��ߛ�P_z����`_������\�Hta1�Ky��|a@Yٔ��JRC/������13u�&�(�+�uPĊ�����,���6��U�2�L�T}n����cԆwXlU�:Gi�{-����D&Ř�X���s\S���FOQ�=cJ�f3��O%>����T"��>lf�R��F���.3�Wۋ�k�06��S21�����TE��S�1�jz'���4�Q�"�B�
���<��g��C����}���9�w������ �B!���L�q�^�j6����\8�s3�d�Z�{��.	Ȓ��m�����^�Jk���wY8����6���-x-��֢�d����΍�U�1X�3�dV����nږLQ����ܓ�2����fv�`,���P������3Y�;ꦴ3���dʯ��z0��S��ɦ�ߓ��|�r�/������Bd����8�q׍b��1l����ym�m�`Fz�ۓ1Zk~)���05���.�������=>�ss� ���¹���Ϲ���(�\��dzsS'+oڼ��:c{��+`��eFw~�{��4�7D�ƽJ�r�&bAK$d,��JT+�u�{Y��=4�:�z�c{��Z2n����Q���T�k��LV�ڃFv�����AA�.D�M�k� ����*��=dbטۇFW!�7���bߡ<��&E)B!��\���}����u�n��3���{+��i7>x�����1��=GςB!��Oʇs���ۀ�GQ�;���B�d&wI@���nS+L+j��0,Q8V��Nh��uAXfAY��m_��&��v��}��,��RT���P��b3��k3��OnX����5E(�d��j{�P,�Z�i��6kphZ���������<!�S��V��[�c�Xճ�xxǇ�*;�:�&��?���-bf~	'��^��Ss8vv�N����J�5i4�7�գ�t�.�:�'n�EkG1T��q��V��I�'B�S�������#�ǁӘ[�BH��$5�S1��c��"\�!���pa����aKez�km�fw��]ix�	RRӻG��Z~�J�.��4����"aKvW�j���� �Ldb�����zc{�J*@�Ũ��]����mJjl�'-D1�+�T�vs��q\��N�p�kf�kFB!���ǧ*!�����B!�BH��ȕ�t�j-vMfp�x��Ә�'��-1�'�<���~�{�>TL��B�cnxW��eF��L�Q�u}��&��FUC�jf�5�vhcf�^�r����ݿvx��`��[7����:�A�0r�0B0V0�}`p��I��Ã�r�g9��Y?$��?��4��i�n��;7���k� [~�51�_9�����E�?y������O��Cgq��,H2��� ��\�s��x��x-6�-�������Z[9�L{�M�{�����x���c����犸�`�|Ջ��<mcz/`~�$r��\��������e#\)M�A㻯-�Ԡ2�;��-��Zntw��}ɧ.�ڣ��M�4�f��EmI	Vb�r%ik���E&v�}H|��I�>1�#^I��Q���hWR���:�j�bj��X
�:��"!�B!�B!��nd��B�p�Vc�u�t����fΝ���D�0��=�V3�7���&�c�j�~3��6(�O>�=ʽM�M�9�z`�9I�
u�Qj����Ѽrj�mk��6QV��.6�B��E�n�I��M�����A~`5;׃=�r����޾���B�_�;׏ᚋ���'��%[&�ͤ��c�ɦq�Ʊ��]Ti;7������>v��>Y�'Ѡ�="�ϸd#�}�f<m���?�v�y��~���O��B���1|���+�<��M���f����ރ��^�e���l蹀�󧰰� �D���he*V����߰�Ml�S����CFw�hezV]G���n;&)L�,՘VT�s�O�Yeh�Nac�8�AlbW'���Cfw�%�d��&���0����(��;[�3��K������#�B!�B!���88](��*l^5��Lѷ4���)��]V#���5���FwQ�P��r�8ؘ�eFwy�����F���]�n��J���e�Q녪>��=x���fv���Ԏ�Y=hf��	C�C} ��NhSC4Ik�������\���f����	!�=q~�:��_�Y�n���~�+cC}���͕��}���S���W<���/��C���������W_�k/^߶�v��=��+�V���\������cG��2!��Y̗�f�Lj3��&���y�,Ma��tE�Ɉ�(���R��1��S��	�"1Kjl�E�;�yU�
l/4�7�+W!�J�fs	Y�>յm�I�͘����U�Lĩ`[T3�x����8�(QJgb��GQ6���M�Q*�!2�����A�����|?�?Z��ch/�B!�B!�B!���|�p���.�(a�0��sN�{�W+�d���~��=��=X?T�E�w��]w ^�{�Ψ^(���񪳹�=ʽ�M�n��
�������+*���X�Zb��$KQGT��XI��uDU8�&���M`6�
��u�\s;!��/'�*��7]�kW��p^{9	���k/x
9xw|�𾘣�C������Q�F��o#=x�5�+��G������W<�oBȊ�P~S���|�p�ƱfhOY��dzΝ��RQiv�z�L�*�*���4�*Y���^�����yϦ}b��:(0�����6��L��^ӹ�^�'�V���mz#�(�]-Fy�.�ٽ"Z}�A�)	�{��+:9��Iu��ڇW�B�w�g��Jǝ��!�B!�B!���5���zGq����. 7��	:���n��nW+Tރ�((+�����ʕE}���n�e[lg�{Ts��OdX�]����EuD��]V��{�EE�Pdh������^�4�G�
�S{OoW�ƙ��;Z��)�kƝ�	!��D}�%��s�n�;��w��t���)�&+�{�Sq��������S3 bhpW�y�0^���xo���p��1��%W�-�
�� >��Ǹ!dEqj��{�9W���n�e��:����i,�ϋ��&"�+,Y
X�fw����R��bUX��o\��^iX@<Ѫ:_צ���ٴ��%GC3*)�K�6ս͵�,j��nh��Ae��(���b�F�j��=���
��'ë&1��C'S8q��ω���;��B!�B!�B!�dn��	:�Lj�o'���iy����R��^/����~ӻ�(2��{�x��r��nۧ��c���hr�5��k��uD}Qox����=u@O�0\W��Ek��M�jC���!c���><2���$����cy�O9_9��B:���,n�|3^q��e�0����,^��x�;��ޓ��w�໏�xr�����~�<���Za!��e��ċ�������o<���EB�Jb!�w$���)�X�K��T���y�N�Ep{Ba��J�
W&��M���]D�@JCX�
��������
R���8�uc��>8^5.ܯc���jI3��l7����'��Į>����u��&4�������dr��^*����(Jc8t��!��(b�!�B!�B!��8����NUt{��=�f����N���Y^?T�	E���
�ҙ�m녺Zbr�j��>���qofn�^�c���uA�����v���j�g�Za�����nXO���02>���*��dG��;<s�gBHg�ߛ�Kj'^y�0:؋���⪝k+Ǐ�Ň��#ܷ�H�=l�Ư�t	�u٦��� *�=���]x�5�+� |��af>BYi�J)��5���1\�6�-9���a��4���-�"V*lv��X�"�0�]��0�#�'4�{���
V���н�����o��)�_{��[��6��ɡ��c�}zs{p��ϟ�P���E'wl��afكb����1���-�p��t�Ts{P��R!J�_KX���l8�A<|*�c��t�#�B!�B!�BZ�w'�ޭx�,��/ �0;3c��nb|�mM�~�{�@�@�PT�E)�vY�구.������}��ă�*-�1��R�킱Bf��C�aX�Zb����n['�bnW�ڣ�bUR�GGP����><x���s���=!���ɦ+)�y�16ԇ�Γ�L�}ox>p�t�#���thpGuk�W�pq����!�z2x�3�����"|���/|w
E�@Y��犸�H����Ć'�IcM���Oaaa!$b�j��R�r�����njt�U���av���'j������@�L[���^�n��Za����?V&h����{��]|��j��5m!�/@����$�uƚ�m��&"�N��m'�����c�ό���,=�C���b!�B!�B!��.�-���CNM�|�ƚ��x�Dk��͜�
e!X���, +n V4��:ˬV(	��d낦aX"�{cL�O��oS��Z���X��`��?.z0���kV����cIk��:���hr���I�ۍ�6�X�=�P��N��a��B��랴o��˱qb��S���_�����c��7�� Ǧ�RY�w���چ7?�)X�¶6�ed�����W_�����%B!����ί�Lj#��&��9�g0;=U~#�lQ�7���Fw�uRF���U@�
���Mg�P�B�=`x��i�aa˗����}��{Y[m��R)�ar#{h����+�"Su���~�5���New��⓻���.����o��m��Q�^1����v�����02:�|�(����y�ܿ'G�JR�$�B!�B!�BH3��
��غ*�'���
�?{��Vy���-Y�{e/�w	a��B��R�h���Bi��Z��(�m)�z[n�C�-���=BȀ �vl�{H���#ǉlK�lI�����p�y�<r�ǒ�<_�N��6���=R���s�0Q�=��a*k�Z��Za�����q��kzI�����>������m}�������-Y5���K-���| Űz��'X?���3��(�.=�S)�����@�-�5��X[j��U���84�.p�7VΗ��}[2�LL,����Vy��-����p/�ˑkV.�����_��/>F��~������� @����M5AeS��b6�ej�Y�z"∶K{�>	:�޻&�����8N|��P��米�]�w�1�%'�R�K\�=Q�=�~��{�?�y��TnK]|��m-�<����=ں��S��O4%��
��������CކZ�=��dS_A�>�������J��}A�l��Hî�|        ;��ʦ��<N�XdTN��M���(C?a���Á�jtҚ��WO~����6~�Y�Gؽ�}
����#�<̞��`*wMdOt�h���������� �I��Y?�c=�`�}��}�r�����h
��z�!�ܹ�yd��&�C�ѭ( LF��\2I�|�L�[M��X-&�`�4�̜��'ߕ�>���d���_W-�,�8Sl~PC}O�7V�O,��?�����Z  ����XR6��.&�(��o��ިx��k��`GG�2���{'�'��5	5�
��{�<�u�����Uj�/���}�u�%>N~��(N�;�S{!ѭ�g��	O�	N{�;R
��?�`:�:�P{�ɦ��u������6U�Ď�;5�`{J����d�	���"ǭ�s�&`���#���hg2
       �C�?$���ȍQ���i͗�E&)w��i����غJ°{_A�T�x��t�v��N��=�x}��5Ã�ۺ_\�=�5������L"�D�n���7A��h������{��P(+>��|1q��ۺ� ��Z�&�Ǉ�5X;LV���46���(��ФU���E2�,W08�
\򳋎��^�&w��}	��j�#*���ɷV-�%SKCW�˭_X&ϼ�]���z�� �\8j����ʦ�uާ�e�7,NiK������L,�O\%���#���D�P'�Tڄ��;�Mb%�wݯ�4�m}8��<���a����6$���&	��ݒ�-�� nB�`{��	���N��C뉂�]������M�ɩ�����ړLJu�7~S?�����䖪6�l�I���;D�       ���-���t���nv��"��r��n����ؚC�Za�uB��c��^�U�]��m��cG���ܧP$+�~��$X/�uҽhV���}��ِ� V�A϶�����>
`�O� �ą���[G�8��놩Vp�V�s�p����k���ϑ�啈�#�|��:$~���[����+�R�Z��sg.�(&�-��)[+�P7b��w�,��&Ў�"�b�x�>:O~���ew]�  RV�a�e_P��3���K��$��)��l�����@J!�>����hKGeU*�}�':Nm����7$������{�(ڐ@*�U�>��I��G�8?\Ov�;��T'���5	��]�ɪ�ǉ�����s�N�9s�M�٭i3�5a	�G�w��        }S+��[�wcg.���2��$��a��[���A�@�����궦�O[:6�@�����?q��T���w�jH�=�h�u�h�ۺ�F��|��b*{=����-�:a��Þ��Yr�y�3�dO�I6XCT��`���X��5�d�a����"������~ ��������K��:L�|���/�H���^�󫟑�=����q�  goKX��#�=�+�W+4�XOD◈�EZ[�c���Ǉ��	��tO%���p[϶����{����J������$>,��~��{��֨��gx=���SZ'���s�)Q�`&�������or����
��O@�:��l���A���f�؝�Xe���E6�F����rO��        ����n�wu�5��\�\s@��Vikn��a�8V�����5О��a����W[l�y�Gہ����zvo�}��:LL)���`K��R*����~`1A[*k��Ǚ\7Li1��a�}|��۝.�i����&�l��HxE� �lS�s���K�4/G��Q�8u���/?�m��r(:��96�\w��tZ� �����s���{~���ܦ�A; ��#"kBʦ�Y��@J��2�k�B�Z�U|�M
�zOd%���U���ڵ��0� {���P�Γ���x�~�0�޳-Qp=�q�!���2A��-��3Ğ`"�@���`{�I���(�{�r{$bsKc�&�Չ��H]׳�D        Ȍ�MaeS�L��rZs���:;�c�����=��X���n8��{϶���Ֆh�_[��Άnߓ�`|�����H�z��5%.���8�uî�@�S9J�=�:b�������b����Εc��̲�6*�{��� �I����g���$H��sF���\��W���M5�l���㐛�_�42G�E���ɘ"���ț� h�{�wwl+u�d�� ֐�"��I{[���='�MZ�0qeL�&C�':�~0�}���>���ݓ��S���٦U����DP݂��ݖ �?��m�ǤTgev�8\�Z��.V�i3ʦڰt4v=/��'\       ������I-�U"��L�X:�j_K��B݋cůfr�0հ{_����6���:a���E�k�}���n��-��YOLV+�zb� {�uD�8�^��s�>h��D*k�����g��X O}����r�����}�P��^�\nx�5ٰc�Jɀ��R���eR��㘙���m����� ���л*'��9Jd|��@���EZ[Z�OX�q�k�*���@'�DR
��w<�}m��'k�z�dP��j��| !�T���4���V�9ի��`{l��"��Dm.iYeg�ȶ���뺞��PY        7��!eS��J�	�cE��h�֖��k����ɂ�����ZO�*�ߞ�8�����O�8�y��D��_�k�];��8پ�x0����!�!�8V�:a�`{���0�ͮVf�H؜s`���D뺾g���/f�Q��j��0o� ;<9V��EG�-��)/n�#��C.�>ut������
�k�������w�Ij�} Ȭ_$�uR��c+��f)���i�9�_{�t�}�'�����$U�aw��m=�Ed����z':O֖�m��k�j0���㡆�S��u/}OLI���&�������X�bW���M�}&���ڦ��:��       ���{q,{l�u˄\Á�Xa_����ű$y�} �CY3Lp�/�>�uC-���\3T�s�0�x�놉�h�'��k]1ɚa�0{4fw�s�Ø#u�|T�����îc�@*,f����r��rAvY���9G��O�#ϼ�]�T�}��b��%����?�����`�/j
þP$��D[B�H�����$�٘k1�s�c��b�x�E^�2��wc��򋋏�o�ϋR��. ��j��;���g���+��:L2�m�gT���X�>	�����&�?ލ�&�zNf�:1�j�]$��{|{W[��z�w�$��S�$���b��g[*�Pݎ{���%���'�"�BOj���p����X�!`�]MQٵ/�ܧ��BUv         U�/,��M�Y�e-�q�F)sE�m
�9엠�E|����k�n�a�u�������s�輿v-�c�0�x�����}�t�0ٕ��%v�#��9�1�]2:�)l��v�lkI[���5]� ��`(Ԝ�.X*s'�p���Ե�C�M�F_G�)��i���Ñhk8m����f��e2��V��e1�^�-�؛�t�-����Q�
�Y�@lf�<��'2��$x
N.���[*V�I�����^Ӳs_�����ۑp䅊����`����~��B����1N�uA�ǱpR��Xy���Qy�S~��c��������@��	�F���ؙ�V��r�%2!�$Ŏ�䘂b��%�K{kKlr�8�J=��Ez��y�&2��+�*2�r{�dRIo�?����q���T�DS*ǉ&�����Y	'��`��s�ɖ#a�MڣV��ewsT������5��_�  @���f)�Zēc��(&���:BQ�D��-${�����\�IJs-��1��j�����3��QeklI�2F[����$ϥ���ƨIlfe���1�T�hD���J��+t'�-!c��5,{��z^G �ε"��F��3��3Gl�(�����r�Ar�!�E��h�֖�ߓ�5\7�-�%�>\��q�%kK����~��d�d�4���a?k�Z�Jh�����՝��i[��g��ui�uug�� Zʱ��'%3����^��TYߺ��5�v[G�s�����W5��k��iv����eq�˶hl�kJi��":��
r�isc��~i�g�D�}��B�Ig�v�:��{��4�^nl������?Pq�_�=��QC��=��:֖�6*7�h��q��!�}��ƽ�Km�O  �C�?"�Vu��_M����%ϡNj�@9��C␀D���oo�`G��dS�Ė���`�I���$�K����Ie/7qߖ�8�y��$�H��z��������������6��<��T�ۺ&�ԉOu��bWC�v�P~=m���%*����O*� p�Pm�Rf��csd��L(��M��/4�4?����]>yw[��k
�cb�Mf�ct�C&���a;?uя_X�V���>ٰ�M*�z2I���9�������:�#�u��=,Uu�����]�2FuC}�W_;g��|U_S���4M���M���{�{}Mc  �pT>�+[W�=�9,E21�(��%��(�߄|���;|Ov%h��&���*�5��{W[�}�����o�;��O��DfВ��`O�n�3���z�t_7�/�>�`{��]�="6{�؝959�C,�4Iu��*����� �f��|�R݅�wֶ�+����:�hln��m�:w������5[��������;:<�麸�k?~��	n�~&�.9y��ay�Oe���i��c?,6���_�>�ll�����:��]�bo&�����\w���Jr�S�sOS�rH�����O/:J���il� �����Ķ����\)r�b��|GD����s4(��_:�>e�Ht�>./�W���z�w{�}?Ǳ]��dmɨ��J
�&��(�j�=�C��>���{lf�Y����v�m������7J�Zͬ9,ц��� �P�Vi?~�W���B����2�"�S\���/VV���MM���V	�S��s;L�9����<�^�8��X0����B�to����Y^��"� �٠V����in)e�Ʈ��h�+�]��\������8y��J��剽�{���������}�8���1ڬ�׷Į�  0��������<b5��:MR�4H�-"nSPLa���������h8�OR+Y�=��¤�����%�'�s�4+�/�uÞ�IlOe��W��}��)����Y�]=�Z-bw�%juJG�� V�2l�7���������D ���(7��T�N(=��������-���ʵ�g��|�9o*;u�����]��o���\<�<o\�v���|���������hX�$�*p�-,�=����-��{��>W�����Vn�b�{��L�����<{t��{�'ϵ[��m[�V�gG�տ{A:�\� U�m��v�y��~�*O���(�Y��\�������K$�!Ae����'��WzIp��T�����R�}�yl�����N��z�������;����j?p[�@��sױ�b��!&�U���$�|}���R���ְ4w��rS��/8�* 0y�r��|9z�[L&��Q��6���,-�g�i�g�7I��[F�68cQ�,����1��Z�ybi����ѿ���|�3!�e��ϗ�f���h2���m͑����(c���{Fx̲R���t�����������m͑���{=�   ��@HdgSXٺZ�P�+�Y���;D�֨�L�� |���������',��J�]�n�(����}�ǵ8��(�������
�S�'YK�3ܞ�PVך�2 �*�&�C"&���f�M��Xu��T�F$ج��nuv	��ިos�Y�P�R�կC-D�~[��5Ϳ
O���sO�śF�E���7��7��R�����
֌*pٳ�5�W��֪����7>�h�nMۀ�'�*?��H�:mY�j�}��?����֋o�fm��؍��|D�=����<���w��c\���M�'7�s�\��W� �@~�W�O�{�~��Z�ڿu�s� � n���AxsD,�Nx��	H4�p�#V�A�Iz�c��G���e{�����v���Q��rOi��B
�L&�����&��l����%(Fi��C�%��ף�Ҕ(�^  #��(r��\�ܑb#4�2���y��	s�����{���a2�y^9{I�8l��r���FY�4_N�㕇^��De�/-���^}�s�
�$�u���\����z�_{d��-��T����9�PN��'���1
  yj�}[}H�uk�*�匝yl)v�(� KT즰X�1FC	$���U�Pq��*���|[l�ߓ����?���n8���Ű��\W���v1[�b4�$b4(���a�}��T�FzT`�" 7~f�?wL�?���O�}�qe�7_���c�]y�ewAEE�ֱO�p昂oL,��$�9��?�X������Q��ap���S����ml��q���v�~お��2��|ٚ��������R�����KNp;�_a^2�T.��l՞bR  U�IDAT��o �d|eKtKׄ�Aꤗ�n��(9��8,"sT����e�I�e� !�F�$K(�����Z�H��S�����&��'�dT��������:p�ߍ��4��h4vN"){��"�Y��D&�o�l��F	��V��HkG$Zo�+�KT��}5��  @jFX��2J�cpJ����e���fy`]-^5V�(c�D&�f�xʰ�V����9|�K��g���Y�֒���JeBq���w���1:�S�S�h{��j�<O�e2�����R�Π��9��?�U�/�{=  �ԫ7w����V��-�@�Z +_�ԵA�%*9��������DC!	���!	�u���������.}ȒԊb%]74 ��d�0��^!�~�{����:6�Lb�Z�d���d��5F	�Y:�Fi�%h�F�{U׶�J�	sr� ����c���Ӳ���pD���v��*�z�k2�TT�	������=uݬ1��5�����בc3��,�+�\'u-�'�<,�W��#��f�q����������W��,�؏.?}��;��w?4il^ޣGL+�k4d6�f����Y��� `��&��O���o��}��GtZ�b7D-:�Ĩ�=�ay�r`6E�}T�qT��m2t_ 7�)n�)�-6�Y����j#Q����n�	D�����*����JiD%��զ�Պ��`������9��*  ��Q������J�vM;�#�K�r��{��! ���r�)%�"�&Nr�-珑_>U%�j:C�h�S.;����9b�+�A�ە1�s��ZX2�%_9����9r�2FK����=u�Q  ��t�J�._ �}��f6����wYE&�r7�)[�Se%,�HH�:Z4��Q#�	c�C��D"j�,�
ս��������MZ+yQ,��X�hP`�cՍfuo���iPW,1�%��R�`E�W���z�f���kT�:±J��Q F��e�r��Yy�U���}Z{ፗ�~R�����[��-����/��5��^�5�kE�T��$V�=���.�~��1r���v�U��f͏�X��Bn���O�ݼ�y��œJ�W�vf��q�|�to�l�^�>  ��I�@H�_��J�<  �0s�\���B1�mהZ	��猒�=Q%[��Ou=:z�;�T/�	���r������+뷷	�e�^��\��"?8g���齲aG�`�N��/W�{������u��'���J�   @��Ԇ�R�����/������j�� j&M-������n�Rh3�����u����{��tDcű�����I�u @������%b5g��Ac[G��-{�k߾��+�#���k/>�o�����Z\�d�S��/��2[~��2�����|s�>f�����w��{��Na7^��V�����J=zF��Sf^����?�X.���#$     `�:��9�<Az8�&��Y���G+	�����Y��3Jc���F�}0N]�+������j��o�Q&�=UE�}��X�'�[V H��(�]].?}�R6�&�  �G�Օ�$���<  �u���Ii^NF����n���.?}��n���n��w=~�Q�K�+�w�2�ث�LR~�6��6w��(מ}xF?	�����͵����ޖ�������P��7c�K&wT�K�<m���ѷ     O'��n� 5�����r��{dgm� uK��	�g��d��N+�}�
��l�[�=�p{�Y����2���=|Xh����%ܞ�؇����?��5��    ��X�t�,>�4c�����~�o�{��W�q�e��x�/~f����O)���ǽ���yW�T7�Ȱ	�_r�,�T���cE�QymK���G���U����Z�=|����>����	�c2�'�+on�+�����B     @w�'8��	2#�j�Uɾ��]��ZX*&����	�g�U�,S��N�k檍��6�.�2F3F_}�2F��S����#~���Lqؔ����1��c�    ��_⑋O�����^��{ss���\���0�_��^�����{��Q�ح�u;mf���Er�}/H$*�5,��'˪��3�X���?�����/^u��`��**��k[���gf�>ݘ�����>_�o�'�-T�    `�(p�	efA��"��Dn{�J�:�|���(W�R�,��qٍ����Ç�H8� ��n��~V�F�h&ysLr�2Foyd��q�@}����hf�Lrթ%r�c��Q     �1f�A�]�H�fcFﭏ����޲�ƫW7���O�􆻞�˱3�-�ͱ���f�+�5˦��/m��}�]�!���yY$ml�<�ޮ�o�l՟RQaPK��q��<����/�Ŕ��s;,r効r�C�     .�l��o��� 1�r�q�<�nC� �?S,E^�O��&����������]|b�x��0}�CV,̕���kg���IŒ��>f�͑��y���6	     @&�=�0�\����zus���M'-؟U�n��̧����,�U���b�#ݏw��3�M�RY�&z��Ys�	U�J���4���oϩ#����Kg|7t��'����9�58v�(Y6�\^�\)     @ߖNu��1i�_C>T���q���ަ�v(�4�s�H���y�ڇ�R��6{\�,��ͦ�K
�Տ�d_sP�ۢI����=k���[ۤ�5$      �4��%7-��F��v���z���[������}r�/�8}t~A:�f1�7�\ ߺ�E]^-X��	%�X	�t�^��{������$t�WV���������aI�'�v�\y��j�X�    @�,f��wLZ�Ր��$k�̗���t�^��e�ʐH�l2�9G���O�tgT���
��jQ��Q�g�=�W���8���a3��er�?�      ���r�X-齒_(�����^t����n����_=31o�;�hT:k��"�̜1���]�7��_v�l1ӻ���-���=�n���M�>�xɪ?D�z��E��Lc%�"�C�9z�<��     ��Y�s�zji�8n�G�|�^�[)��I.]`d�.[d������LuIYcT�8�%��j�����;j�[
=A�9�-��V'�MTq     �qԌr�?�(���Vn�ݝ�n�_�U�6�]��D���m����t>�%'ϖ�7W�(�nW!�M/�E�K�������[�w�U��Su�e�����5+N�=�����ч����.Ս�     �E�Gp��\�>��OY�'��Op���z�V�?��\��3T�w��<�>���ϓ{�Y#��ܮX�/����i�kWl     �`6�+'�J��<�ޮ'�s��_�䑊��ѿxx��j�6�<ד��)��uY�Z�w�j�%�M�Ks{ ���=�n���Wr�WV�2灿���`�w�i�Ƴ�l�/�0Sn��     �e�8']u昙y��:	���qE6�Xb����.q�k���L.�Ǫ�C?��?��V|^GU�F9�<��z=Y6�->�O!�(     �֙K&��BWZ�ō��\��g
��k��{�|��f�<������(�_��&��}����8o��.H�K �g��~ɍ_=�i��|�����?�u��Z������1���[dgm�      �8j�[�/.�Q�ˑw?m0F��d2��).���fcT���,��71�:jz�
Ba�6�,���>j      �8�f��1S��o}\��f�IG��Uۿ{�Cǜ�`ҫ�.�)���V��������f�A�_>-���n��?U|���Cr�+>����-\8�xR:�W/���g�M�.     @�F����Q+dp�x
cT�'��^���魆��9��{L���:F	�     -�Z:Ir�����}�����/�����=���W�����^�r��{�FcZ�����/}$Ս�����p���o�m�;�����h�}���
�;���t���r_��5,|    �J���3s�C R�5K��"Пi�X%�p8*#YY�Ur�i)��!�>�+��CT���ig���e��@���1
     ��Vo?{ٔ������n�:��k���L-���3k��3��t�o6uVq��S��*�Nʭ9rr���iln�ްL��[����p��:b�c6���FeP�}���co     Ⱦ�	Q�U��,�^��4e$�>�1�WV�A&���J��d�G���c5����j:d$�6�1�W���ʷ�      �)ǉ''-��c��`ϝ7^��Y�f^���(�^W9{|Aq:�?y�X���7ICk��Hup_2�L����w0��l�}�O�:k�@S?����s��?~v������	s�����$��}     �ktA�&:1t����H��)LߥT1t�k�H��)`����B���:�o��(w     0T�W�� �[�?��O�B��G֮O����U�� ߭�e����x���ߛ%�tp?{Y�~X^�p�k7}����E۶_�Z��iS�rs��[����#&���(      ���-�*ϳ�>.�=�Q}+��C2�Q}+g�2Fu��Q     ��e3FIY�3-}7��#�ZO�ŭ_[��{�S�^�h�7����%��O/~$�`X�I7�1�.�3�(-}�k��>�ٶR�6��w=v��f�Q��OY8^~��&	E�     ���C�Mϊ�|
�<zV�e��\�W7�&Y��7�(     ���'���W���W��K�6߽茫'<���3��jݷ7�*G�(���g�[��Y���(Cz�~es��~���5�����O�=��7��^v��}�lr��rya�     ��j��vh����x��nM�$�0��7;���Q�c�    ��*�ˑy�S�zkUS��iW	�n�u�N)���b6i���E�	���&��8lZ�޼���{��N��w�=�roe�7G�S�#�    @���<�T=#�<ƨ�1F�1�s�g|Dlf^G�,��Q     0D+Mc*R�yo[�y7V"�������?�����9z��}ϝP$c�ܲ��E�E�%SKc%��F�]�	2�o�f����.���hJ���R��     �y&����H�h$��g|HF�<�6�ǨQ�뛌#�9�;3�!     `�\�	��S�����n�t�_�}�o����*w*w?g����&�]ܗ���~7l���K�m�\���wA�ǡ��R�ԏ�9J�              @�f�-�b�C�~C�����r� �~���5����玝5�D��>n��p�YLr��Ҵ��aU㵂�����ۧ�ᯏ�8o�Z��>v6w              ��:vVz
R��i�֛.?�eA�U5/j��r�̚^�ot�K&����U��Y�/>�TV�M;�ko�l�YѼ/piC�M�ˮ�e�O��R��               ��`9zf���F�Q����JAV��������o/;k�QZ�}�2^Fn�}JIZ��pO�����zUc��<s��1�iٯQy�=\3g�               �K�R�qh���u�n���
�foSۗ���Gv���E���_�$�p_���{e}k����K�U����E"����q'�              0 �KOA�O�#Ȫ�/[�u��޶`R�-��\�+n�Ե�%Ӳp�X�b���ټ��?����kk������WP�e�'��Ѡ^�B               Џ��4�S���1��n羦{L*�E�>��B���BQ���M,Ҽ�H4*��?����5��-�t;,�O�|T�(               H�b6ʌ�����yW���\zrP�u��c~^�⿩�m7i���	E#/�>sl��}~�����+׼.�����큫=9V����W@�              ��F��B�Z�����.�s���������勵�w�X�?��,ܵ�Ko�izB�W�m�ؿ>Z<�d����W(����                �t��Q����5dvu����se���}�*pI��&��IY�y�Mk��mw	t����e�m�=K�              Nf�!s����}����x����H�Ӧi��c
��͕�IY�O.�ռϪ�����8�M����wF�ѫ��f}���:m�Ԗ�O�               '�˴���k�xJ�+������?�x���N.󎜀��R��}�i�X�;7_�f��^�)t۵�w|�G�o�               ��[�؛�i��pD�C�	t�������@�>'�x$ӲpO�_v_��]�YۺyL�{��}N*%�              �������������^]#Н����y�]�����Z�}t�K�>�Z��
t����we�i�}L�[               �X:�{�[��ҍW�\���7�I�>�\b6%�H�d-�^���Ls{ r�Uk7	t��C�Uv�j�gi�S               �Xin��}���o	t���W_�qi՟� R�uHe}�dJV�n�E�6m����"Э͵/�a�Z4�@HZ^t              e��nD_�V}k�ne�Y�]��>��騼]���+ЭG*��t�+��6��TǑ� �
               z(�uh�_4����u�j��(��Z�Y��٢�Y	��95�8��l�ZCk�nt��k՟�l��Y�:B              ���]vM��k�n�ֹ���F�Tv�ײ�|���?Y	��s�������ZS{�Ne�Y�]�ɱp              H��qfw_��I�k�`�?Z��qh���KV��4TpB�t�#ޫu��U��               ��qٵ&����]�RݱQ�>=9# ��[4�3,F.w�s�`�Q�>3��              ���i����m��p�]�k�T�����bҬO�H��n��	��k��D���b6
               ��������6��u��ŤY�֖��w_�p75�8��oW	t-kp���              �dNC�2
�
t��=9V��٤}���Ǔ,���!u��]�uZ����              0�Y����Qi�^{ Rv���d� uV�&�+�G�Qy��"�@ע�日03��              ������e8,݋D�a-�3G@�=�hڟ�`���ϭ�zU�@��&s��}B���              B!m�*�����dԬz�*�~,�%+�t�%;��ReG�]��F)к�P8*               �.�����l�t�n5���/0��4|"�d6��-�2�!�3�              0�� ��h���0�u�=
K&e%���4�S�6t�l2�jݧ?��X              �ґ׵��N��٭&����:2���J����C�>QC�@�,�W�>�1�               �����C5��Y�6�)G�kW���|�Q�﹪�= ����{�/�y�v�q�@לV�x����              �p��H�ۮY^�%O�k��2��l	�tT�v;m3��粕iݧ��              ���B�Z܋s�Tp�9�ըy�}DTp���׼O��:N�k��G���:b��               @o��>�P�]|3�f6\��?Ϲ�k���f��u��8ʤ�ܫ�%���`Ь���P�[�����<�ͤe�{�               ��#k��1-Wv�u*7�6I�>�6�K&e%�
Gd_�_����T��W�[g�X�<$�S�w�A�4�2��              0��#k�[�V��V�u��.J�����J��jp�ZL���,���	tǛc[�u���Tp              H�*Y�����N��wO�G��Z������ɤ�ܷ�m���5�3/��y!�K�^�QZ����I               �X:���=��
_d��4�s{M�D��Q��W7k�gi~���TTD���)׺�O�j?�               {�Z�#-C�E^��{w<|ԏ�X��@W�<��Z�������Z�=�Ie��V�o��"�@7"eO��vL4j�g(��ʋ.               �D;+pO��i��N痔w�]���u��(jޟ�ܫ�$��Ԙ���tX͆����*��#Ѝ|��\���T�aQC�               Hnke����\�r��|�g��+v{��W?�����?�O����)�ؾ,�uel��8��ܰ}�               �ow��i�Oд�)��q�z�Sqթ�/�
,߱����E��=�iY��6��<�>cL��u��˗�YWq�GN*��j��Ɲ�              ��}��N�>������r�_][�>O�>7ﮗP8"��Հ�;�e����Y�q�M����rx� �
\����`�              �SY�&u-~)p�5�w|��!��<vش1y�Z��1�HEV��|R-���Q���肜˅��.6:����V�{�              @����FN�7V�>���+S�����H�U��Gf�Q�~���F�!��_P6望�c4�W�o�7���}�\�|g��z��<�U�~��Z-               H�Ukp����q�nR?'Ȫ)e��h�g{GH6���UjXY뀻�j6���V9\+Ț	�����7�              �L��F�"F����_��슇��T���⷏^<���Ժ�w?��P8"ِ����[�ʅ��м��
WW��⊵�����7��8wb�8��m�e�v
�              ����U�=Nۢ�%�9����?yD�jAV�_xK:�}uK�dK��W5���[�ִ�B���r��F9�P�qFy�04����ō�Y�4              �p���4��f�/���"�͊
����??mt^����"Qyi���^ظG�?n���ΟXt��~�̥����A�\�cK�M(������`�               ``^�X)W��'F���-t;֏}���5mT��i(H����X��l�E�}݆�i	���X�xj�^*Ș�ŞߙMF��mjȻ��               ���/�?�����5�{���oV�[wS���!AF�p��g��_�����!��up�^�,�w���1����tZ��߻㉛tř�i��;�`��������ww�.y               ����;;�p_�u~�Ύ���iWQ5����4Too���H6�"���[��p�uڌ�s�R�Ҫb�:������aQ=��v     �
t.�8@8V !=�S� cT�ᨘ��Q�
�G�U_B��QcT���      ŋ�*���êy�GN/�B�=��Rq��i���{+�MG��zo�t��0����Z���Sf��nѼ�#��λ���ι���	�ƹ����u���v�Ɏ�f     ٣��p��L�M�|Bo�@X\v�@���s�E7S����0*N��z���a     �����;e���5����z�T��滿}t�i������ �nf�}����i��Q+�/�R|Oźu�X�<$�ܵ���e�K?����     �����l�S{�2���t���pl��::���U?���A!��B     @O�񩜹tR,_��������'��KV�+H��Ş��KZ&�6��'[+%�tpW����e�Ii�����{�]�(�'	4UQ5N���:��7��oC���q�     ��m
�7���^�4e��i
��B�/�
m�4Q�V��y�_�ڨi�uT}�/t�j�q�     @���ʫ[�d��r��VC�GM/��;�z�o?���M������������>=��eucg���٣���1�F�������w/:���ɛ���f�]��������%�    @�U�er�]�O{�U)cT&	tjoC��t{�1:w�@�*2�U�d�h�@�*y�     y䥏�pW��X��E9+��w~���������zԲ��U^�R%z�����?�cg��t<��B�N+����}��7u퇂!���ǿ|����꿱�C���v     ���N����k�̝�P��Nƨ�c����<z���9     ��;�)[��W����L(s�����o~a�y�!���~���ʟ���ғnW���%�GAj�ܷV6ʋ���13G���|��4g|ɋ�֕W,_��p���w?4i��Qw��ƴ=Ɵ^�P���      }ؼ�'Ч���Ե2ݵicT���^M0s�.�@���ò��p�&��u��5��Z     �����&�ŗ�N[���u�w?�č��|D0$Kf�Z7���IW����ʳ����]�]��o��f��*����1�EMV���J���ΙP�v�ב�1T�◧��&     @?��tH�?,N�I�/�;5����> ��V��lQ�hD�_���)(���R��EvG���P��4��{��l��.      ZZ��V���F�O*NK�V�I��S�'�o�U�ճ^�O���#��.I�c�����$�.�۫����w�	�Ƥ�1�L-����y��z�`@ήx�z�伍Sʼ�t>���� ��    �5����mrܬ��� ��Q���[���#���k�����Ey}y�1��׿��EN��+���    @:��_����%M5�%�e71��?߿���7_z�'����'+N^0�2C��A�m�Ͳ��]�'�����̮�N��/��If�{�%�$���Z�RPauW_�(�e�(AX\��R�f@B�&�!!!���3��{�eqeW�����|>��ɄDN����s���N��䷸w/n�!�{��]w׵g|��/o������޻ޒ��.r�g�    ����r�{b�V4��U6�����eq�?�|��w���9��2x͓���k�YK���������1�,7�   ��7�xx��]J=r`�nF�xƅ�����Olޖs��������-���e����X��7���MO,�/~dB��#���#������~�}�o钛�v�C�i����RR�:    �ۂ�ձzs]�`Cv*�S�J�o���+�9?�$H��Wʣ��)xͪ�s袵51vX� O�\u�H_�d]m,]_����܌6x   ZHk,��mh��5�L�t��I���Vuo�+n=�#���}��M���_�/Nd���i�w�a�z��9�������^s����/����]�w}h�!�=������U1���,   �k��#�xnk|��!A��6c?0{{�FSgl�'"�����o4�٭qƉÂ��E��������k�7�������3
   ��l)���_��-z�	;�ܥ�ˊ��v�^�������W��gԕ�J�[tu{]CS\vϜHQҁ{���h�q��ע�.,(�c��K�o�gط��c�7�t��5ŏ�=d�Н[�\���{^
    mO/����C�m�Yۢ��1x�9˫l�NĴ������ы�*c���u��m��e���!x��+�w�-m��9e���k=   в����x��#b��-z��#��+-.\��7�'�⛧��༫�������'݊Zn���{x^��Z)J:pϼ�dc<0ky|���m��t��g��WN���5���t����9����ߥ��v0�5�w�}s�W   iklj�k������l�h�;f����\���s>3*
Zt�	o���)&O��o��0�~xC���Q-���7WY��<eF��lF����Y'�4�mh{Uc���   Z^��ϯ��|��_}���JK���b�%�}��'?���.�����-�niK�m�[�/�T%�g.�oN8fp���>t��}_Z�q��_r�a�q��,�N�Ko;�	C��ثU�\�zuC�3si    �C�!�مq��=�����6EM}S�-]_��߯e������ͱ��.��gɺ�xtnY|h��A۸�����&^Y]����&�
��Ol��Z��   @�X�jk>z>刱-~�A}J�>v�n^y��~��/�N����~Ȅ�6n�?ti�m�M��۞����HU��˪�����?x��_�>�>|@�Ž������z�U�	���ר/�V�*{Y*j��S^�o�   ڏ����=�[�]�����s�*�7wӓ�c܈��yP��u���2��=xs�?�17��cx��u�X\�.��]���=,7���ַ�gT����   К�~��8`��3�����Q\p�!�]8t���}jޚC���Ś�d���;������&�k���l�����=���q�S�Ƨ�*�ػ����w������m���M�ԥS�ǘ��)}��(},�dߚ����Y�a[U    �KeMS\z�8�Sãk�V�N��k�G7o���9.�g}��QQRlF[˦���Z�������O?=*���ֲ~{}\u���ew
��=���E�f����RW=hF  ��W��?��\\��E���-~�lcy֬�[�v�eS?����0+:����sď{���/-���-�Ե��=����޻�=F�k��u-��g����=��'����sN?����ιjʷ�}�����l�uVw�X��Y   @��pMu����q��C����m�h���Xu��+�/�cM|��Q�B�WQ�ܶ&�#o��Mٌ���8��B���:�<:eMTՙѷk�������;��vB��V�LY���    �-��X���R��	���9���wh�3{]{��Uˎ�ZG^L}�巎�uP�;&�2�K+~����6~>yF4�����U��]r�����}8�����Z'��?p�}9����W~�3?ѡVf��?o�g���M9`��ݺ����Wn�=	�   �}{fAE�*���� �{*�j��o[���wf����F�o=D�ق�k��?���_T�;3wEU\���8��!aD[NenF9%7�[�wf֒ʸ����Z߂^�Hhul*3�   @ۺ���1nD�8�]Z휽J�
�>p��,6픳.���=퓷F2iRsA�.w_vĄ�_��[[�܍M�񳛟�Me5����=�q{u���/��U��/,(��a���U���z��t����w��+)�����Tڭ��+���6~zӳ�   �����GUMS|��C��Uߒ�6no�����[����3+��ා%���m{Uc\x��X��6xw��R��M����B3��e[��{]�ь�[��-�=�6���RdFw�����gwu    H�o�����=F�k��޷��C��2�O���pS���v��h�~|����?f�e�ٹg[�������e���hw�{f֒��܃����m�s�SRt�������i��«��׿��[N9�1ڑ�\O�L��3�������7��o,�   ����̲��8��!ѫ�k�c�_U��{]> �ɶd��ϫ�[�����ۣIZ��6~}׺ذ�����W+s3�&N?vH�iFw�W��įsϣ����\\��ڌ��aFw��k^{��R�   HG���ᙸ��#c`��z��n��O~����w���+�U~�?�8e^�3�]s��F�y�����ui�[#�?kE�:}q�'����)ϼ����O6�Mο��>���۫7W�:�ڻ�0o��o];�I��?�������}G���=���'�����B�]�9   ��g�����+�G��#K�w��9b�-q��[�_�cd��nX_���8pt������{h�����M��hHw�,t��������W3�^d3z߬mqӴ��hFw����s��+��G��w.޽lF�z~[�2}s�6�    ����i�}0ztk�츴[a���Ě�/�1���K�V}��o��|$������C��d��i�?�����_�������C�����ٟaĀ��s�W3�K����u���=��O���4���`��SG��y��;�{ri�{��������v�   �Md�G~��8b|�����ޥ���SK���5�l�%�j����1.�cm�[����^����6�fk}\���l+>;^yuc\t�k3��#�����|cm\�Ȧ��x�]Eοm�k3��A�8�.,]���G7��I�O   �e��ܛ���}�(,h��{qa:~���m�����^�������M:픊H�/������~:vdߏ�4�W�o����~|������M�~����9Ν<#~�����1����2�OI���<<���V�xmٽ��T�{޷?�R[�y~r��c�.>s�Q�6���H��O.�   @Ǘm$}r^y���2>��8j�>ѣ������T�?�%f,��iY�r�9oeU|d�>q́}�o�v��i�X��>�xnkL�_n�p+�ft����h�9����`�mX��.?��s3jD[^6��������7�޿O�*1�oe���Z�^�   h?f,Z�:3~p��(h�U�E�]c�]��?(�����[��zK�%s��^wˤS�Z���o��>jpi���:��?��`A�6�C��zsE|��iQY��Q������)~|������20R���>=s�ɹ/O�ȴ�K7�-ް��ʆ���=�S�Z��U��u�?�������c��>3��%q��s   �\*k�⶧�Ľ�o�����������J"����PW�3_��'�ŜUb�VV�������x`��8t����b��R3�W�cֲ��.Z�ͪh�u��7ŝ�m��gm�����#���q#<��������,��<ں�k�b�[���f�W~F��݌���܌f�M�����(   �>=���(*,�3N: R�{����}r_^yL}������[*��\^{c�u'�8iR����;O�߯w�{�7�σG�ӿ�kA�dcYu|��i�����90��ݨ�o̯�?�s��^;���SR�;�������#{�vsYu��+r���U���64>��[ɲ+�v����wү���)�ۣ���K���YR<�_��Q����M1h�kw�\��5;   �Ϋ��9zi{�ػ(�ک$�U����Fׂ�#��d�j�ax�ژ��*��9�g��,�}b^y��ۣk�siL��蘡�bH���ڵ��hb�ݚ�hM�[Q/���_�B���^�[�?���{e3:�4F�ftp��(L�3��]��f��U�9��3�m-�`��9e�����{���k}I�64{��\3�}/�����h6����    �w���<����	m8�^Ե˸���玣s?=��z�u{�����k˫�U��=__W0��8��OX�f��I����yt��.{�ҳ{�޽K�wЫd�~����Tm�^g^�d��Z�Y�Q�;QYS߻nZ��_�F�e�zv��s?͎CrǗ_��Sg��u�͵��Uu���CqQ��®��
���U'�N_����m$   �_l*����fGY��Y�6�OQ�v�%�Qڭcp���E�5�QV��+��� ;�m���M�ّ�.�ػ0z�׌��f�}�]�7eٳ�*w�U5�g��yi�R�O�\�?2ٌf���1g�17�5u���^�[��h겿��_.���>��{t/��E�;��g4{��^ݘ��   �4����O��/�URT�kD�~�/�cB�8��_�̜9QQS�\S��T���P���Xڭ����k�nE݋��~��ެ�\g^3-�ok�q{�������OǏO����MvEG���E�u�{�=2?��;    �LCSĚ�����R������z3J��]�y��e��ٝ!    ���"j���:(����zv/�;�U��c��/��];-6��DGС�L]}c�}�3�c������Ô���b�*          :��箊�۫���}J���1k��8��������U����v���5;�l����wtI��TU�򳛟���          Ӽ�[����_|��9�gк".��|4d�t�!������X��<~x�?D������T�nz&��/          :�l!��^�X���1q쐠�565���7?�0:��g�-�_������c�������5q��3;�-          xseUu�?L�:b�������.]���=���ٟfĬW7DG���̆mU��?��o{�.��UW�W=07�<�j4w�;          �6di�Q|ن���'�>�������q��g�����:E����o��o!��[g�t@���=x�o(��n���n          :�g��/���8��!{޻����W⏏�M�`u�	�_7c�8�w��7��/��0<xws�[�/������          �m��q��O��w��|l��ѽ(xw��My!����E��3�Z��o|&7,����Š�%�ۗmk���Y�          �O٢�;f,����������sD����7����-������:e����_Ys�m��9.N<tLt	��������yqg�ɦ�=P          x���?���8|��8��cx���{l���9�~[UtF�:p�T���e�Ή��[���ǰ�����g������          �D��}Ƣu��C��?`��ѽ(x�Ek�ťwώ9�7Gg���׭�T?���1aT���G���w�]Sss<�����cU��          �V}CS���¸{��ġ�㓇����X7=� zqE45G�'p���g\�d>p����~�0t�6�?�Ҫ������          v��꺸��1��%������k�v�|Y�eq��⑗V�S��7	oӬ%�ǘa}�S���#��]�#��m��^X�L_�U          ��m��q��s��̏��%N>lL�[�����Y�6t�����-,^�-οuf\u����~;űw���{DG�pͶ�kƒxtΪ|�          �%�Wo{jq�����o��q��]�	ãkZN]QS��]S�y5^]�=���o�������-�=pŇ����*)��h���|��Ћ+b���          �����«�Ǡ>%����kD��7ڣ��Ƙ�h}<��ʘ��ڨoh
ޚ��jjn���?����w�s��-Y�=� �6oM��j�[          ���۫���䏑z����>4&�4 R^�^^]�/�O��6���vz���{����,X�?2�����20��=x���֦�5[*c����Ҳ��ܢ����&          �=Y���/�{���8`���w�A���b�!���K��Y�>喘�bs�\�>������D�-�P�?n��8���j�=F��݆��Y �[�s���[+�յ�b���X��,��[��          t��������#ӣ[a�5 ����C{�N{EQa�?����|��tCY�ǅ����]A��%poA��"�����g�E]ch��گG�S���޻�(z�v�n�_ˮ*���®�����M�M��u��+<ʪjc{U]l����۫c���TV���         �3��m������e��*���JcH���׳[�)��K��WIq��-.,���.�=�uu]�k�����khʷ�Y�����WǺ���~[U��iy�VVW�+6��          `�jn���옻|sо�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          HBᆩgw	    h'.���v����HPCCC����ۃN/7�����"=��8㌱A�w�E}?��/"=r3:.��rϣ�rϣgGb���g�y�    h16�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��۵c   �A����Q-�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,,�ъ\�    IEND�B`�PK
     �]�[����C   C   /   images/ba153158-cccd-4fb1-9320-38bebad1b7f9.png�PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK
     �]�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     �]�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     �]�[���4�|  �|                   cirkitFile.jsonPK 
     �]�[                        �|  jsons/PK 
     �]�[	���Z  Z               "}  jsons/user_defined.jsonPK 
     �]�[                        ��  images/PK 
     �]�[P��/ǽ  ǽ  /             ֕  images/0b351edc-7875-4477-b820-546ce15be531.pngPK 
     �]�[$7h�!  �!  /             �S images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.pngPK 
     �]�[��n GV GV /             (v images/5a738b76-89aa-4728-b8e5-f09c859dbb14.pngPK 
     �]�[����C   C   /             �� images/ba153158-cccd-4fb1-9320-38bebad1b7f9.pngPK 
     �]�[�c��f  �f  /             L� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     �]�[��EM  M  /             zT	 images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK    
 
   h	   