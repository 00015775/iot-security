PK
     @^�[�<��s  �s     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0":["pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_4","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_2"],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0":["pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_5","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_0"],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_1":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_1":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_2":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_2":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_3":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_3":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_4":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_4":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_5":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_5":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_6":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_6":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_7":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_7":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_8":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_8":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_9":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_9":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_10":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_10":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_11":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_11":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_12":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_12":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_13":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_13":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_14":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_14":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_15":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_15":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_16":[],"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_16":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_0":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_1":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_2":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_3":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_4":["pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0"],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_5":["pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0"],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_6":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_7":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_8":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_9":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_10":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_11":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_12":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_13":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_14":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_15":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_16":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_17":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_18":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_19":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_20":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_21":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_22":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_23":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_24":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_25":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_26":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_27":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_28":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_29":["pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_1"],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_30":[],"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_31":[],"pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_0":["pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0"],"pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_1":["pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_29"],"pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_2":["pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0"]},"pin_to_color":{"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0":"#ff2600","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_1":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_1":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_2":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_2":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_3":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_3":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_4":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_4":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_5":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_5":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_6":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_6":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_7":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_7":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_8":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_8":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_9":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_9":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_10":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_10":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_11":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_11":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_12":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_12":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_13":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_13":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_14":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_14":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_15":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_15":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_16":"#000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_16":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_0":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_1":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_2":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_3":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_4":"#ff2600","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_5":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_6":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_7":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_8":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_9":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_10":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_11":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_12":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_13":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_14":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_15":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_16":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_17":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_18":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_19":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_20":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_21":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_22":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_23":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_24":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_25":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_26":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_27":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_28":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_29":"#00c7fc","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_30":"#000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_31":"#000000","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_0":"#000000","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_1":"#00c7fc","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_2":"#ff2600"},"pin_to_state":{"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_1":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_1":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_2":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_2":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_3":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_3":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_4":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_4":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_5":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_5":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_6":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_6":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_7":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_7":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_8":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_8":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_9":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_9":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_10":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_10":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_11":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_11":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_12":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_12":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_13":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_13":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_14":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_14":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_15":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_15":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_16":"neutral","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_16":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_0":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_1":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_2":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_3":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_4":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_5":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_6":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_7":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_8":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_9":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_10":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_11":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_12":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_13":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_14":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_15":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_16":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_17":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_18":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_19":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_20":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_21":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_22":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_23":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_24":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_25":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_26":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_27":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_28":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_29":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_30":"neutral","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_31":"neutral","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_0":"neutral","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_1":"neutral","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_2":"neutral"},"next_color_idx":3,"wires_placed_in_order":[["pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_4","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0"],["pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_5","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0"],["pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_2"],["pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_0"],["pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_29","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_1"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_4","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0"]]],[[],[["pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_5","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0"]]],[[],[["pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_2"]]],[[],[["pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_0"]]],[[],[["pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_29","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_1"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0":"0000000000000000","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0":"0000000000000001","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_1":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_1":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_2":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_2":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_3":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_3":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_4":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_4":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_5":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_5":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_6":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_6":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_7":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_7":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_8":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_8":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_9":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_9":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_10":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_10":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_11":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_11":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_12":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_12":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_13":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_13":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_14":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_14":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_15":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_15":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_16":"_","pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_16":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_0":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_1":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_2":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_3":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_4":"0000000000000000","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_5":"0000000000000001","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_6":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_7":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_8":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_9":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_10":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_11":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_12":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_13":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_14":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_15":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_16":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_17":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_18":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_19":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_20":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_21":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_22":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_23":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_24":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_25":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_26":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_27":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_28":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_29":"0000000000000002","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_30":"_","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_31":"_","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_0":"0000000000000001","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_1":"0000000000000002","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_2":"0000000000000000"},"component_id_to_pins":{"c761db77-2aeb-4e5e-894d-70927fb06784":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"553cb021-004e-41a4-a0f3-1f1baccab3bd":["0","1","2"],"a898b99c-4f03-4cb3-8c38-65f83c4f7bf7":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_4","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_2"],"0000000000000001":["pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0","pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_5","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_0"],"0000000000000002":["pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_29","pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_1"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2"},"all_breadboard_info_list":["ef713389-553f-4ef3-8c4e-ae27e235a732_17_2_False_925_355_up"],"breadboard_info_list":["ef713389-553f-4ef3-8c4e-ae27e235a732_17_2_False_925_355_up"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[1356.25,492.5],"typeId":"b269da49-8c00-4ebb-bd25-5859ea0c7cad","componentVersion":9,"instanceId":"c761db77-2aeb-4e5e-894d-70927fb06784","orientation":"up","circleData":[[1337.5,635],[1352.5,635],[1367.5,635],[1382.5,635],[1397.5,635],[1412.5,635],[1427.5,635],[1442.5,635],[1472.5,635],[1487.5,635],[1502.5,635],[1517.5,635],[1532.5,635],[1547.5,635],[1283.5,350],[1298.5,350],[1313.5,350],[1328.5,350],[1343.5,350],[1358.5,350],[1373.5,350],[1388.5,350],[1403.5,350],[1418.5,350],[1442.5,350],[1457.5,350],[1472.5,350],[1487.5,350],[1502.5,350],[1517.5,350],[1532.5,350],[1547.5,350]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"2d7cb472-066f-4306-872f-cdecc946e2eb\",\"explorerHtmlId\":\"e9503054-5667-4f99-acda-29509149cbf7\",\"nameHtmlId\":\"19e4d613-6efd-4ec8-b7a7-175ff44b25e0\",\"nameInputHtmlId\":\"af3a1ee4-803b-4e1c-b5a2-9cc0bb627783\",\"explorerChildHtmlId\":\"dd622af1-c564-4f2e-a208-41fd449ed125\",\"explorerCarrotOpenHtmlId\":\"13943eee-45fa-43b6-b8f6-87055934fb31\",\"explorerCarrotClosedHtmlId\":\"168d702d-1f99-4614-b60f-2cd9cd669ee4\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"01e2bb24-6c23-4f1f-b771-37a4581ec2f4\",\"explorerHtmlId\":\"a163593a-c2f6-4caf-9dbf-13eab7bd9be5\",\"nameHtmlId\":\"a97429d9-5346-4bb8-8df7-1c2c8e7d79e4\",\"nameInputHtmlId\":\"e4bbd91e-593c-4741-907e-294e7b88c5f8\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"6af55ef5-d33c-4a42-a55e-ef5c39e01150\",\"explorerHtmlId\":\"4db22048-98d0-4063-aa20-e125885fa3b7\",\"nameHtmlId\":\"7aa756eb-39dc-4835-ae45-6650d452bd30\",\"nameInputHtmlId\":\"9ad5711d-e8a3-48e3-b3a6-223cc332ff6e\",\"code\":\"\"},0,","codeLabelPosition":[1356.25,335],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[965.9075245000001,132.50997799999996],"typeId":"38af4144-8c5a-4c1c-8860-ff9e0c7b1ede","componentVersion":1,"instanceId":"553cb021-004e-41a4-a0f3-1f1baccab3bd","orientation":"up","circleData":[[947.5,260],[965.4655,260],[985.951,260.24]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"DHT11 Temperature Sensor:\n  - VCC → 5V\n  - GND → GND\n  - DATA → Pin 2","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1251.0029296875,200],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"a898b99c-4f03-4cb3-8c38-65f83c4f7bf7","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-6.06147","left":"872.25000","width":"715.25000","height":"666.06147","x":"872.25000","y":"-6.06147"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0\",\"endPinId\":\"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_4\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0_0\",\"rawEndPinId\":\"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"887.5000000000_365.0000000000\\\",\\\"887.5000000000_357.5000000000\\\",\\\"842.5000000000_357.5000000000\\\",\\\"842.5000000000_665.0000000000\\\",\\\"1397.5000000000_665.0000000000\\\",\\\"1397.5000000000_635.0000000000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0\",\"endPinId\":\"pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ef713389-553f-4ef3-8c4e-ae27e235a732_0_0_1\",\"rawEndPinId\":\"pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.5000000000_365.0000000000\\\",\\\"902.5000000000_320.0000000000\\\",\\\"985.9510000000_320.0000000000\\\",\\\"985.9510000000_260.2400000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0\",\"endPinId\":\"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_5\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0_4\",\"rawEndPinId\":\"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1052.5000000000_365.0000000000\\\",\\\"1067.5000000000_365.0000000000\\\",\\\"1067.5000000000_320.0000000000\\\",\\\"1592.5000000000_320.0000000000\\\",\\\"1592.5000000000_665.0000000000\\\",\\\"1412.5000000000_665.0000000000\\\",\\\"1412.5000000000_635.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0\",\"endPinId\":\"pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ef713389-553f-4ef3-8c4e-ae27e235a732_1_0_3\",\"rawEndPinId\":\"pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1037.5000000000_365.0000000000\\\",\\\"1037.5000000000_327.5000000000\\\",\\\"947.5000000000_327.5000000000\\\",\\\"947.5000000000_260.0000000000\\\"]}\"}","{\"color\":\"#00c7fc\",\"startPinId\":\"pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_1\",\"endPinId\":\"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_29\",\"rawStartPinId\":\"pin-type-component_553cb021-004e-41a4-a0f3-1f1baccab3bd_1\",\"rawEndPinId\":\"pin-type-component_c761db77-2aeb-4e5e-894d-70927fb06784_29\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"965.4655000000_260.0000000000\\\",\\\"965.4655000000_290.0000000000\\\",\\\"1517.5000000000_290.0000000000\\\",\\\"1517.5000000000_350.0000000000\\\"]}\"}"],"projectDescription":""}PK
     @^�[               jsons/PK
     @^�[�.��  �     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino UNO","category":["User Defined"],"userDefined":true,"id":"b269da49-8c00-4ebb-bd25-5859ea0c7cad","subtypeDescription":"","subtypePic":"e30496d1-6e1c-40fa-a66f-2add70ecdc94.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"a7fde0f7-2836-4f0c-aad0-66dcccec46ff.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":9,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"DHT11 Sensor Module","category":["User Defined"],"id":"38af4144-8c5a-4c1c-8860-ff9e0c7b1ede","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1615224e-fb94-4bec-8b91-0567bb6a6470.png","iconPic":"c64d4bdb-8b24-4d1f-9af2-aab9cfab9f47.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"17.14286","pins":[{"uniquePinIdString":"0","positionMil":"210.61667,7.20952","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"330.38667,7.20952","isAnchorPin":false,"label":"Data"},{"uniquePinIdString":"2","positionMil":"466.95667,5.60952","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     @^�[               images/PK
     @^�[�R�W�  W�  /   images/e30496d1-6e1c-40fa-a66f-2add70ecdc94.png�PNG

   IHDR  u  v   ��:   	pHYs  �  ��+  �	IDATx��	�ם�����w�}!��l��Zhz��@?aK3�`l���-Ü1���vws�c�w������=��-,��lt��#��%K��� �ElE-Ԟ9�ݪ�����̈��ܾ�9A%��q#n�ȼ_��"!�fs]uD��$�\B�0$R+�B!��� &�t���4H�BQ�&�뿿6�m��#�B!$71��_�yd�䪰��s˚�u5��NC��-�B!���&��E��]S($7	!�B!$/�UaGQ� �7玕�%�7��t����˒i�(���F��C��B!�B��EaGQ��u[7a�����������!y�ђiF�����!�B!�&ׄE��l��emM��8If��?�J���2)K��̙3�ih�kB!�B�p䒰��s@u$��X^e�������r!�B!�&W�E�A� yD!�B!Ğ\vu`�KB!�B
�lvu)R���B!�B)H�Y�Q�R �b�4I(z4����±ȼP(6Mb���hB!���d������gL�ۧ���ή��^7n�DB}���'�;"��|���)*�Hqq��_����}�Cr%�$���';e��a6m�/J�l�V�,7D�Z�Kk�B!��Ad����������'��s/^��󘢢"Yq�d���������_:}2�D�\_(����uMN?۵u��.�-��-��77�B�w�B!��6aGQGH����6�>�-^���u��f�Κ"%�ֈ�,����3�z�����v�.��]�X���vٮ���@6	;�:B�XL��D�~w�>Ow�u]s��ڪG67�%�h|y9��1���2���ns����,��v�.�e�fڪG�G��)�R�zA��pϰ��S��]��o���ϧ��lvu��8t-}х�İqsi���u;+ݼ�(nr#�!�B�lvu��0qA��?A���B!d(�vu��(���˥�:+vU�ln�H�gB!�B�@�2�6E!9JT|��K�b�<�uk:�S����̮(U���]��v�n�+�Ѩ���z��P($�)��a�l���n.@QG�����S���������:P^^������%_n�leڞX�3S��F7��ܺa����tww�},��%2r���8d�l��]/���������%W�^M{_�pXƎ���e�l���n.@QG���z�����ܬD��Ç���9������v�T��0A*jj���Zjkk��#���m��l]�[�ym(~����EZZ�?&ҙ�ab6v�X�%����]��v����D"ERQQ�քTODQw5��(�e�l7�vs�� ����Ւ
��w�Tg��@̝?^.�=+'�~[�����bn�!�ʌ�!��%1��?�=��5^�?�W�1y�x]>n�T]3C��~���4IF��D^&�(��yw����\����Q$<�ǁ:v5�lݒNҔt&hzb�/xL��.�e�l��v�"�	�y"�v�.���l&�Άx�\B̝<|X>nj��C��Q#��j���s����i@��a)���R,��v� o��5)�6M�/�s�6w��3&���Hn�h(�(�C��Y����<1c�l��ݠ��
7R/&�l����t �Έ�n��s{�Jǁ�2�s��e�q�t:��]�q�`�.�H穓����rd�T��?�/2�����^�3���J$K�G���D��>Jy�Oz�'3��v�.����^�p!���k��Γ�(�e�l7?�O~�qŕ+W佷ޒ#��i55Rk��+��K�"�G�ʸ��"i;}J�ܺE.�志ًɄ	�8 &M�E �f�#[�xQ���=�'m^�M�]��v�n����J����a�l���uDA���.W^��\?�^�;&}==��qWq�ʱ�~"��2e�!�a�I/a�͐�#�B!$#P�%�~�{�D��'�*�����(~ �$Y_V&�엽O=%���i�K�h8�$Y�f���B!$cP�8����C`���ʩS��[Ɉ�"�|��4��?ɟ��*��B!����Y.�񆴿�[�PV*�t-�.��7������+�ň$��7��/a=K��B!�d��Y.O��_�5u�r���(nP®�Hξ���;�]'�.^���B!�BR���@���;;��Z���C�
���YR"o�h�L�9S&N�*Ğ�"��.ٕ3/�pB!���AQW����_K�'�'��Ύ����G�R��.����e��մ�B!��"uHgg�m�\S[#�?�P��;�,���W_�O�/�q�&	���e��θt�B!�d������Rc���u��Rˈ����K�2��P!Y(�B!$cP��?u�|~�ti��J���Q5���"= hj��UUr��i�&`�+�D�Hӯ������L��,P�n��J��3fL���W�]��v�n����K�������]��E�fu2��J���P���}\\/;O������ ӥ�v���r���y�g��4!�ڪG6/o�޺��E�^�g���r�5�8�L{{�tu%@�v�.�e�^���\.X���gp�8��v�nf��F(�
���pD:._�l�(Vֺ�R�% SB*+D�AC�;�Ĭ�������6�4��v�.��8��c�:�\ii���vB�v�.�M��l�����x��T��I˙3���6�غO��!��BrO��Ӻ��;���^����t��vb����g\�.�e�l�i�^�v"�q;!e�l���n6CQW`t��H��2^�`8"�R�t�!�)���$��uk6ׅB�-n?�DdĈiM�4�b��b)�5�]��vٮ�v�"�,�iND5zB��ő�]��~�� E]��z�Ttg���7l�E�p]tw&c�j��ӱ�Iww�\�xѓ����]��v�h�+P����]��v�����("��^�v`�#��pcţ�^��}A�1i\�5��#���Yа]��v�n������]��v�:BrXʊ��f�Bٺ�9�6Q� 5�$�B!YE]�Q\��<LK]J�BrSM$������+����M�B!�B�%7f����ha�����\1�r	!�BH�AQW`�"ER\^.�L�:MuN����z��7�>�5�Y)��fs�@R�1tg&�T�p,�u�|��X�j��t`�l��]?h�%o���n��׋�]����+0FL�,��[q�X_�d#�XLjg��X�B����[����ۿ��)���:t!%覊ϼxe�d��v�.��/�z�]����f#uF̈́	r�w���L����b�!���O��;(��q�JL���}�3�x;5/�D��pmb�B!��E]�1a�l��g�IyMMV�:�>c�<w���I���"y*��&	E�FCrԼ]8�g��i��p����B!$7�����m���Ei�L^�{��U��kJ++���LF������6 �:�1�~�mB�C	<cQ�톼9 �Ƙ2Kgϐ9F�׻���!�BH�������jI���U����<o�Mz����/۬u=��9g���ds&���|Ff:���[�çdE�.�ґ��M����>-�&��i#���xE���D_?(�9x>�BH!BQW�\w���jӯ�v�Ȭutݱ�|�s�B����R���2�<�z�{fLTbo�S�$W�3�g�ßW�BN8��M���E�e��?S�B!�E]+��[�T"}�Uֺ�hTb�2��[��lc��k	���n����D�]r�52��F�_j�\ �®�!;��h�{v�.P�,��}�8�K�I�/��Vgg�kt�⵪���l�

����%K�x]F�-��@�A��Jw���BH62e�k�@�-���z�{��qawǌ��#D,q�"��Ϥ�CއuNY�6|Y�ϽV���wBH*`+���&�1���
� ���P�6[�*ʔ�0�	��xcz�O^�J˳>�-/�����KnW}��e�p�X�q�k������~5h}���Xi��l|�ׁ=PjZ�����X~�l|��� ���E���1�����u_f�3����(�
X����"���[R9r��_t^��+����z捴����,%]W��Gwi�|0sQ��6��(ǧޜ��%�W��^�p4�z�N�M���G�NT�~�0yHֶ��m��#)�]z��������k�'��k=Ld1�����'�j�j�O���H��bw�R��8�lu)Ʊ�_^?ŗɽ�O ��O��BM|�=����^-00&������t�w='ZLڡ�����n1���O��y|��ϸ/���>�p6�86W&~��@���-R�~��v����𙄢����t�����d����~Uz:;?�]�4]W8"��o�F��:���v�o�-�zE��ًmw䅣�o*�n���������u���B�_k�>��>�)�ښɤг��W���	��ǰ�a��ɒ�Ƹ�$�1�!��ˣ���6_�E�_YA,�Řઉ��>�q�jf���)�t��z��p]О��Ax��%���7=̖;e�B�|?yٓv��8�����x�u�/�PlZ��|�=��z|zu��f��M7��3����7c	�m���~�}�o,)�
�������o�������Gv}}�J�����/}�+a���Rv^�����RЙ���Ϟ��o��ՙ�x��#i��%z�ݐ�A���uB[i�� �u�fr�uz��, �yjV'c�z�����gF	��L�1m0�_Y��0��x鎨,9F��1��A�d��m��7�S��w�����ǈ�hA����B���ĸW���Ό���z}���8?�+������1lN��7�74������񷖢������kk�7��]�0i�\9y*0a��^����ZXi�	;��N��!�4��������M�T� ����g_2<tC
�̮ts���~���νmZ}� k!���D�ڮ~�~0�����X�(7[���t�u7��>��
��ۆ��n�����z��A�,fk�c|`���S�l�����_��,�;�/�+�)T���3��H���.�ʊ�"��%6���#2j�t�w_T	���������ꀅ�S_]-��Y|I���&���];a秠ӄ� +�<*s�ޗ�����Dx�Y�nH���VgGܽ�C�:e�o��,c⌶!�!Lp]1��>�߫k�����/�ԡ-sL�H��7Zܩ{��)����DL�7������G�[Q�^N�16�����\@�v1Np~]/|��G�Xt�N�PI_�v���9�c:p�xy��ݍƘ�k��J������Qň��kE?$Ľ�,ۖ�E}}���7(��n�?l����q;e�\�xї�)���t�E�/���~#-t>ⷰ�X�]P횅]�����?��>$O	
L�Ryr�I�����ܐ *%f��ۧvGN���ަ�_b���ya�:L�0q�rB�bhD�.�ؿ)_Z2H8@X��DN]+�
�Mu �cU�K��Ճ��X�u��	�����"���@�^�D?\~=��y@ kwD�}���xy�hGd�wf/���OQ�Ǹ�A�-��a��Ȭ�V{�Pԑ8�c�Ȣ��[�����+R?m���?�I���tG���Iф�x�7T{��m2a�A[�~]�� ۅ��-*����t�vOO�1��(k�%p�n���S�$;h
�IM�&A��K�i�x=�18`��dj�O.Ov�Ƥ�j��Ѽy_&&���t	
s������o.��N��^�� ��NFa��^6m���!~��g��D��8�y����>��I��'�;�vPI��3u�Eb��X�ZN<(��~Jjjk�j�h��N��h,&��R���J����	�t��!�ۓ�v+�.*���%�,(7@��p���+AYhnHzb��?0Q�F�vu�3��`"�[��,�WɅI�~=Â3���A��*�@z�D����&���_�gɚl���������	���w��_���Dj��$�"ᆸ�2�X��D.��=��9����ɍ���#�D&k��5%Yjo�5�y:���2i��㔂�쎘�:k׻�y�,�B
�� �{��}�8i�Ln�YW+������w�?.��|"��쑳o�!��=RZ^.��s��q=Ʊ����װʕ�+�fϑk?�X��e�HD�r�t�K��8���}pD޾|�>���rdu1�KL�G�:����x=�/D7$�~aԓc�V��l��˥�BH栨�������'��/")ӢN���y��+r��u��Yi�l�7WTT$+n�,��1VUU%����y+��g���d�	��KW���.9�Ijc6�v��,���fx�r��nHΞk��v��Ep�q>p9��h��=�p�U�.�[
��5�t�h?\�
�)��_I6�1g�h��ٕV�F,����������,�q2����:�f��m�GTIEE�||�^�@е�uH4���Z�(�ힱo�V��mF��Ew.��+���Kn�O;�a-,R�<~�]�`�D9x��,���\�e0��ص�����$;�|��6m�<����E!��1#�K������ܦ���H�(l�;8وj�V��n������2�&d*�?��]3�^|CV�5O��x�lX|�<���B����`\��w�,���������8Yy�Lyp�̂'��oճ/I!pǌI�/Ɠ�u]�`b��{���d��7��|����g��9���A�B���ۭ�����B��v�]� qn�Ə���L��g��>,���55�"�&����Sn��+WL=N �
a���)#j��X¢Y������T�>&�:B!y���a�T�L��g�������d�xϝ_�B'�t��fA�?����X�w<�$���[��:B)0�����<����i͸��g��up3��E�aJ}���z��#��{���8)�����վ��½u��I�u���JQG!�NL���7('T�s;2����	q��!$�8p���\aÀU%(��q�J���B�/`��=a��{_�s��:x�s7Ld����e�=w%�,`��G(�)p.\h�ʲ�5��L-m���nSK̻vۤ�|p��)˥��5/�5똝�J�������������l7V��o�ض�m!�b� �N\nl�[h�P����Ҋ_n��]6{��8[���<NNCQGH��'����G"��_���M���;���.�]p>9�*�	^���t�ty�ݏ���L�k��-�J���khX���E'�@E���g�(�qR(�k�vi�O7�U?~I��_1��.��HP�ȏ��H~}�tt'/��S�ejU�oA��G_> �p�X�I�?u�W�[%�X,�p�k�����O����n_��n$q�ӧ���{떑�v�G�{��A`��(~nqY(q@�SP`]̚�GOv�"�]��B'�~���.���e�/���3��.5ur�r�ZR�����b!��F�3�BD���	����3����v���ue��'!��������/b�T�������?�ӌ��N��iWM�{l{u��B1���R��Iv�/\+\�c�z����B'H�s���Źٹ?��+�cϿ��1������E!�d *X�t����)�����+��%���.7�p�l�_s{:���맨���8b`�we�1a����@d {��	������+�qR(�q�K7$�5?)!g���B2�v}��!������z�WE��K��@�!^.YLl�v�|!���ڤ*��Z�nj�6N
�|���u�P�BH�����
��Ec�K&�����VAa�6��a�öX�0%=��b�L������m��84\�$�������)))�p
	C���3�t�d-���\O������:gwV�"R�9
���2�&��{�-�T*�L�}����M!$(겔�HD"���]6��P(�����z締C��;��a&���pE����e�C�Tbě�dm���fApB�'(겔ʲR)-��������d�7i�<�ٛ��B��%����H��!vo�O^��Y/����!�;��:��U&8��"��(겔_:#��?����.I6p��]	LB�� ~A�,�5����q1�R*���z�3o:p����!�!҈�JG!�E]����u��6N�td�Ő� �5K�u�u��%IQ ���	qg�m������r�j�Q��R��[f����p�BH!AQG!��#v�jAǯ�
��t�<:���Æ�d%(�|۷��MQG!y	E!�d��[�Mi;���f����B����T̘('.�����(��<}�qu�������8S�BH�$%��^OV�ض��
<��{��];0��Dۄ����	�
�W{��vU=X�4_C(��L���	�GL�d̮U��X̟A�nX��y�`���i?����X�q;G���m�,38�T���"�F݀�����	�VӇǅ�6��!I������ yPV3h/ȶ	!�I&��CVg�}b|�Y��`���w6�uy���0n(��^�}�qȓ�i�dJOO�yd���¯�L>q5�}@�$V7�T�h�D���"� x �3N�}Z��$Fy��W��{�V���>��3�Y��2�6!��Ȕ�B���0�x�6����7�E]� +/n2u��ȸ����y��3�Aԩ�}	�^B��%e�3X��%�����G��.�����j)��	!�E&�~Ga�H�/��bN���|����Ж8�Y��MR� _��B��{?f�a��o�b���e�B�V2%�0�ł��{(��S	����)E]�I�6��z�UΘt��͈xB�3�?>�u#�OB�q2)�0'���]�Q�Z��U���k���u�ʠw��x�+�a��l>�M��u��;'n<q���..O%o�I��m��t�
���po�>�}ń(�Br�L�+�0�p�[���y!��E]��ڌ��p9�D)�9�?�3��e����n�n"�=k�b&| ���a�����U�"D�'��KdR\��Ƃ��AY7����i<ɘ�曰���C��/1�a)�ൖH5�h�Qt�X���g��F'3�%�c��
��`���	!��
��+/1']Q�7m~71n���@5�uyN<5�W���v��TQ����e7�Nɞ�O?����,��?�_n���Cr�\3���`�Vp�<�wu�Br�D�J�՜��q��06����:Y>z�P�9�Ϊ��-���������TC��cIC��N�n�tC�NS�����RQ�����}���M��*��p�'��BH��J��-fڃ�A���aP�--� ����R��ytd�?I�!VzEƗ�%�� ƍ�B��%��q�<��a�k'֍�U�@�;�S#���?qi��K����B!$U2i1üT%�3�=j�nr��3D�.��C���������@Ow׵�����	M��e�� �7���x��͙(�%�����,���칋�օBl�B!�ȴ�L�+ю����_�f>CQ��p����8�$&l��R�
J�J�.a鸎��!�BH�i��99�O3�:B!�BI�LY�̞d�J�e����:B!�B��m1�xӮ�?|!���c�^�����ˢ��E!΅mRY>8�㔉����*�W;�.!�B��L��`�����.�X �X���7|r�U:;:$bI���t�ty�ݏ�Ӈ���.!�R(d�b�6��vj�Os��|�������V���J,I�͵ӧ��ߟd����P`2kEե|��!$����5y��bҌڱe	1>o�Bm�<,$�&��,�zbng���I�Sk���c���=o�6����Xp�Ȥh�}>�����.�4o���z���.C7��m�r��s��H&�Le�b��2������#u�(��|f�ZZ��b�*�0߸�v%2�Ց�b�f=i��b!`Y+��Q��DYqL9J$�ʛ�O7�%��˄�2&���p ��b� �͢"m`тQogm��^��˷I��K�%��1�'�wӇ�n����7�������|���%��#�B� z��Č1	Od1�d��:�HC.��v"
� �����Tn��T�G_����a����)���1���1�zhf�����?���
s&����Uj�J���y���e���&+n�)e�E�7����E�3�q*V\��������	�ځ���{+_k�Q�B!�dL��.�=n!�COJMԭ�hݢ�_eU���@(b_N\��W����O��2-�v�?�D��?&�X�Qh�� u�z[��,� ��D.�A1��Fv��Wj�J���Dyp�Ly��)ٶg��>xX�_9��0�^�tve�Z�)T<�3�J�~���4u��!ݥR~5�:,}E�i���^J��$��x���%v1fLL!d�D[��(ڃ0H���#�c׮�f7MXӴ�(�����f�mq܉b����	�K��`a,Y���Q����P,rpfLTKKg���"�'���[����a�S>�c����}���93u��!�\$��h���@��*��#3nS��l��irz�ra�t���I8�h���5��w!��;���范N�qfں�8>�
��]
{��X̠��&�ɹ��iˡ�J*17`�3[⬨�+Kn�[q��LZ��P;06��٧��x�}��1c���k�,1D�t+��%��|���� �"(1��.�]�:@QGH����Ł,:�t�Vǧެ^w�T��7�O�;s���%����٦��ٲ�J��d(��I��]0X�Rbb�Nh���c��N��ר~���cj���""�1b=D���t��\���:+����Ձ?��)�� �~��[ԙ�w�E!y���*�j�NX!�(�!~2�,��d�.�~�}C�4`1�;��D�, � �pf7Ns{U�`��=s�%�S�K$ˀ���x�G(��s�X����'��vt�?��PI>�qS5�P� MW��AŨmzz��x]:����tK�uG���巆�7�s��S���[�^o�$S�dsL�S ��A�	�f��k�N�J�'���o fk������X�%�WZVv�'��.\M�~e\HH0��rLN�� �V2A�W��+?�!�OT"c�9\9��0�5i��-�4��3����D�Xt&�t�� .�IڡV�׃�Cܟ!�e�4.�Y1���w0����O��P(T�F�4S���y���|�d9�`%��z]"�O+h#��p��7&���,%]W��2\"K��6���������^I[�9i�BR�L� K�X*�	� FH%4�ǯ�׫Zl)�K��&J��\faf=�qX��ݢ3]ډ�e邔�� Z��x"p�2Q|B*B�Jz�*��N�X��awp�_!�d���}��)oߐ��I��$n�ü���}�#!���y��Úf�P�tnu�$�W��֤,��;W����ʄE���U���#�B!���$�ʹ!Obֲ��$w��#�B!���S�}@��J�W&PV:S�ARP�B!��@�k��X]eIa@QG!�B!9E!�8S�kdʈ!�B
���˕<+|NQG!̜	�e��{���D!��B����t�sy%�&N�x5g� *++�kkk�������B�Pv<����BHA1{�(y���dճ/I�@K!y��o=�
�Z��Qd��^Z��>���Mdl���Z�A�2c���`��/�ׇC6�-/�5h�(���梴���~����ˊ�v�RG!������_�|����D/�2s��	�a�u��z��^�����,kafʹ�m��P��r�O^V�v>�y����a�;��\�k��/��lqw<��1u�B
��Br��-�-R��,� DX]E�_���[��.��D�U�A��3 �O%}2>A��! ��@`BB�xj0�ԢB!��&u�`py�����Ġ��9�BDc��uS��s��B!dx(�)0�K�x�2���->�YӇ�Ӳ�Ab��2g`L!�BHr(�)0`�j����3?|A�l�D)���0�IR�hft��Y4ڶw�l%�Rq�$�B)t(�!I��S�S�E�o�Pg�T�Ol����*�bF��g�C�X��~�B!��:B
X�҉UӂLe¼�:ٸ��x"s��d���@�S%`I��G!�R�P�R`��HY��F�(��jZ}�e��.90h_�|��S�_?eP�:��B�]:�!�B)4(�)0��R�N.�o+�t;����z;�N|�*n@�ڃ��N8B!��ᡨ#��� C]8U����+�,n��A�i�I��-v(m��%�A ��9�PG)4��ר��S���s�$�r���B�N_����`��3g�hc�^O�33�c}����#B��#� �{�W�����!�l����ֺ��z8��O	D�Y*!!վL�a>N����<�d��k�h�3q�Ԕ�������!^�>)�Q�/_�p�}t��LQ��3dh?�tv��9tR	�|�#'<~�]��;��x��WdǛ��n�^6��g��;{ze���&?}�C5>w<�L�9��cϿ��ͺ~E�.��a�-3e���������^���������}j=xl������o�_o>�m��-���F�c�1c���gʉ˭������w4,S�֯xj�:v<8�~�g��Ot����r����\x���#��?,�[�z�\	�Br��U|o�z��l����<g��=i�Ng�L�T�[���v@,&+o@��S�Je������N�Pq��G$
��FGw�t��Ji�a	�'C}�=r{�a�W0y\}�<C��H*✀I*L�1��}�<cLn!dr�eF-��O���ƾ��0�Gm3DF>Z�0� v�k�!| � �c�!n��t���H��:-r ���t�s�{����o2����Ȃ�t�Ѷy=��zX�1V���m�1b�pXf��m+�c����C��1O��Ա����|�����_���*��G�|y���~*�qS��'�U�Ͼ�\m�q\xb|��1��u�B$��%]���nҵ3��"��$e*�$�ʙ��Jg�Y˛!�7�V���]��"���y�1!���K�k�&�Xc۞�s��R�������P�-ܬ�Z��*�cb�R�Q.�X �*֐��N�=�}�;�v�Nm{��59����q�և���hA��7���v�6g��ScWO��2�;�B�_�	(�!����vJ����HQ��yդ�k�L�6|�6�EJ"���o�~��l߳O�� Ŝ�'�R}ѝ+،vc���a�^�"j�,f�����x `;/�{DY~a	6�_�,^*\�l�X��} C�����"iuK��cv���p�4o�s�;���h4$�.�wʫ��&;|�YY���ߕu~@�O�;)!~BQG!9�.9�.`2z�;����j���>c镪�	R\Z+d(�
�Z�e.0	�t�]j�Mna��f� ��{,G\�0δ��������"��e�qiE�~�&�W�yQ}�f�8�M�|#�^�m����/�c��Y�#�N?X���B뵘�k� sL��c��b�������a�1AP�عUϾ�����S��Y��[�����/�ԭ|z��{�<���xL�'�W��?|AV�2k��D�b����;��*L��:B!�Ģ}���+�XL�Q'a�3�>4&5Q5�)�-䏮o^ły�v���L%w���+Y����d�!H��}���97O3D`œ��k��XQ	D��Ԑ�Xv�!T��J��uvV+�cL�^%bf������sJ�����������X�;(���ڕ�����(��P�B����Dj믑�1I)..��2���弜9sH����ȱ3%�H��bN"��@t��CJ�m��eɜ$#[��|���D��L�������E�hK�C��	I|'X�,�#�x��x���P�B��~�)�9d}U�h��>�_Ξ��L��))*�P�uwwK��I�9�_. �	��#j�4?����g�u.��̩�3�ϚIr�qL86�����H2,����鑋W����_ƷQ.��Zs6S-�N(�!��b�r��a9{r���t�!�
'�
�u��\Ǯj�m�7wL��7gd�50)��ʤ˪]vH$��u˴�$�����Y��FKQG����B�kƎ�A���������qR?+�.�4���s��</̍d(H����eu��{}�v@p_��ms���O�Bc��3Q�OBܒ����B|e��OI��c�u��T�^���1�tV�)�/�N��d_�㪷���X�襰��'�l�S�Hh�,��9C�j"��hn��Jة���e�p�5'@��Qܛ�p�EB}_�h���Ol��qW�,�$?��#����f��핎N���>ii�Pƌ����1a}�R�@D�>xDձzͦ`s"��i�;F�8��W�Ώ,�8�g�	1����b��uA����.z�
c|�S�c��2�Ȕo�@Hn7^Ǌ{Vr회k��AĹ�����B�k*++����~�\��WN{�vb+�}��E%׀0���aiy����3���c��u� ұ�+�0I�5ˋ�(~�ъ[f�b����*&�~Ʋ�Ya}�M�˼�d�b�E!��G�d┹r��>5�[J�륻�\Tu�@�/�\� `�I�M/�w��
��ҵ�Tf�ŷ�v=LG�y����>B6B,�|��܊;��ç|Y{m,�t��C��BP�m�b����k�6�	�/�K��c�I�:B!CGJ��l��!RT*�'�$��~(}�HQ$&�e��s��~�#��v���?��{�᳷)WQ7�v�l
b�
�b��7�d�n�������(����Y-�ee�neUی>I�X�5�`Q�*N�\c`��X,���p�������z��1�����B�@�8�!�p�9�N c��㇫0��z�m5&u�AB������B|�f�Jع��Q� �����6)��H(��r��8r+X0�D�[B7`��:f�n,Rv.�$I7)
&�8���M�2���Բ���dܫ�:�K�!�&�ւ֩ �c�^&��k�����9"�za�����0���N��� �-�)<�I5�	�@���k�W�߃v3HaCQG!y�ƥ�b��-�ʾ����/�����q��?�S]����hTB�L�+U��	�`����Y3�������25at
\)!x��X��8_XU~�A�B�ќo?�,�fW*���8K/ĉ���|N��s�}2k2=zU~V6X[q�ZHa4q�1�u���P�B�3�"t����¡6);s����$*�Cm��CG�����=+�b�ܸ]B��J�X��m��l��3��):#��K��v"75�o?h*M�)�Gp5u#��7^�:klU�V�L�sŽ��ӽ.���_��K�-�ΪJ
�:B�a���wjI��WE��UX�u����".O��e�-`1D���2�� ��jw�:Lt1��&ᢅ���+��"
�6���ǞE	o����+�a�M4�f�W;p�c4[1FP3.�v�n�R�g�x�JG�BQG!�XX���=&�?��L�:Q�a��붵�I&&�n,��(�48&XQ��I,چŷ�up��c`"����'R+��U�l�
. ���ڼ��eELtTɍK��Lpq@��q�
��Vu�l���y��B$}(�!�Ȏ�<��d]*@�!q�SWL=A����|tXG���qn��̻��Ä}ת/������l�3�*"�m{����J��v"�q�C���h�����b_XplڵY[�i��-j����5A�KQG!����q"\tz�\ ����%D��	���mpզW�Κ��چ1Z��\6�G�eV�Ź�춧
�ϟ��	k� �~�H��(�#��۩�����E�N����\;�.�*��z�i�CH�ˆ����E!�bb�C��N�e�t��ǉAܠ&�Y膋qD<�W�7T��o<���Ȅ	�O�V�+��o��6P�M�uy�dXE���ƣ{�i-�0n��ֺT��%La��$��B ���
[���uK	;��cN�ݖ����	�7ե��q$
v���r�� ����|g��S�~1t/�C$c�ML)������t�/�18�����S���⌱`���
�_�?-�(�!����t�b2�	0q��C;���,��aӋ�;u��:u ��*9
�]@w�3q��"��Y�L����1��W�b y�5q
\kO�Bk8w�h%��ͮJ2K���B�N�����l�v�
�򇉦������L�� ��V���N@,jk�)�x)]x�����uA~׮õ��F쵅.���+o����C�`[;�M����ݴ��,A	;�:B!d '�s$x�u�f���|����!LSu�QL���f�<%f
0
*�]�ᒉ>�+ӣ����A��ZE�3��RM��qg�bF�~���r� �E!�2�5{�p<��{�@�͙8ʳ�)�~�R����с	�q���d�Į�5�NHc��!��_������!�c����DU�.��|-5p�gG�w�vu�B��#Q�'�n�Ŝ��&�n-^&N���k�O�פrmR��9q^�Z�`�Lep�4�\�1�"��~�� �����������gm/�񡱳���"�㧰��#�BD	���M�[;ae�n�q7��gJT�9t�?���7{�?��87Ba�1�NU��i���%y�\-�r	��9�l�����3�{�Ə�uv ��J�r���cOu| �p��CY�<�K�Q�B!b��.�t~���L�MPHۭ%�0�K?�����H�X��:�Ŏ�������~Ԯ���~Ƨ��^�J]qxk��7�J�o�!�(�!�q6�Ǥ<�0ۻ~����z&�Dpp�1O�~欏Ȋ�WY���c��d�:?���͙�,f��9D.�,���uy����BqȕN�ie
�ab���@1���M'�Gkm2;V��n�]��k@������e�;l2_��hg��SH�_�L"C2����B!q`ep.�r��8����D�l����If^�[x%�(�!���ضBE��IA�)� ]��$��ɚ�U�:���	Ɔy���u1Ib�vu�BQ�:�^��{[����&b�PDz����"��lz�Kf�Ry�vhgIv���)��m:aE�.u�Ȓ��R��B"]aGQG!�8�67��0�|ͧzS�=(��a�m�>���Hn��5a���;h��5L�e4t�7���iRM�����1XDQ���KX�En��V}!����u~�U��=�N��]��\�6�#�(�!�q6�a̙��l��W���t�yX�|�)�e��L��}��a?k���).��p�3g�D�Gs.	�Ar<�CM����F�)�C8I���~�����*q@aW�vu�B�8���7wC�]�~���&��|o��M,�k�Ǆ�N5�섃X��j燨���c�G?���,jҭ]�(%D����ڸ_:)�ˤ9[&��p٥�/�;�:B!D��.t�~T> +�V)LFw<웋i�,�}��ʱā���u07k��	���_�m��֮�&�;|uw�<`�X����B qY��Qa�����s�
X��
���iҘ�)Ydq�%s�=w��Ch��hY���<�bj�X�b�L$�Y9� !�N�:��U��J�u�<�+?�����n�[�p/�f�˂ĉ���#�B������ŕ��k^΋:�+D��`R��=w���$���[f9�>մ�p���K �:^�Y½���&�i"��?�]�_ԁU�ڻ~E\ܤS�n��#��% ���K��6�O_p�\B�`D�"�x@}N��T�E!�2���f<��UWCX�y��/sU�BD����p:i�eԜ0���MYo��y���jy
�R��1�̶W���A׮s
��Y�q���@������3o���>�᳷Ƴ�"��	RH*��B@���?��a5X����k`b�{ս��`���G�DpA3'����%��;��	IV[#�J����������@H�p�m|ة��� ��&i��u�_WV�4��W�0k������v�C������6A�/�	;�:B!d <��S/�&��8�)� ��N�3pG��	��aB��J�ɂ"�oV�򖙆�IO�-�$�A�
E��Z�g����C����)p{5Ǫ�t3kj ��\��Z���f�$��]D
��E!�bt')��!W��zr���eF	�����mϥ�?��W��q"x���T��5՜��+^����[f�6Cȸ�7��;r&�,��j��s#v ���z_���n���
ƼS���E��<�$K�#����#�BL`��$f.%A�x7�.19�0��]�F��W��o �pP�@$8.�Hq?g�(%4�\���M���&c�f����\��u�E׮�L�v1vS�/k��X���ͩ�����5x�/_w�����{�1�>���N�Q�B!6����Y�@b��քl���L4a-YѸKe#t:��a��4q��x)3xx������F�i`��Z��o�FݷT���!�.Z���2��}��k���ƳٝSa��(!�L`�:7]�~��9)��XK�����j�xVaGQG!�X��w����L�1�#&�n3]��'�zB��21�,� |`�r
�t�d&��6' �k��i<�EV?�~q��e\K�?@��K����V��S1�kdWcd��h�@F�T3�&(0�����!!��XUl�����E�!DX�{ ���T��2gC�;���4��I�Y�Q�B!68����lv8�:X}��Lpa�q�7@;X\�ʊ�.�Ļ�
a�=M�lm��6�M`�k��*� B �ƣ�\!�!�>��p�*U��N4��w�\<qcm��ƥy)�����O�-�(�!�0�[9���lv�Y��v-��>��2���u�M�r%�V��Lgu+耛x)+�������	��$���c1��)�VAg�L�v�4[�܂qk%b���m]9��_nBR��BI D�]�M20��s�$e�ʄ�!�J:Y.SqC���q����D1e�g���K�A����:��"=?���7�U�}�����֮�p�����;�[�Z����:k0n����;�҉�n�:�k��̠�>��D�mY��Ld%�E!�� X'0�vc���l��Qj�dZr����(W���\� � F�Z��Fw��TeلE�1���4����������P��3�6�86�,�Nȸ9w�h[�O�1Ch�Z�eb�ly���K�Wh����$�,������J�*17`!�cJ��e�U��u�B�0@�����*�]1��ㄏ.U8���F%rp�.]�$A&�v�[���"�S�T�)��#X_��t[���y���Eg���jz����.���ע7�[�y����bH�[(�!��$�M���-3�q�'�^&	���uN�YтΩ`.1� ���ۦ���[&���nAp�x��3�?-f��t��BQG!�$!�T�f���dq��#���aW"e��*C^:V'�[A��J؁�b�w�V�]F?�}Щ��d�ѭ�e���B3p�����s�}\��7�N	]X�P� �l�@I܁q�4�3kL`�.�$?��#�"+���ݓ�(V.�TIsU�Ģ�!�V�*�J*�5
IkW�L��:p�C���H����O��(�.9�}�hA>Lܛ�I�Y\�b�"*]k��t�F�tNX�(�`�귞\�G 1b�C!E�bW��[`�k��g�^�@&��^ƒ��0Ǻ➻���\�t�A���t��#��F��[J�.I��Q7Nr������*��#fI���ɒF�TɌ�1R_\麝�!�||����Q�Q'9���Όj3$p����px%�4iX��
��(�84k/�=����5'/�w����fe���W�|��G����K�b���"�p����핮�^)�8�~%���_><u�߀����E)-�����M#MkHi�}'?��[���^^7Y6�~M��j�B�<쳮�Lm��;X��[��m�"Cȉ�$j���Z�(M?���e�vA㶦V*`�H��@y6��L�<���k��C  >�g�z/+K���V�v�V첏zJۇ��V��O�ȑ��F=k�:��Y�l?ky'$�B,&�KS,�i6��ɴP(<��	]
�M~E!��?|A��m�l\�@	���Nz��KKd��ý�'/�t�Ģ�r���?wD��kd�\�������-쐒<l0��uֆb���9�G?0�'�.qh_gI�˞�����x�r��N=;�=��5�F�!,��xS<����fi��� ���ZJ��%��C���iYx���R��d��C����3x��a���/��,��:�0��~���D[�Xט��l���DB��ZC�N��(�!$C�������N�x%�aB,���ݷHm��4�sƏ$�^��=9�P8"��r��n�T�ǬO�����˄)s]�ǿ��Aaw�;dGò�q���̠�`�>2ǆe;z�şqS�yX��/a��
d��x\�PBB�g�z�Y����k]� .��I~?T����j��6����Y�k���bL��=�I��f1�� ��h����v�m� ���E7�?���񇷮k6~����T��l���F��E!��l�Q��~ ��	���y^P5�Z)�?d���7H�كr���R?z�2:9
Yo2&n��9����̡����6��v~��������+�]�_�j*�>Ix��:�N�uՈ=�GK$Ա�ec�#N���������}Q�����f�9NJK�d��R\Z��1hA��)���C�Pr���p����'v��.MW8�"f�f�Xhc�_������o��5EJح���#��D9� �%�^ď�ȱ3�ܩr��o���D��HIi��D(���#k!&x�f�C\�zg���N'���9����\��:7����:	���~���Y��� 2p��%&�-�[C�!�c�Z*����Xo���z�p ����UŇ%Zo����_= �P�P�w���>��?K	W���0#�,�������9a���v�:\�s��M��?~a��W��񢓜��4��Ƶ��+�5�4����-��r������j	G���弜<���Ս��Q�����i:nO�_~e��]��z��EŔã%���XL��D�~w���խ뚍o�U�ln
K����L[US�BH��0_���#@��Ek��_��ܤy��vB�z��s2f\���a�G0&���������nX|[�-R�:m{u_�ʓ`ҌI2ĂrI3&�w:�^};�b�`��u���Ч8s?�2��Å�!n���Tv�\*��J��(��\Q-q| �М,�q,��q7t}�:�g�ƏG�Z��S�ں~�w�04'ځ�����h�$���87��קt��z���Ei�x.�*����HiQ��A_��W���uV��ij��ˈ1Cc��jF�����KW�>?y����������<�hDD�U�!� �y�a�߿wt-}х�ĺf���Y���E�pS���BrX>�Z��C��MU�4�D"���c�%%�3�� �J`Ʉ��dV�l���.}P[������eV��K˦_���3kL$��Y����eW���09�v�vq|�L[�2C����u=
��?5�(�	�ڰvM���>!��YJZ`=�����8f����Ht�:��,������];wXX�̥=r���>%��Vc�� %eu���%��J���:/nw 
� ��6=-~t[�tX�vu��� �%2����e%���'r��{2f�L)-���s.��&���z]�M��ܮ�G��}Њ��a����~<�O)A%�	
�DD��:�\&?{� ��c��Z*}����Gb�Dq|v�y��n��S�����U��Bf�=ރemH���ǃ�f���\�'��;���^���k*,}ϼ��%&F��^N��\m;穨õĒJVJ?x��7���w~<�D]W_ty�NaW��憈��vu����Ee���)� ���RZ1�vQ9s�}1j�T׌�&�*��ٗ������aV�@�`�	Q��������@�ud��y�$ی���I;��~�m�|rV�� 8ஸb�a�@[oͥ���J��5?����4h��cC�S�o�|cH�����C|���a�������hF�ˏ�O�O��i��8��c�z}N8fm13����Y*��"�������S�9(��~¨��<�o�z8��GyE��Ec���7��z�������9X�𛇤)^�aF%�еu�Q	�b�<�u���)u����	%�Y �t����}i�,���>Ǡ��.f[\Z/&�(gO�+-����q�IIi�tv�I_o����O�{�;�P�N !X���R��6�[�E�%�w,�ﺯtY�������/���1�|�d�8��+%��g���h^���&Xo�R_���eþ�YdC|Zף��P뿶���X�;�h���|���}��e��rN�DKK���뤭�tuu��+��	1)���~�QY��{q�b�3ǔ[K����=�n�d����ƚ�p�7L�:B�1�J��hA��a�L�aW��i�I�)9{� �?���Ĥ��Lm���Duo���t0��|��d
��q�h=D�]�����,���'�7����\���J���f���땓�ޖ1c%ma��^�O��N��*ɬo�r�zEW_�A2��uͱ��׆B᧜~���Br<�D�8��/�K
���?�}� �1�k����늴�����΁���W!�d7(y0i�͆���!����}g�Y��j�n�����y�����$va:6�R`�\�5�x�d�b�|&�.���]�#[�8��Q�BH�J��A�Y�d��(k�����3Ӡ�mEu����D RT*�+a!���\}�n���Ⅳ�且�����y-;U��lvMkHX|\ǉ�"� ��	�w�E%{h��uu��#�GOo5�����E3�v��B��/���4�όk(!�"5#o����?_^Q+�ܤ^_�xH�B�bє����&�ıX1ǉ��.l��x�D%�%􆣍��0E!��*e�R4�'�)�47A�-}R:bp����}�iU���"Ο�Z���޾��K�IiɈ���KH1~D!�xO8ҟ�S'�rC�!ގv\��{;������W1N*�[%U ��bib*Fn����.�4������e0R&&M�E��A�#[�8q���#�"_�����@!����<2^��¡6	������{]�]�>k�+cw�;Kef�j<;�`]s��k���@e���'%b1�'��fH�Ius�:B!�B򈯿|ɲ搐�D��&�2 4Cu�B!��D:��$%B���Vq�ِ��B4u�B)h��A-��t�*�: N�?��APZq;�����7��/a=K�Rݞ��B!$�h�u�O�!�xE!������ 0�wm�z	���m��zw?kmB�(q����뺯_HrT��E�%.�[^~K�;BH�PY$��%�2`���⠬+E!���+��$��M ܏^��jj��B�B�@QG!�� D���\u8vZ蜃~C��pi�	!����e��.�yN���#�B���X &�MkP�ސ�F�`��N�BH��T@BH:ٜ��BI���ar�DX0��K&�7���z�1�-�N\�F���_8P~S���y���:�E!�Y9�^�\����*i�*�X46d۪X�TI���B!i��	�c�U�u��]v[�t<�NTq�Lԩ��-R��6x��<�|�?�bжX���2-�}�D��|�D�R��`u���ie��:X"�Ȑ �*z�X?����^aB�VB"�U�l^���u;%(��F!�<t7����?\U"�G̒v	K~�F�TɌ�1R_\麝�!�||����Q�Q'Y�tH�a�v�?�g`�N��6�_��Ab�襖�k���w�L&,B}fp8_d}����j>?��ZQI�!$�	ǔ��
Qg���u�B����zۥ�r"1�®��V*J�=�w.�|��oӇ��a�J5a����2�-|m��ji��e{~a��c�����8&}�Zܚ+��gt_�<�4>�ϛE1!�d���S�f󴮭�f�8��on�����(�!�$'�������#RV^#c'��zWϼ!��.] `�3��Q�d	S v��Ѯ��7�����.��l-`~bv�8��� ���A3Ě>��%���f�����[r;E!$�)���$��uk6ׅB�-n>JQG!FOz�3��A:6
�[�����R�/]0d��P8"��r��n�T�����;}|�L�2��>{{Z%WЖ2;+�ov�.a�]�p�2� �jVЦ��m���ǂq�q��h���$��S���猯#�d+��ܝ�غ���F7V:@QG!Y&�:)��pC$������%C✴�&�n]Ոk��r���#F� }gʥ�K���ϘE�-�t���D��oZ}���k�������D�K��)�N[��p�i~㒢��̈́%�X���W��n_��BL�n���S�BH�0����DJ���D�v�3'��d[�@���;SΝ: ��V��K��~���VKQQ�J���k���H�0�3K&b��2M]EY�u���a�� ڍ�B� KYQ_�Q�l^([�5�&J��F�i@QG!Y,m���n�=�o�*�ރ��v�H�O��P("�&͓����sU�Z�ɘqU�%�I>��tN�g�GB�}B!��&nj	@�A�E�Mn�.5u���������b��=�o�j�I$����Hoo��DJ%_��Ji�V�T����%����K�ߖ1�u�l��X���H!f���}ts�_��p���.]A(�!$�Ѯ�p��r�gd+�q�DN�|Oƌ�)��5����t ��M%�p�L[gFתõ�u��@G��g�A'OA;*qO�̖�w��#��v��U�����'��*+�-k6�$EqCg���B����zx���Kx��02)e��%�Ҋ�2aRHN�x_F��&�5c%��צpis�:'�"��ە��>�(��|LUV7[�(�]wO�ډ6���LQG�5`E�b�k�o]��nl�޺�t���Ѕ���*BQG!Y&��7!6�Ƅ>�K�F�"ŵ2a�r����r���w���VJgG�tw�KG�e�]o��I52���޽�u�g��u�F�$ ^,RwH�)�%ږɲMHv��e��Ue'k���k��5�d+n��$Y��쌦*+��dU^'��b{[2�SQI3�K6%Q )RE��w�{�y�n6�@_��sN��S�>�o������v��t%@��_n��Bz����������ņP�3}O����oeQz�~�:m[�����p��4 H*mw�l����ϳ������ηӦ�MM;r�pW�a�#�@L�~�P�͚e�=��/���
j��*��knYk]�A;3zԎ}��M�6?7c�T�֭=;�j6�T�ۛ�7�W>��t�s���_�|~ۊBzl���O�*��a,������������i�80�ʫ��7_�$S�KYz{g�=�U��ڀ�2������6m˅�n�Z��q�����P 1����j����cbjɕ,} �֨��W�Tȋb�3�����2�5;=b�G�"*g�K��c��t�c�!�/�R��r�M�����3�v���3Xd�R��9���{ k�ͫ��G����v�s/�Q��1 �$.����v�]��j�'�P 1��AA�����2����{����w#w�(��uZ��y����}MXSs��F�g�֙Ry����
��z������n��_8S!����\�.u�
�? �vu cj$�\s��qK��5��2����q�W���*��ī�L|U�������ﱗ  A"�@���-5�MN=3>�ySKl_�˞��^w��0���vk[�9����옵57Ys.�Ukzn���3�n�bm��/����{�  @eu s
n~�O8pxq��V\jޗ.��0�����/�~a   �u �R�p�W��+)e�  H>B    $�    �P    	F�   �k޴iӖU�VE� Z[[������է��   ���:    H0B    $�    �P    	F�   �#�   @��     ��ޛ���eT ���徎[��Z�j��ի;g3Y����c�T}�Sٴ�6Fg�   �W���s�����z�W֯_����ı�U�����7    ���K    H0B��L��`G�}�   B��d�[m�k�   <�:    H0B    $�    �P    Q.;��u��~�����vz�Ł��   @b(�m<9hI���ӹo	,��    �Ԯ;>d��ٺ�졲nW��2��    Ԍt媧@��u    B׵�����{��6p��\sYɷ��@��u    B��w��Ĕ���?Y��?]���9�y�;B   ���?���~���\t���t���L��m|�ƲoK�+AKK��}�n    *Rn��5g�������r�5�<��/�ۋ߷q�   @��J������7t��w?��^�2    ��k[/��_eMM����Դ���q{湷,w�m���\����N���=j�<��B�+����a�    >2Y�3���eK����q�'��С���_�;?og�L���P��׏Y63oa"�   �;~|��o�tA��+��L&��)�P�?>d�ׯY��#�r�6B   �:���ǎ��|��K3��w��(7�@'�:    H0B   ���}�G���     �u    ��ɡI���;粖t�Z[[�-��H���s�mj	�\!�   �o�k�O�wy:�d]Е�)�����;�r��(7�+w���P    �R�-�$���c����l�K�����fs�Y׺�&B   �D;�����7;r4�r��x䰅�P    	F�   �#�   @��    ����]ikϜ�F�I7���+�-�   @,��pq��[������)нv�'m������    �V��j��    �Z�� ��    �^�����    $B�� ��    $�v��;hIu��P    Q֍��Փ#�TkΜ���:    �C��Ɠ��dg��޲��X=B   �D��@��u    b���T�#�   ��zt^��P    ��9�y�;B   �X���+u�<��֏��ڍeߖP    �֜�F�>>L�   �FC�   �h���B�~�U��T<�LMM�˯�g�{+��"�   H�L����m��e���G��i;t�e��(��   @����ö~C����Q��z�2�L�0�UT��
�   @����c�mn>s��+�r�"�   @��     �u    �`�:    u��ФM�̝sYK:c��-uY��    ԅ7ߵ�'�λ<�n��.���N���\�P    �R�-�$���c'���3�pU��u    ����K8j���Ѻ(��    �P    4{��zo���V���������d�   @(�~�N�'����OX��N�uǇ\����'� �   �����^��G�x��{?�.Wo���rN��J[{�5�L��F�_X�m	u    �s�e[z
q
y�.��]���sz�Źo��z�@���������nO�   P3�C�e_����@'�:    �V��.�@'�:    �Wo�.�@'�:    ����a;n����/u�8���)��tB�   �SW��Z%���S6�wВ��
,�	�   @�/�ޟ���oS�uc'����w~i�/�@`�G�   ��S#n/��]v�9�xrВL���Վ]|} �G�   �������ꮅ��!�   M��6���	�z��e���z���-�����+Υ��@�]�喪��   @(�]r����.�i�q�t�����l�(:��D�#�   E��?�kn��+�]w|�:��)�)�����N�niPρΫ6��    N{�uo�t�.�����w]�{�����i�{��W�>�y
v3���˾-�   @���J��y��PKm]���^���U��ǚ3C�H�Ǉ	u    ����׏�C�   ��)�]C0����)�g���۔�׶^h�o�ʚ��Ǜ��i{�����soYP�*��   @�|o�F���'��K�7����[�ߦ\��ٙ�Q۲��Z[Ϗ8��v��Q�f����-D�   8��i>���-��i�KͱSo���=z�����ö~C����Q��z�2�L�0�UT��
�   @(v}�	�3�P��
���_8����r�x��*���ǎ��|��K3WT�E�   ��6W��}�G.�:�:    �Q��6��(�s�4�N�/�KW��8JG�   
ma�M�5gN
C�.�1����U9��q�    �B�(��!�O<{�������1���){��̓C�6=3w�e-錵��X��*Wu    �a��[i]�վjq(f5��1��?1t���t�]tAW�pVT�z�:    ���2�ݯv�-��B]�6����e�+�d��؉a��6\EUn!B   ��OL�x��=�Ɓ7��pԼّ����-D�   8�4�n�P�B*�@��P    p~�V�\)��a����    N�ϕS�R���חB`5��42B   �P���nh��,����F�u�:��~xf�x��]�!�Z:3o�n�m������nK�   ���i����;o�7n]f�i�����-4��n�]�ɺv
t���oO�   �5�S�/�3'
t�̡��`Wm�B   ��P��d1�zvA:!�   \����K5p���0�ނ]P�Nu    �@���O�u��G�V�,�^�]��Nu    �a�Ŷ1X�6+�����;�T��rY�   @��G	��]��(�u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#ԡ*�O��G^6ki���dldU����   ��UI��ܻGlÆW�m3#�  ��P�3gθ�qv
t'O�4�p�   ��P�@�`���iq155e�N�2   ����������1   ���-����Ӂ�_{[��tz�   ����6������V�ܴi��ޓo   5B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�5���_e���N	�~���O��mz�k;3d  ԃ�-[mt�U��:4�������\`��~z� �����w �z0ٵŒ�P��06l��S��x   �"�   @��     �u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:4��-i�⥭��ߦ�������   Q#ԡ!��ͮ\���6�m3    u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P��0�1;8�	��F�L   �:4�S��Gf���#�   �:    H0B    $�    �P    	F�   �#�   @��     �u    �`�:    H0B    $�    �P����)e���~��Ρ   �F�k�;8>k#��@���l���u�)�� CݦM�u   �B]�8xf���ա������   ���     �u    �`�:    H0B    $�    �P�Ě�����)�d2���d�W��T*e   @#!�!�����,�ͺ���͹�u���   �PuH$���@�)����X[[�   ��P�DҐ�r.   ����9tn���   @#!�!��(����9=s---���j   @#!�!��JGG��C�W�$�  ��X
v�.�rl:c���Tp�x�   �8 �   @�����q;u��Ess�uvv   P�u��ɓ'-n�w݆   �W�:T-��N�����v   P�u��l{��u]`]�.���fl�}�   ��P���n����{-�f   �O�:    H0B    $�    �P ��ؖ�6ٵ�  ��]�-Iu ���n��  @4u    �`�:    H0B    $�    �P    	F�   �#�   @��     �u "u���?�j��Z�lr|���W߱7G��> h<�: �Z�����T��e��Ykon2��� ���     �u    �`�: ei��#G��d0�FO���>bsss��MNN��![31S��gfglv������X�>/~�)����N<�b���-��,^�������W}��S�vf����}� �x��Pw��w���ޠ�o~���-W�u��kÀz� r�/���)[7L��>d�����uZ0�^{��_�/'���P}ڤ����]�7��`J�3��5{��]} Ш�6��(��yPw�>i-��r�PO��T ���ٮ��zkoow��袋������>|������CCCv��	�Fww�vs1
"���U�V���DC�'  ���Cݢ�����3��9rĀzSm Q������mݺ�.��[�~��.�`���y�fggmffƅ�~<x�~��_�L�D�P�
z���� ��5D�kii�իW��U@�K��O~�~�7~�� �.?p^SS��]�v���7o��o���8���ةS���^������z���� ��T(Lz}  c��0���G��m����*i浸��[յa��f�-�И��o��� r�ڗ��%��C���J��
&�y�ץ�^���v�m�ٱc�\X�>�"�'  �.D�Sǭ�����!YRss6;9i-s��8;H�:�� 
����k��~���f��׍��K�N
%���'���_1�DD*��/��.dEY���/�b������v  D�!B��h.I����5kָOÑ,����u۸q�ǩq>::z�r���� �s����	s��%�Vٴi���SQQ )��A$���!�q�O  p��ujt��4Tjݺu�a�dч jH��4I��S�+5�h�������=DԋT��QHa��+�t���ۿm===���]�A�����W���Q�  �T� ��� ��G�Gv�w�@�!���\�e~��_�����+��f�>	v  ���Sj ��+�����2�q���Y��'O�^�k���y�%�#�P�;  j�P�� �}�v��?����I�ya�@��O�ľ��o-nĝ/� B}�  �%B��J w�y��ܹӭ��\�ri��B���z���/�2� B}�
� �� ��� �T~я��D�O�  Q ԅH��k�˹��Z��A>33��V:.��}�)�xa�` @Tu!v�;��K�m���J���_C{��뮳���߯� ���g��7���q���l}>���gϞ%�#� BЀJ	 ڣOa���'n��JD.��"������kK�A$���e~���?��l};v,��  �!�huk��72\�z�n�!�Z�p~~�������̙3v�7ح��jO=�Ԓ�)�=�βo������p� �  ���� ���O�n��7���w��7ߴ���߱�^zi��`Ah��ܼy��a�'  8��9���j�җ�T�D4gR�n��u�h�����K���_�> ��u 577�=����!��a���\5,R��������4b}j~]X�	  �F����o��۷�U=�����p�|�w�}��/�l} ���B��H���h_�z[�g����`����~Gջ444d���'�����>��`�  G�Q*�r�h�m.����s�aU?�2/#�%׶m��p�F�U�BN�<iw�uW !���> @q��)���<�b�I�Z[[]��sW��A��g?�ن�U�|����ȲK���> ��u����][[���k�mRhԍ7���A|Æ�����>���B�yVP�	  �G�C(ԛ711�z����d��$���>g---�Un#�.��N�8Q��P�gU�  `y�:�J�0���\��B^�a���f����:;;�رcv�m�������oO}����  +#ԡ&�&''�'��wG�7>4�Id7��Գt���馛*
!�繪�O  �2BjJ+�jHZ{{;[#���?�qzO�h��ߐ\�nccceݞ�<W��	  VF�C�)ȍ����իݰL���*��_~9�A���ڒ����%ߎ�\��S�`�[�  �4�:DF�1�"*Iok����>粗�o��Sc����!�R�h��+�����Q�竴> @iu����t];=���!K���.���K��U@�e�֭eݎ�\Z��	  JC�C��%�%х^ȼ�"�������,���  �!�!���Ӗ4�k�R�>hа�rP��UR�  �4�:Ć��iULŵ���|�Y�����Y\%�	  JC�C��`�>v��J��i?E���y`�<�zI��>���> @iu���MMM��Q6�������cY���  �(�;�ӧ��   ���f�繯�l:�|�l8��tֺS��6�ZO*e7��Xu�%��i��   q���e����_�v�u�kj�M���Rf���u�%K  @\(�ͧ2{��=P����3ۛ�i���r�.�'�pG�Cli^�u �ѿ��oڗn�΀ �N��]����K�޳��\G�?Ͼf��OJ:6k6�ͦ��=���A��z�v���hv�n��P��Ro���K������d&>���ˇ��o���^��9��V��7�x���P��UR���/��8�\��cU����>�����Ѩ�:bK���������e��5E_�k��N|c��>�}��s������7��t���Y�]�kZ4%�NǾ��Ԧʟ�;���[�Z�9sư4�k��r��,����W/ƨ�GaN��8�\G��t~*Ѝ�gz�����3�ܽ������Lz��`G�C��f�<�B3�7==]��N곸J�^��3���3���6�����M��\G\�t����7�^�����<��u@v��s�}��������nG}.����gjL,נ ��:�Fs��3;j�<�����6Y�{������!�I�r��	ۼy��W&'�·<p�@Y��>�Vi} Pk��N��=X�r5���}�*]<�P��S��*����������]x��o���q[�v����Keݎ�\Z��	 @-iۂ3��U��s�=���J�a���_��(�h�JB�+��B}��>�ֽ��z�����z�  �mz>��ط{8{_߮T*�p�7%�!���g�yƾ�P��3��~��n���O�W��U�sA��5��_��^?b��F P��Y�~�.i�����-���P4��'O��N�^{-�挎��ᾕ��Ҽ:��W��O  j!���[|�[�s�uH���GC�^x�����mnn����uvv�O�ӊnO}�����U�g\t�nsC1�����,#�������.y��^�]�}��s��]w��n+�ձ�Cs���y�}�C�.`�����/9��W����7]m�_�t�Ǽ�g�������=N�I�<��	C|���?�W�����λ^��^瞽���Z��v���%o���}��ӹ�O�n�ۭ�^Uʹ^x��K.X�L���'�]�,=Ϟk.[|.�>� h�K-Tb11����d҄:�z<���O�=����C��z��ۦpV)��,էzYM}����h5h�&9���^�2�0G��>�#�X�ԈU S��u�.�u
{���Fr�S����]c���j��q�k�z
t����K)<N���+�qc��x�y�����U.�K.��^�R�\ra1wN(�W�*�\�?�{C�;�����������_�^�<��dm�bD[tܿo��!��:$�B]SS���������SO�G?�ц����{ϭ���c��1�>�
�>�QC�	O�#5
{C����rz��^G5Luu-�֩q�Fna#S�X5�ըu�s`}w��5�������!�u��U#</�U��u����a�ნ�PJ=�K�:��
G
T{K8G|��,(����s]���u|�{�������?�=��\�9^��J����ō�f��.�pB 7L�?��m߾�aC����
j�o��4�����>��8���,��@԰�A�5J�xv��\#:���5t��o��P���hw=u�������{
���!��{������F��:��Jy�ѹ��T������[ι�WK=�bCKWR��J&���Q�L� �뗿��k|_w�u9�Q�h�����'�ܟ�S+a~��l�`t}�� ���z;Dp��z�
�\���?�R��+�=�Oe��}T���^��R����+�Z)������T�ܳe�#�uC�B��YN�+�\_�ia�f���"�!47�yuᚚ����뿶����j��`
]
!���r��Ͽ����o���L05X\/�Ĕ���G
����<�K_5�ESw�BC�ͽ\��+��a����\,u�_���{�D��`ņ�\԰��#����W˝����A��z�^a-@���_%��������T�a��^��:$F�0C���7�\�cǎ��ի]�l}.E_�;�F@>�*�]�5���䵜��`.�R��0�{���?S�<*}/��Q�B)~�}���'&c�=j��?7x�綐��/~8b!�G�78/���,�}��s��{b��K}h�ܪ��Y�y�|�:$��Ԇ�=��Cn��64D�VgԊ�~�i���p�ҩ񪆈�����_V������]_t�g�B:�PWw�9��ł�B���o��C�<݇�~5� �I�~�(�����z+_Ƙ�S������9���ߋ
���M�u����,�}��s]��yr^h��w��4۶q��
��L��ҥO�C"dzY3�N���~���.�s=ӰH�T�����|'�2���}�j��3�O�Y��q(��!
{'\p�}�o ~�\a�ׇ8?�-(n��>�zF�CS��<��{����o���r�l���m1p����Ntn�+<�6�z �R��{Ҋ�GW���BŞ7�G�C"�|��Z���/�l�z�c��������v(��y�'�\jh�p���r�����]�6�2���0�{����[e�Rz�s�@��o���Ph�[f�e:�ԳV���Gt[d,(�Gn�\�/��R��r=���=��7�x��n�VU�g��J,����z�b�S�k�n+�xB��g����v��׻/4���l۶�n��&knn}�`~}����e�]-�s�̅�rC�)֐J��]��g>rvq;��T#x��N��a�����Vl��R�p�մ^�7cY>�-L�������W��=`~%�b���=�Z�d��]de�����:��A��Be�|b�g��C��&R�S��:Ğz�OW{��1��G>bO>�d]���n���m����裏֤L_�����π�O�}�F5DԘ��c���QH�G�׿U�m����_��b��󸫄�I�W��`�J!;.d�PJ�큘w���JC6�r��r��W:��y���CQf�
[�}�R+k�BbO��h�	ԞBH{{�}�pAdvv֒n˖-��/~������d�W>�gkk+�����n��S�������\ H��Y����v�����͙toٷ1 �O--|�y����$���^��K\ �bޗ�^R�ɡpX����߽��}-^6T?=� Ј�Y�b�rz˽��F���zvq
 �gr��'BZ�+S�����F5�,�@�(@�rMλ�v�uO��=��Xw__�z˽���E���]j�߻��VOD���'>���	�"��[�e_|ql��s�ƍ��O=���q���X�ƽ��Wc��l�<-��a���G��޾�D(A+�2�G[S��"�_���+�J�䦄:�ZRz����;���-[��U�V��>�1{���ȑ�/@���cw�q�e2���8�P̵k�&�>{,���4�o���t�?�-�}��{r{2��~�o���
wn�gd	�V��w����Ҿ\Z������(@�䚝ۣ�[�ќ�SI/��[---,�CSSSv��	��[\O�+����Ԯ�.�o��W_mo���=���G�@`bb���F}�G�c
U��������Es���[�ma_1��-?�k��ƾ.c	�`(4��L�ڤya�������j����L �t�}=���|-�U�����ޞP��R/�z?z]�p�M�6�s�=���n��Vף������~x�������g�*]F��Q��ˆkX��zs|O��S�SO!�0�燺��%�wA:���{�O�)k�O��ξ۷{�ej�t&Wfu�%ͥ��.���v:�v~��2��)*�/M��뮳W_}�~�X�P��P���!s�s��
r^��'  ��J�MM��;��Lz��a�����g���5������.G�S��52�k�f��뮻���_��4��𡡁'O��|��jP��ѐ9�ysA��#�����E.*�6�^X8C�mǍ[�����Ш�4Գ��;�r	� ,����k(��\����@'�:Ďz*��hs��to���<x�:::�s����Y��)Z���k�uy_q�v��i������˙���t��o��g�J��Ri(���K�+ĉ������^5C45oם7�ysn���B
Q
z�c�r�������������=��
7|�ֆ�Q�	 ��ԋ��o�{�k�J���}]��T<�����@e]�ɤlUkk(C\F�x�7'��nsaGC�4G��@��^�_��_wD���>��[92,����z�5�\Mժ>����ի]��^�T
X��la��k��G=X�S ��_E����_��S�{�����O.D�Ebr�ٯƩ���R�/%�ߣ(@2�-���uܷo�|*�g�����?�]���-@�:Ć��Ԟo�;�����W��Ұ��f�n^�(�|�����v�����GV�_j�G���/mr��".��R�k��"r~��[����܇ͷ|f��jU����YAY��~�z{��W���{,��Jܐȼ��n�d�2}�}�G�-Z�zs���_�>�|��[~/�׿��u�.��Pņ�Qn2�V���GV<N�r��@mh��fK�,�~��L�ؼ�/u��65omjڑ���s��2��������+��ȻvIg�FFFB_eT��رc��W������W����y�fף��ﭷ޲�G���ZR@�ܶuw�w6�~Ӳ�FU��N�էz�4�qfff񶱨϶ա��`T�S���D���W���PV��^{>��Bd�P@?ɣ׵�zM��<��p�����f{8����Ke3)�?.�mږqݖ������q��S����5���[��.����̴k��z	8�t��o�iq�zP������ r�m%����e���LOQ�*��j9�M�N=cjt����]_�=?|r�gG�R�S�~ΠGa�R���zE�U��e���LK� z.����v�]���RB"G����+>�ֽ��5�N�BH�-�QK�]k쿽�s��|�O��읉�����1k7�\�QK]vm��\}��U[��P/�B��WM
�P��ڹu�婜Z���Q���ϸ�Q�79wC.s�_ϱ^�Q�\ũ�L����~�?�"B"U/�Ns�^��K*�J�%�쳿y�9�Gh����e�Ƈj���7r7�炀��X���9�[,��E��nS�\��:\=���.|�Q�\ť�LHh�U�s � h�:DBaNC�V�.)���ؚ�v���� C�R����q,�H=�@�a���F�蹪u�~S?S��T�z���:�\nOI��M��{T{[���,ן_���'�5���^˿hL�C���{����#�F�_�R�/saÅ���!U���蹪u�~���v�EE>�y�|���U8�Y�Q����>���^g�ޤ�ʿ?��ms����x$��+}H�r�3��C�׊�"�HB��E��n�΅�W�{��&�b뙨�P3������ ����O��x^�����M̱�E%�>����C�G<���yznK��(k�)��TY*[�}�a�FLX�*DUn=WQ�����ܗ�p��^y�� TaG�K�g�;{�x��:�s����"��Q�QL�!^�W8��-�p476��k�Ø��-�*��q��u}������[����.W���?��~��^ޏ��?�A�;���zE�CM�;�b@�����`4Z}��Cr&5��/����	�f�¥6����h�o��j�y5Pܢ(���k�}�3�1)Ć��e�Q�\E�[�yQ�CZ���X��X�7nue�įt6^<o�ӽ�_�p�[�=e>䨞}o���?�¨g=W����P���|���*pz��<��P�P)�i�z�; >�'����y=F>�(x�J�qmp�aFn��\�M��Ay=�E�U#��E)���qs������~��^�b������\����z��ʵaЇN�}�=��ĉ��> ���>�C�g��.Ե��~��-H4����|�P��)�i��0��"ņ �rטPO^�q5X��X�<�c&j��b�Y-ʍ"HG�]�7�WR/s��S�>ȅ߻�7M���6�p�@�>���d!�[������Hi��Fa���繑����U����;�T-������z,n���ߋz^��P����g�[�<9��0K��[�P�b���\j�q�O��	�c�a�]~�)z�~�q?R�*�O��*�P�v�Zͮe��R��z�%��7?�i�!�a.���O�]�y�����p�?����ͽo��^a���
�ş��{]&a���ɇ��^c?3L�����ܞ�C�5�U�ר�zF��z��k����)+��9���8 ��FB�m����U4&� �'��F�_|��SQ�l��A����Qܜ�\�8�����\X^���y.����De*$�h�����sɯX���lj��U*��9F��?o|�Q>/�`L�<�d�zN����}�E���s\�%�5����Ι���{~�d͞o�u!����Ş, @p�<�\�*�@��V3��7:����A�:��[���WI�����q�XT�_ �phg��}A�勢L)܇p�,��W��
{��X�)�*��u-,7��^��*W=Xz�U=�!��Baa��Z���3Y�����#�: @"�/*��e��s��~uK?���Z�����*2o-̍�����a�����'~�<?-��/k]��� �����
�;��!��N��[/�F����P H,���Х��9ao6��?�%5N\�]�5S ����Bm�a��i��ד��	�F�~��r=Vn�b�q(��H���|Q�%�K��É��n�\ʭ7>��gB  �
����Z7��Z��HX��}��6Ȁ�XX��-E�+��綰a�/�os&�x�S���(ʌj�Z�y�6�Ν_n���s-��E����r���P H$�s�����\�j����σ��\n�Ͻ��+��޲��\�
��_�����J��T�]����.���	jq�(�\NT���-�s�틋���R6�\ʍ[�Q*tB� $�r�D�f��ׅ�"���x��v���ܼ>y�߰��9Uf�\�P�ϛWX��w[F��s=�R��"4>H���'�Q�����!�_�ޯ,�K���:w)�r��R�Nu �D����Ԟ,~>��G�c�sH�z�
;~���h��}��\��y.X�\5�t�~��9�z˂|�(�P\��_E�m�P��ԝ�!��\ʭ�ߣb�Nu  Ĝ��V�e��>�x�r��;������[#���}��|(势O?�0_�\�$�)Q�?dY_~�B��~�iX[�P.�&�r�Nu!�>uڣ��6o�L]��OOO�xܺu묵��  ,n���?o�u7��,�^����-����(S#̇J�x�\�<�2��0.|�s�2���Z�F���+:!ԅh�@�����Y�k� �M����Q������Q�r�J�
�5쵪u���C�h�W��e��\ʍ�R��   Q5�)�r��@'�: !�Y�y�k�R��L��Kg���R���oO*e7   ��@'�: �\��L�ؼ�}���9t��ж�����iG.��J�]n   H�r��R��Oe��?�{���N��=8m�7���u����R�=�;  ���$�	����/�H6��3����qc�}�;�]��i@ >�y���͵س�Vʥ\ʭ�ܨ|�חr�ܰT�!B��А�>}�&e]u�U�?oܸ�ZZZܶH��A{{������Yss0�F٬�0ה�����-H�v���Z{�@����p�i@k�N����ǼW�}��C��K�+��܇>o�����[�Q�U�!B]T�����.yִ��ի�=nvv�2�L��)Ѝ�gz��e��U��7w�o���9� �  �C��Nu!���6�z��������B�̴��^�e���u����|��^���H�  �� ��6B��ު��A��C�͡Ӑ�0{�
)ح�������3   D"�@'�VBD%c!̡+��bvܿo���b�!�AI�Rn�1�R.�_nT2���[G�!�@'�v�m[p�����*t.���9��0L�D�Kgf�mbb�����͛��ň(�r)7�r������:*7hA:��Pw�С�ܷTP������fK�̀�L�gz#} �vg��ەJ�6`�$���٭[�R�T+Ɩ�G�r)�r�/7*)^_ʭ�r�F���u@�e��}m���>v���KoJQ���?��K��[�r����K�uTn��
t��w��dR�~��~cnJT�� ��R.�Rn�����K�uTn��t��w ��*���Kg�[2iBJ�?�'O�����ߺ��@��R.�Rnr�mM���[G�+�@'�}w �*k#Z}���}#�D9���sDK�t4��
�K���\S���[G喪�Nu@�e�V�-V�����   ��U�BPc�tf�bFA3E�  D-��      �tB�jl|.~�/�{����   *E�B     �@'�:���4۶q��
��L���  �"�   @��s�b1�K�l�   �u@��2@���   �H�:��b���ۖ�X�e���U�V�t�5k(�r)7F�F��חr�ܸ!�5�2�\{ߎ3�ܽ�b�9��5���x��u���i�\ʥ܈ˍ�^_ʭ�r�PD �uA*�.�׀���͛˾][[��^�Rʥ\ʭ�ܨ�����:*7�u@R)��mg_���݃Q>�u�����ЀT�ԫ�)�R.�V_nT���Rn�g�: "mM��i�p~�ξ�T*�׀�R����z����P.�Rn��F%��K�uTnꀈ�ޗ�G9���9��^:�"�N[ss��:u�r)�rVnTҼ��[G�&��P������L|c��,Wa2�vP�l6k333�K����r������:*7	u@��S�<�}=�o�p-���L�L   �B�T�n�hJ�� �)�5g��  ��: |��{��7���r�:  @}!�1�`�^�u�}k�؃_nUʝ}]��0�+:�n�=���/{̧:˟�>4�bώwX5(�r)��r����~�ߣ��Q/Z*���oߎ�Tf��7wTsn��t���H��K�	-7*���K�uTn��v͖�Y.��<k���y�_�|;mj��Դ#w�   ���1�����w6��Y��X*3�I�`�q�lӶ\�붬�h��~   @c �	�^���nwޕ!.e   h0��inS���    
e����&ԕ!�B�pvh    �IY(�R��PW����S��3    �3���GU6��c����}�y3    GC/'�����Dط{8�{��T���     G�GY>��Lc};�hch��   Ț�Ӣ�Q>B]F�3=M��   иr���o���� �Ub���ѝ}
v���   ����.�Nu�R�3�Yw߷v�RYO   @.���Lo�C.��4�����ξ�uM�#e���   P?�r�2��曻�[���kQ�f핹    IEND�B`�PK
     @^�[$7h�!  �!  /   images/a7fde0f7-2836-4f0c-aad0-66dcccec46ff.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     @^�[Y�u�= �= /   images/1615224e-fb94-4bec-8b91-0567bb6a6470.png�PNG

   IHDR  H  p   ��   gAMA  ���a   	pHYs  �  ��+  ��IDATx��i�|�q�u���_��M�HK#[�bˢI�A"C���v�	$@;$�����K>$@Fx�h�)��XD�RdE�mj!-J$EJ\ɷ��{g�r�������,��;s�S���̜ӧ���_UW�Y!�9ә�t�3��Lg:ә�t�3�2g:ә�t�3��Lg:ә�t&Og�Lg:ә�t�3��Lg:ә��
ҙ�t�3��Lg:ә�t�3��3��Lg:ә�t�3��Lg":+H�,L�HK��,�9�ș�t�3��L��3�[t�K��
R?����E�0��� H���}�>�:�	7ӟ��"4������(Z��|?%��̔}z"�Х��sR�=��K���C;�6���쁔�KC�TF���������s�7ç���k7�~^�q1t����]�cN�)��� �QZ0�g=_�o�7��|���.a�3<c]y����b�����伵1g�ڕ\�0�7��Vn�i1 ��޸+.�1��Z�^6�V)҄|��-e�k�\�z>��+�����U�U����|gϝi;�c���{�g�L��a\�(2�!��O 5G��%恌a��+ �,�+#�4n��U�]�N�&�'ګ�G)��M9d�K�<�d�_N������Z�"n������$�.)H�+�"��W־��ھ�jc�4|xm����4�������'t���:7��sI�(r�NeX�B@�z�I�	@g;��mXL�ic$�iG�T)@)�k�	�ey��0��s�Z\)�U�FB9XF�Ss������ʳ[^!����`]��i�r?8m;/H�0H�l�6$L������������{=�z����so�|�rJ`w��>7-m7\�w�����t��W�w��޼em��<��R�6[h_��|�>;�@ �(ӊo9���R!�)�g� &�ymj���{�Q-�a������':�ƽ��\�����){�9}��v��V[��7?�޼��z�e����Wָ��"�v��a���`Oh��6�k
0�(�r]!���(�1=n<k>2B�	Y��W��ךs�8n=u��]u�j ���f�e������>Ȳk�Y)�p��6$m]��禉��ɞ�o\o���GW�l���.�7�'�:?�ͦ��ٰ�%Tx�r0Ɇ��C/�qr��*� �8���	�E�	e>��}���概��$�r�]�1
���7%�Sl��U�=N�(r=KL�ϡ�QJ�0���?�+��&�#F�:�g�,���=ӄ5iX��A6|���/90 �W���y墇/i�� �Za�+
��f3,N�ң�y�s���O>��ʏ?^��3O��^�^?|���ޣ+s���5�����N��7�_;�x��^�l�	9����u�E��݅��b�i`kI�t�lvT�/������~��g���@0
�d.@���\UhE�B׏C�Ne,���s����T2���r�q�ʜH�P��o?��\����
R��}�'�/h�֮�2�U{���н�ط߻��;/�Ͽ�2�}�Ë�y�����l�r ���c?0�|���=�˱訥����r�C᜴�]`�",Ǡ�N���X����m���v��X�§^��������|�'��[��b��AAv���ag�ϥ�/�4ӆÜ�-v�Y���"�YU ���	`�]���rl`j��8V�~�D�����uu�vUg���'�5���S�.�����{�j}�2�{�y��μ���+_���O�t���+x�J�p���G�!bŌ�[
K^�����A��z�����z�/ߕ	(ɣ�$��(ykPD �Q#􌛹��}�y�G^}�5y}��xb_|mc�?���Z��2�����?ɼ�`��gގ�)����3�( �҆g��u��8���%[6�}2�Pc.�����	����=�k�Zu�>�iظq��*������/;�z�
���Ë�������{�g.���;^��}�Y�"� ,d���y�|+�;�@�4��kY�ć�F/
��$":ÿ	b�u?Q��a�����4�v}~mͽ����_x��?�;���g�񤻸|�~�9A7���?�&�#��z=�gY���kG7(>�zl��$V*@^7�0/q���	�p*� }g�u����k�R��Tu�߉{�=���*j=z��V��	 �G��kKaf��ve��_����e�ld.Nn�Dn*�3�E�44���R^�x~ȡ�=�qƭ7�c��eȺ{�oV�|d�������{��{�_y���x���o]�g�|a>3�G�7(L�7�����G@�� �E����͏����o|�/���o<�}����{oyeu��G�����j����"���*���k�x
#�2$p�ec�b(���J:^�zU W�����D���I<��)a��dab Z�k��e3��닶��&{�c�TԞn�$(|�e��r�RK�`&g� I ��֐C0%;�>v+ǃN�m��4 q�}	��ӧ뷼���{����������r� ��\���~CrzX�	%���&Xy��Ս�sl�?$�5@l({: ʺ�1h���҄�z��$������X7HuC������۬�ڑ:���E�~sO�]ëx��yۇ����Z����e׭ر	����'hѓ:��C}���m,c����]g���J�W�.���i�3'�7jѯ��S�_������7Ü� z`u���Gr��i���b7����k����_ys�ڛ �݃�͚��/�3A�^7���t�`|q����,wuF<4'�.�q�QR��'������� ���@��tJ<$#��=d輞��M=>���\߻�X߇~���W�um���O𝟰��߸��ozǽ0x���J��:�r�O�Vr�!@#�DB�1ȩZ'��y�7��Zh���2�M��#�$��у��:)�݀��<��>^a������WWW���_y�E\��\o��^tA�r;�M�0�7�y����av:�O#W(�V��b#ƛ�_���k�C�����A��ҽ�N��w�]� �A( �$8�3]���(4zg�D��~�a�}���Š:?�v���<�hw��_�<�ҫ.��� \� ���eV#����w���6�1��� �V�hER�%!g	������4Ic�h�Q��*�3:�GQ�U�����hl�y3��<��P�����ݑ�>ּJgH�C�<�$��RL����<�Օ����R9ypo //~��/��/_�/|�=��?��ů�����/���A,|fH�؄���P�NMAr��ˍ�w�~����y����}�_�����W�����=��x��U�__�ު��7t+�0Z9�����0xJ"�����f!ӫ����jM8�K���;�im+qD�E�I|Ӟ�G�u����G3h. f��Z^��o�[�t͎�騫����cϧ�����E������W?y�E�悄�f@]�l��>q=��.*@�}�˶ �������^�;$^`9ڥ
�UYM72
�����H��E�`�t�j^�3�����o���?^�ܮ� ����yc���� O��{��k*�
F{�='���gl#ǐ����:�ij���X�bۘ�S�+q!����~�������\�W�����_�z�����qԀ�\j�cj�A9֫���!Э��j;U�XW��������i�0��f(�G��\�@g�V� *��'g"���<�PØ����^��7��>��iA	a�2����{4a�A��0<��Ut�����b�Iq�jsTNG����R�c-{{%��~�Ɓ`�1�����8��/�M��Ǜ��{|��x�9��`���H�5��G��5b&������kE�oԹy0L\�#�:�X�!�STow���\A�
��K���l�lv^9���ol83 �Kg��bm�/���~�{cp�ȝ������R�Hۤ��\��e_+���'\O1_����/ƥ������.lP0����"�<ߌc�+A��Z>/�x�+����跰�+�Z,KR�T�k�����@��ύ���������~���j���kx���W}�������?��^���;/�_z��co���{+p�3�4�D�� 2^m�;޸6�������g^������?��O���|ӗ}�����7=\mp3��� X���7+�����S;���O2`�Tmב�]� -��3��,���V���i,p�iL{���y�-�fEa�(B�������d�V�"^�ť�����,�a��x2;t<$ٺ�v�{�+��zP���<����ݵ��²l{�.�>��� ��'�̥J�^�G%�,�d�cU-|	�#��i��
*�����Y�t�q�����Hnܮ�!�ӄ�j ��a������\9>�-a�g��J�-Y|v��@8�c������Y�ty��l�7�`Zs�]��O�a�4�
B$��d�u��ϧ�_��L�i�v@��%~b�{i~Є�؁ɺ�ul{҂zml��Z�3 !�����@���n�՛��ƫ���s�>ݘǛ�Ţ���������s��;��E/�d�7&�E_�Xu��e{�x��y�[�2���v�B���p�n�lssj�rƊaιM���4�0�.�M8�I�]&{646��]iX@9����65��(���i��n�r��`L}�ǆ|��2�1U�W`��ڱ���I����A�6��7Oܖ���w��כ����}�-(��$j[܄7q(��|&7 ���� ���&��s��:���Z��u��x��`�V�<�/���F(GS��b��L*J�Fj!�畩�YH�r�@�I�z�l��������Ý� ��e7��I\]|v�=��W�>��k�s}�ʿ�և���w��'����w�����U�qg36�D�� �t/~���k?��G��ӟ���_z}�߲�˟\=|��O/l�S�Ż~�w嬂d�" X�Y��t�©���V2�d�<}kaj����"}S���{��Ga5����{�Z,,�qh��6o��E����B�������ӝ�@3������xY���l�%i�:��ￔ��ҧݳ�a�����B�(/e d��3�Q,X#
��%��|L#�ud�ڃ�~�p�t.�.K���͓G��4��(J�!+��hX3�	���
��X�b���r�>4ǹ�������.8u��'p<׸�;��Y{`+ʏ _�,�į~E6E�׍/A�X�J��N��q+Zv3m&��x����xiো����U�E�ɇg���E�.!+
�XU�K�����ȭ�l�=y����.L̘��F���V݁�pջ3KO���ހ�w���tI�{;�V(ִ+�7�x���Pk�N�61mK:4�טè�HZQ���d���W �7��K��3�ѝf[
y����@k���Ms,����W}���
RI#ݿ���ekD�`$���ϋJ~5�ٱ�+Zj�m
�E�$V��[�������"ä�4�!f/fur�M�!��*N��z�v�>�������݃�����?�~�?���_��{O��_}������m�����������?�'������_������y��<w�`�t.�>��Z�B�� � <.���U���0���4W|^�w�����lŃ-��+�w���RWTq�VHmI��m��	��oA9���  ��"��ltX"�x$w��+N�,D$�p�u���V�&���4����٩�x�M�wy�ŝ��˦��d0(��]##B�aE�6�9:K�Ω�>��h/���&=�����RݒȎ\��WQ����M.#oqmH�)ʤT�mI��M�덪`T{S�5�Z���
�1�&�+�ޠoh�û�9�w5�0�����%*.���D�Ƣ��#I	m�Z�2Pu���hɻT���p=ٔБ���+:+2/z��(�D�o��z[�ye�#C��l��e�h�R��@��B�ɋ�����蓚F=�w��'_A��`�%��GKqQB�Z/��5wE��w���4v��꓏ᭅ��o�J�_���ksh��%���0�ܹ/y�FS����!i���.ɮ����p�ܴ���|V�w�4��\<�������߸������v_�o���w�����~�����v�^�ܣ����}�;�֧ͷ���w��/��O�
�n6��;8lV�!��F��ު����tS��װy�x��Ԙ��T� +K�td̯Ɲ# 1w���� �l�AHq=�sau�a% i!�A�E�5I@k��)�RI��u0k����#Ę H۵�t����۲� �,) �rKу���~"(�]%@&\�ʾ%�l��}��f	������ c�u�lǚϭu�1�7� ��-�*֋����*S!��WnTT9k�P�l�Q�,��UQ)���J �ѡ-��B�����,�s`��>�u�������l*�I�ԏ�U�7��i��s0q��]K^W=��Da�A9�^)2���#g|��lIa<�!� z�B�q5�শ�j���4q��r�� �adѥ�\��.Mإ�ݜ�&��p�-���B9a�q���,>5��iq'�:*�	�p��\m.��\K_Z�"s�[I6%{H�e")e0��[�g5��y���k�1�}'�<�0����ƽ��?�d��>�;�oﯟ|�Ϟ��Vn{��<����}��{���_{�^z�ަ����3��2}�"�c�)ti�s������x�M`� �Rf(�ܲm
�%���~k|���vӔt1ϣ�d�������>�W|�[�q�c�+[c6�%�p��v܊�7PgqS���X������R�m���,:W��?�pm����T#Ƞ ��-ѱla���0r��A'cl<[�?2���W[�]���8�i|��4���!(bp��]օ�!jQ:y��'��f¬eժ�G����}�#�W��b{AT%��Bg����MUq.��K�L��!PTCR|H��4�����
:L-�B��)�6g�V�#�*B�N�Q�NKJ�9?�xp�(���J��t��"���qzU�=�Xw��3���'��a ���#,�?r/�)����B�u��p�g�3ʸ��<�Lg>����`�T��M�^��K�}{!Я����#.��������\ͭN׾	��ȵ"���K{2ĳ�dv犍��jǸά�2� �X��{j�B�����?��|��5�CG� ]o6����}�����p��_|x���/�+(���m-�sE�B�������:�LNl�M/�t���l]QF��d��;��� M����C�eN������3y���,�R�����1��E��ӱ�XT@
u��àˋZ�Xp���C�uNj����H%83�b�f{�VT͹,z�p��P��hReph-Z�d6WG�l�YL(�I�Z��T�xx.7�3�-����q����T���:h��q~���Xw]<EeӐ Jr�$?��j�KP|��AXȭhXDۢ$	
$^�@� ���җ@e�����!�e-�Hwj�%`�:���<_��.�oFg��כ�]4v�1�L�v.V,��<O����o�5��K,L��-�E�y��x�л�����	)K0Q��7m{(�:3�4��'�c�[A�L���ତ�������f=��a�Ձ<F��ӡH�7|��C��c�Qv���j@�>���;����9sKtt
��e�������Ǿ�]?�z�-��淿qpa7���̪�0�Țk�����mx�yZP��p�dW�s鬝�>�l�lgR�����P��]�$,m��Q��~�x8�O�;�0hS�i�o��k�b���o[��?`��|Q��S���8�?�T1���t>�6�YfW[��f����uW@mw��t��:_���X&�w��}�0S�+o�v}�@>�O��mkװh�P>Q&kj���!��1��e`(�t�K�h!O�!OT�;yʐu�� t�PIo�Vǝ�#�e��rYrG�3��9]�a�Ԑ����ظNCDm�Я���	{��j�)�o��t�\�B�������|�>;�����:���n�o(9�N�9��[Q���� *�lȰ4�E��,���,ҏ��(׊q�K���3s�5��-x���Y��R��rl�Q���}/`71k�񈀥R��d�+O|�Fk�� ��.�o�V�'���Cw|��NAz��<�#��K�=��_����+3(G!��������Ɏ�����u�K�T)̙� /e�e )=#%k ��M�n��4��}��{��>l|ߞ�Z�. I�	`Կ_�"�9�	A���1�p7㶧P���\���~�qݣy� 	]4qW�ܭ�x?������7a�9��N�s�@��|�F��Ҙ�M��kb�s<�)��A�h�7�zB���|���� �?�wM��t��;e�-�+^z;ٺy7&[�-h�"��‼߹����y������zz�wY܄w�����;I~gR����[�!��t+�~���*�����٥̄hr#����μy~�̳���ݱQ���0��pl,�u�J=��j�h}������95ٕW������/�� )�Rc��0�5�-.ٲ>)���T�P���Nεv�j$a,���g�n��r���:�<�n��>i�?@�#>�hw�;O?�C �w��hp���^�tt
�k����#��\����j�>�{O��9bK����B`�g���J~��{�Ĺ�6��|ߥT��1E	<`�Ӿ�����喆�h�3P��-�
AUwض��^���%[:�i:L�$���j3Ȇ;Y����~Z0�ΊMgts�Q���>�m�8/}�"eWW�u��A��Q�s�A���Z�QVA,uEk�%0{ʱ�Q���~*�5�k�lÑ�#����<Ka����Ax�"�ֲ���V����5�0	�ģV�X.c�9�-a4���9�+qx�	E&�`@^c�|��ID��ј��N�$��t۪�&ymN��Hǌ����c ��F��u~��'�YWh��4�h��H���߭�������.�]��A�]4S`����dƘc�@�c���mQ񲣧r)�^��o�O\I��v�94���y�R:,�4Oָi���bv��Imu5FF�F���uݭ��Avv����;�"����(���W7��?}��?�=n�Lo/�}������M߉��K:?x��|�#�vA2Ic@eFc2�����c�����$�*�S~ۆd����W�e˕�VN�QU�T,�i`rd|kH���I}(˪���X���U��ؙf��f�ǣ�T�T:>z,_������F� �P���s������BYv)���,y�2)�Qe��)��20R�R*}f�ɧM�^d�Գzn쾼G+:����1��u���L�n�p)�)�R��5�M�.3X*3r���t��^os�)Y˞��3)�����p����83Zɮ+�F��a��Qّ��aMٗ(&Jil+�W�ށ���r��F�����bV�7F��v�L̾i�w�����cЪ�j�׬8���@oP�U���쭌���S��xzi��]����ҽБb]��^��N�P0،�W� .����30����;GeY�jw)\o��ۢ�1�_�V���D&��BT/T@Ƃ��:����2o��w����練:[`@4
۝n�bQ�,pl4��	򎣨bu���*�q�R�S�Z��o�8m�dlC���+�"�!�,�t�!����A�)�46ogy-�(�hqIa��M6��p3�S�'ʽ��1�R��L7�W���`ͪ��ɜ��!�+��2k,]O����=(�=*�������-G� ��N۵�p��r/�������I�(͓ �^�-T&-��$�>�ֶ�K��~�2QVk���}���g�u��p���e�)�zX��"� �!�,�WilT5���C1�hy�Lf���N._�6D��CM��N������n�A�:%��H���`C{RS&��kJ�|F���I!�5�ף|>�4*&��Z�_<���s-�\�F�>0�8�2�$��Ɔ-&�X��BIҟ�n�Wֲ0oo���g��=��[J����;�P����\h����3�p�i�ؚ�{�&��R������ �u�tC�$��4}�D����_�\>�4��D͊, ���C8G�-1�!p���9>��Mb�b�N)����;�Ft������W���n��NAr�w�rʽ�VCgmzZ�($ G�
}[[�幋r
���ƶ�K7����!��W9s&��^����I
���\UL0�8A��Kቦo|u���T-�-L?J(��l}[�+��*��V��f��]�C�n%M�f0�c#�^5f}���� 1�%l�B�7TD�j�E���S���q$Ĭnb~Vs#�E^�S�C4@,�g40��?�q�+(�ҚW���t��1�����u5h�iG�at��|w�r���貞�G���vηI�g\$�o�=͌˱�\y�OM��n<6��M+]g�iKi��$3>�F��(%�84�xjm�z�t|
��3�r�Hл�S>BC8�.�e��!�F�_�VE���띏��1s�kˏvqk�-�9�䘇	5���{� tX40K���M�[��H?���p��s�UB���G�s��)<��oU�Y/CG3AY�eZ�;0��[�@s�؄۶7A� � �ʢ(�Eb��[Y[��]�i}l)ژOc�~����������t`vE;�1�.ي�}չ���� ���vx�9�b�q٭h;�"4%[�F�2%g$�r[ �B���1x�o`��K�^tnV�����\[W�� r�Oq�;19Ϡ��W�5�a���#��H/{���̢�Zg�d	n�:Q�c,���!����BB���t!^�!��ݝ�&������5�\z�y�Q-]�7�`t�P2o-[���2b�9K77a��B�i���_�����Lm����{.�ı�f��Xü����GIy����̛5:d�!ky�6{����K����\͍L���?o�����M�P7�v��c�X�X��������k���v���G�[�%�HM����bޕ����Bbv�v��$WI�`���{G� s�������:��`�|�� \����=�T�F�6kE�v�r&�.��h��lY۟R�1q�(��`�B<��cIѭ��_X�te�0^e��a���׿mwfk#f�şJ�`�dJQ���vav������Z��H�D��Niup��}�e�Ǩ��r��?��i���T�,���d��X��s���R��X�R��� 놩0�@�|)rN�����t ������UF�B����&����:��	���O�~6���SG���iG�z�@�=l��*��y�B]ې�V
o�@g��9P�(���^�:W��N��i5��:^4dr3 �Qy=�)��a���H�T=�(����
�^>/����gEFN�v����9���H�A%w.�,�ۂYv*�mE�mZCޮ�*�N�@�؛����3�u����D����GnZ_t��^�=�t�
R�H�t�s�(���LJ庴�PE��Nyk/3�D�bq�-�p�tN$���ǎYD��u��)�G�R�Q�RT��@PPꇖ�F���C./c��JFL�@�F��<)G�@F� �yr�Jg��c�P�]B���E�Q����R�M��ac�i0��D���sX.�h�G�/?mP	TU^�ḿ_K�sԹ�����HvҲ�,�^��/+\T>F�1���w�����+af�[M<~����=;�QXRX1�x�QVר�R�(<3��_��q]J�͘&vtH�s
��k6^�m!�x�{��y���ql��,�=`�����~2f�/��.R�a�n��@��7�a�����軣S��	˚�D��̛R^��+S�i�jK}*+���9qn��¥ai3`�4��>Ƒ_��e����OњW-�����TY�ŚW;�����ނ4��rQ���D%����f`��Y���D)v��{��Ƃy��U���tvi��t`2l�J�T�TeEB�o�Cі��a�6rk�H�b5���Q�,�z$>���Mw����刣�I�������	!}a���p��銍��~HS�Z�j�15���U#�R��������-Ol�&6_E�-v�s�"�g˜2����G�@oQ��%*�r����ر*��5�;֙4�C��R���G��+ҫ<n�A�NA��wr�b1�p�����B����I@{[V�S'���T���y�.IC�4��g�b)����E*,�"K-���\U�y����2�R�	ϸC�5R;�)�0Z���_I؄a�+snB|�(�K�������%�2�)����@r)Z���]�v�AKP��]�s�=�(!+ہ"z�2����wQ��(�LTd��G��fc��?%e�4u[J=u)��9O%�_
w[�lܴJo3�K��b�s���HUڰ/�K�m�h�����Y��@���v(��и��G���1�ae�(d���k4�����I�Jc6ٴ]�}t=��\,�m>��ˣ�ٿP�e�$�Iǧ ���	D�P��hrd�0ALV�qV%�S�hܯ2%��tf,d�F�:$>J�H _,7J*«ѬW�2·\C<5�).�1�����4 9^���턗)^�X �j�lOe����3R
NLN�%��b��s�	(����3��������-�(S!���>oU�P󉍢e���܃P�WC~Z�lΣc?s��@�����T��ƀjA��3n]ʁ��R�/�#�P�RЏ��9��A%WH�dWv6؝w�66V��!�)���R�h��,��@A�OII��-H9hx����c��\9u�g�:F����0�H�ԛ/A֥Q1�t��ې̩CS촎��z����yɍOt�f+2
�<*�Sj<>�k5Y��qj��$zW[4�y����*H���ua�:�2���R��>�d��/�$N�����Dy	ێ�2�h]��>��x$�������K�x����|��T�]�d���;�s�� 1��WX&� ����L$��i�f`I	B�� ��VQ�.<#��r�>��2uI�I�(���a:,���.*Ɉ��hu3[�7l&o��g��Vh|�+�'��0��<��'�û��J�gc�b#Jm�϶���,I�)�x,`���uy�G�+W5����~艍�}�A� �mJ�!�XF�򳄫bTR��@g�R�b������߷�����;�;��A^�Ƒ�gbNv.����-�Ԧ��+����k)&���+�v�kk���Zѣ9�|�+���h��$ ����4�-�v�)	��M�K�K�c�G3�<�I�l������D����<47��ظvC#wa	O�2;^�����7HG� e�� �N��9�nK>P�\�k�BA|���y��mi4�$�J)�[k��
��\Ej�Z9wa�+�I��&�JũY[�� � �T��M�連8�ZU��ӎ��	��u�R9O�2�Ȭ�aw�\�t�"�9.�.�әB������1B졭��*�iI)"���&�PY�f����J.}@ꑰ* �L���[ӒLNM1���l����d����>�͡b$8����ʺ�]�r"�G	�<�JF�2/F:j�s�ϥ2�3g@檒,	�Ә��%>cr�~�j))��5ezS_3�3���US=[#��E��rz��s�J 1�WS5K��Y�t��n4�I>�cy,��sǧ�ݕ�藹V[�S��܃5����>k�H?FM�̀���p��.\�s ��#8y���C���/P==*�bЁƨ0eQQ\+�4�=�>��m*�9�L%��[��%��(�.5�����t�G����aJl|���1<1M����Ô/��f���;S����m��6o�p��x9kn��RA��$z�c���"i��q:K�����1ߘs���2�?7K��-�B�nQ���JU[M}��Z赶O?e,�u�����i�}1Ov�ib[��'��s���9�~Ǒ��8���~��b7$�*��t�fd^q���ze��U`{���L��GE�P`��tM�jǘZ�C�5���&�����hއe@��ژ3탠��&�'���R�O�n��G� a���aF1"�-b)I�1 j�i�rⱁ�Qp����3��B9.~A\P��|0�.4��^��mIۑ"ߗ�C1񅨑a�3s����׽�̨Ăv�Uυe�΄��$�00���LϨ��y�`*X�����}�Ƌۍ��aO-7�a�=TVal�O�y�$K�f[>6�J�/.�Iɴs׬<%=���KKw)w��b�p��0��!�����{�(��	6b��f��2�84-�i5i��]���h��o�Z����BT���	����*����u���$G(�$�Hjl�6���d X��*��2���m���9/����32x̭�T�2j���D�)
yn �qZ
P�*�䐌5�I�i8��EFڕA�O������������n��FMQ�����%����ÐT|x��M�*�dw�v�a���߸�oD�l�쎹��X�rr���ŻLS3.ډI�P�MؐA!r�fy�q���qq�Q*H<�a���5-ָ��N߁2�S�0�^w|������a��Ҿ��;{�K
A\�2m�p������֤."�V���) =���.8��p�K���	��r�x ��dkJ=��[?�eF����<�;�e9��E,W���3����3�NZ�Jp�E�+]ꖸ���Xh܌;�d�5	�L������I�O	;�%���w.�b��ϝiJ�k=V��d  ��;
9{)/h��x#˳�+Ub�Q��#7z�2ٮ���A4e)x�t�&�/���,+�i�E��}�=��Āgڍ�l[OY&�0X�b=t|�����3�&���_�E�t�m1C.�ĺ'�z>c�� ҁ1x�Ly�
��RA}�E@Ό�����3g�3�pK���>V�Q�f@�^�(6���*��z5�4͵�j�k�ޖ�VHj��#n2��[w��U�J��L1�2-�%%�]��/�-�i��R�9���P3�<�/rbf���\w�˞:�&ܚ?�D�;Fb刿�؅S\��K��Z|�9q�yk��ʰ�v��ug��L�X;��
��&>q�݃���|��Qf�&[l��[��T�-�>f��)�����h����v�l�3���I����0���>�t����?���g}g�٩	���h�7�Z�잩��o�p���AH���KB=�3�w������
K�H=+�;��E�i�Ԉ��
�mܨ�/:V�W)ٯ]�P��mb�ڡ��(W���"�=ˆ�e����3Hr�j���d� 0H���F\�Pnά_���,=L��Y�o�4�_�����g�^�v�P��@L<TRu��Q9�Z��"�7���i3=WmN0"u�T��6���$�t~_��%>��5�k�mV��±	.h��W҈'�[���6c�q�:D��D�.jc��<�;7��#Iց�r(��7��4z2x�r��n�']s��И1bv��P��e����Hr`��p���/�����ug�4�oC �h����JH}b��qlH�j���cO�f	(�y���}�X�/qi���1�]�w��#&���#�%
�ڑH^`�QM7���8ֳ��m��]��*�� ��|.7�l�{0�cW�I��ʐ�)�b�公9��*G���Q�qe��=�����G� 9ʴ�]�K�q��ʴ�3%[Zќ�AI:
��e�b��K��*E���]�3G�c�N�]6ܞQ��J/]���T��:G���D#�U�*������9y�F��P\ G.ô�Y^cE!v����Ё�eS��2����߾Fa?�r �It%��/�8����{�z'����N|N���U��x����_�̉�9ۭ�5Ғ�Ȕ��@]E%�2*c�15Ն�܃��ͻZ�
_B�h�(�,�C������*HѺҺ7F2�]�xδ�_i�s�Lv�R#?n��ʄ��g�w�,���F̀�c����x�j���v{���i��}aݲ]�0�o%/���c��g����F�{]j �S[
%-��j�-~	Ǜ=cc�2-�P�L��-�)��)����KrLvM{��%��u�K�z���L��/������������&o�`C�E9�#�'ǫ �C�r��ֶ��a0�F&e�-n�=�֏:i��S�#��;Z4����90��/��4K������-T�w�����L^=��p#��n;Ky��+[�Zs[�Y_5o�����"�̢kE"�[�c2w%7P�HKvI��z���HfUQ��"l�2"��?���b,ٺ�ET��T亣$����a�O��� �q>�
�ǁ��bA���Oi����f��=��t�-�r���=0%��p���w�R��/�
�ӎ&)���#��A�Ö� d��<�����g�g����,#Xj����-��;y$`������T%���L����ŧu?�q!� ��kFɴ��@N�3���p
jw��eS�u����U��R�FTΞk/�uO2����\,.׿�	b3^����v�$�* @+��_E�Fe0�c_�!��)-P�[g�刬0��x?O�1������j_�2���̥~3/Y�ZQ���h���9NR6����g��t�������(��;N0i;}6Ϩa)�b��"��K�2'�a�p�����uI&3��I�X*���1���|�T�奉y��&���%�}:Z��Чd�+�����Z 5���"���eC����~��w�.�ғ[�+|а"6�%h�	g��=d�9Q*�[i(�ևp��@�c)
2:W���N���N��" �ŌU�ߝ��#>�)5O�#��=?��>���jR=�H�N1����/	���4�S['�zN�X7,[Y�2����r������V�L�]~n�ZD%;�AGG��ғO�?�oqs
�2ް&�#����x�Xåѹ+1����˰���L"O�YX*;���ǔȃ��5�EG� �h,:I��'X2��/$}�f�y+�����.�@c��SlWS�X��U�,�C�bay�R�P/��`泾$}y�����#F�4"��R���ڶv�]��oN^H&4��E����mĸ�6��f�?�Hc�5�-c�}��m�MB����.S-\�yu�dוx$���v+')��u*]�vʫ!#��ӣ��m�Z�?�l蚠A5�뽻{]���6X��g�`����Q���Z$�$�`��2��M
���p\w{2�h$,�/aV�~� �x\j�3ϯ��l<����t���,��^[�p&ײRA}��t{I��ɍԞ�wM�-���h"�mC�\�Q�Χ8Oz��ʤ�*/��W��N,~sv�Fl��i)�~�ݞK�)�9���'M��Z���������_��8��l����@*�%^�Sv����qN2�?�3|F(b�Y2��-HU�m!B���C����ڧ\�X���Ȩ�ؐ0Rm#`t�\f�AE��Xn�
���$cT6��k�w����l"eU~^��]h�~�-_��亿p8��0Ad����lT����[RtO������������|�xT�m���p�-)*�b?b5���_2���H���<v�@;�i������YDc�Ai�th��b�2BA���$��3JZ�%$�/�v,��v�P��9�h<9� ���)>!x��PEG� � 0K�^��k�@�4&��Gh��)�s�����:L��u�U�儉��(y�}���W\��I��۲��י��L�G!�	�(nT���b�^f���.��}_7��?�ב�?F?
�OJ���!�bl.v�Z�e_`*)�ܴ���T�@��wK��)�p���H�<:p��e=1��@s����Ӟ�d���;����>NH��Љk%8��Mq��^:��w�����:�
�K��a4���CL�r(�i|� �0nhN�H��0�9��Pn���xP�Lq�ZF�K�R@�'+άB���ʁ`����%��2��� ��N���ǑC/���(R9di�a��q�r�@&9c�	��u1<���h� l���T�Ee�蠞.?���8�N�ҵMSRo�˥�����Aв�k�k]v����;C���3l�^Q�󅓗�3H
�d�d[[��e'L��U+Lb�.l����AVw���`TϚ������v�6d���C�e����8Sl��hrה���X����J*#w��CN�(�ߴ��R�oE/�B6~7Y{����XJ��<����(�l����7�ؤC�l�;&� ���IL��g�I0}[�����l��%�,���1\.��'��CSm0�6姰RgUp�$�P�K9�����QӦ����B:���d��˖���/UZ�4��Q
*;As�B빱���7}NZ�X2�H����M�L[�1Tz��f]�[ȝ��4���h��fYl\B��QN�w�Ei�i�a���Z�z��D���LL7�Bp���17( M
H�Zִ�UZw��v�K/W�˳�3mO��I �L;�y,�j�A��4�׋��Ӊ�\����2�u����!��F=pO�Y)zg]z��g㫮v�\Y����wd�B�\��Sq�� ���~�$M�Vg���<77�C�>.!5�p�+Y���+�j?�Ѝ����w��U�\��R��	���[�1�{����*�- 
�;{��R���ܴ�QK�̶�av���Y�F�u�f�.*u4�	����Y��A��U-�c����T<$�ֲ�35�6�k�t��"go���w��x7@[!.�BC[zN�vA�;��/3����9���a��Kν�1�V�lE��weU��9��.�2fG� 1c��ص+{�J��������"�Yn�:���H�mr�YP�P�d>�/����!N[��ߦ1e:i5����]��Ol�ofp�%T
iP�jO��;�ߒ��@�~��;�ޛ���[ Ʊ���-�3���(�0�V���h�WGL6rFf^>�;N�C��r��~W���\N`N���nj�w��-h_G��c�G<�e����tq�WߣU�� @��R�;(Ch�Ց��� TF*��u4Z>�P0�ܰ��v�r��La�)��vB¥�Oj����g5S��z�.V��H��Q��6��ӲxQy[� i��A��ہg�v��Y ���:X=�&TB���5�*Tڃ@e��btV�r*w���
����~'X�s��i�=ӁIt��S~��g`'�g9������9��]}�#�ϰR���f)s!�Et�j��I����R���� �F��8�o�q[��T��ۜ�R
ȡ��4�4{�Qۻg�7n��RA�ɬ]C���vY�(�K�� i�@�^�ߗu����V��4LE�2����tZ6�,Q�^#r��	�v	��Weaⵌ?�J�5i����Kb�b�ĩs�,�]W��ATZ�0D��A�b�S�++H������d�� F3���p�́���޽�㳬,�>��=�0����nʕ�m�q/��z˄J]�43'�D�g)J��bGX�C4ۍ	����Ux���8�Z
�0��xGJ�^s�+<0k�$��X�ʎ�T`�����H�v������!�ύ�n}W�c�Z
d�\��e�5�!�
,��W|�#Zi�t�m�LG� �Q��
`�6Z'[L0���4F���r3���$;��3%��.~BZa����Lh�n�)��W	 b��n*Jz��uD@h�C���XfD?�2�[I��g��B+�V�%�p����.+���w扛�r-�w�s��ș�{�D���31�i���P	BuC�}+�m7�v9�Ρ�B��9��*k5G�r�'��Z��`�L�W)�
�N� *�9!jWE���t�ڐB'� ��
�Y-��x�ځ�zd�Ϟ�9'�����$��
f��GQ$��$�I�`��kq�hFvR������џ6�BY���0Me���:�+_IG6OϴwZ��b�;?9�0�\����R)��w��7�1�h�s�\r�,)�R�_���$(>%�s=�� bH�鈵fDDFov"r�o*$��+�7�SS�p�BP4�S �!�,�n[�n��,���V�F�2�����`�j�i��Q�֘˜�����8� /�T(���D��TT�N��iO�Y�[�5���[��Ю��Yr�dH��c�(�V�J�F�-����ʠ��M���c�2#��Z�]���94���To��8���@~E'Gip�UJ��l��O��;=~�hu��䷋Q����%{���aw�I�-p�h�`�Zg�2P�k��B�F�M�u��:�w��:�wV�N/���M�3�Ul�[�Y�2&{�[��8��	)H�I�����_�rTۚʀ��
�Hj�AL�H��۠f�8�m?���Z%�?{����/��c5�иp�[�]<��v0{����&9����S\L��x��BZ���I�Q'Tm�|��npL���g�w'+c��@Kʵhߌ�,�M�\=Ҿ�c*�2��Q�Ѱ��o~��9tȱu�	�ݖ|��y����O��M����RY��W�0Fl�c�j��ˣ�X�(��5L�|u
dKW����w�h�R��x��Ak��:^ u
d}�{˭�� װ��h�K��E�3�IX�U�k�0i��YRڛ�&��3�Vϔ�*���$Y�kf�K>�;6��V5�� :RX����j5�����&i�d�I?�+�|���{F�!k��PNp��m�ww��g������P�)��A�9@�Z<��IWίmkm�Ӽ(���3�L7p=���{#�F6���l��^���8�7��<&�/?W �b*W�:0@z�N�����ԌOigo�`y�ۊ�2:�ls��uT������E��܂9R�@���e�W���i�<Ӵiy�+�XѢ4Y ��ǩ �~C^�e1��Eki�
pL�T^$�0�.m�6��
T^�)�(��*/hF!�L��r��0�l�e�@hi�1E!Y\�Bޤ��}�1������w5�{@��m��P#�!������؎<���+x&�Uۍ��Sz�j7�1Ӻ����Hw����c�ؗd,�T�Ko�&�bY���GQ#�� �S�L�㷕j.���00f�����[�wUN�%!W���"!��;���� ��F�ZGU�EB������f0��X{w0�x�.K��q.�U�d]I��R���Ch�k�ƳC�|7P�I�c� �����b�*/)+n�{�vgV�dE$=� 4�X�(�ߞ�k���4B�w ���	��j㖾� ���ɉ~�#8���v����Q�WRQ�d�����w-��c�ڙ���9v���s-Z��]�3���	J&�L`���?i<* o17���Qz԰,�W
v2�Fà�D�V��c}�g2���(���ZY���V�������e$�[�]{��f��(H�-Cڳ��&��$a�S'�9)E�-=���ΧԦI��{fw��P�qwW��i
@�qLl���5S�/�eCWe�v���WN|�-��JwՕN�h'j��2��K�f�*(�$�=-2"����d��[Ќ�z���cǞ��\9d�D���ZI#?4���v�;=ƌ��i
�|6��:�ȗʖϴ�d<�c�y�{�-g(Ij?C�75.�y��ػ���.�;��e�B΃��±��>z�w��w"d���T�y=q'�Q�u(TцR4��\
�{}��!n
멇H�^Fޘc>��jG9l!k�	nQ���_���ϞQs�ͶР��?�}��?�3�sV�N��ؕ�*T�Z�?v4P(�
�DU���[������#S��pWi~D��g���e�`���g���k��<^++hX����4S�NS���aF��� k'l����a���U�$/�ٝJK�k��1�"_�h��wOv�c�G� 1��[�|2��hL#7���J��4�A|7�ѭ���Ę�D;�5���֓��V�Ԋ�a���.+G�EN�ݦ�&^��i�c����p-M  ��UR@֔�վk鎱��M�p�4�)w`��ʛ����"1������=V^8�E�S6��$�Z��FQ:�׊���Qq�Le�A��FM�W��yOo�Wj�����ㄌ9���%��N���u�1�!+�x�d$^�NO���P�LgZJa�C선����&(�|��O�셰y�����v0�H���	��H��!�Ӑ �7d`�p}e���-�w��2ZA�G�w�c�6��V;��k��mik%�� �@|�Ah�5����S�KIŮIDJewˁj*G�L�F��cc�a�ޅZ�ޝ���zU�A�~�CR�lY������-���v�%'� Շ���@3�� 0(��v�����|��]��
E�tЊ�ŽV��B�t�?BӅ�c21;Ch&]�w���p�O��ҹ )�������t�cؖ-����B�p���ז��@e�l�"�,O��K��2L��~�;��4C�rqI=�~�B#���0��C�2^i�i"u�M?����-"Ѧ��	fv�;o�`���5b>�@l�AvѼ��en�WE�q17fZ��������/m�0�4M.����ѿ�w&��N�{t��yG��!E"4d�(�HX�,/��,Wȭ�Ȋ)x#{~,Z�a�d���s�m/��y�Y��gڕ8\k����r�>�x�����$}/� ���(+�І�|�����k�M�o-�3VԜ��-��Ә�w�r5L��
y�H-�{�3�"����A�ع�a�!��ZO3~�jZ��Ү��(HA�����T�1yHj�fog�rz۱��������r@�3x�����g��yO�B (J�H��!���E�'TߒW���F�
�����wO�r+h3�i�f�"��Լo�o_T�KZ���yMg<v��O	8���;׾?P܅�u(Ɩ����c��X�f'z&���i�<�ޗDk$&K�����;���n�NFA���HK�¡t�[�Zy�L�A%(5�C�,��ԈձF.�aX�|H��	r�?���ES�"��k�����H����=0���2�tvyA��k�ٮG���Fy�A��w�۠�T�
o<�t�|_I�)v�Ogw��ݒ&#TȠ�%R.[g:=��#H��<T�X�t�rd����ɾ��pVn�m� ���ŗQIK@������]�.S6o�D�����k.u�L��F��s��>�#���y�Ҳ��.#'N���.��JV�]��PLg��A	wT�'<5��Y]{A�P�I �A% dV���U�QO�\K�ry�*�Mj$B����ѿ�Ux:s[t2
R���Ha�̭���:ә� W�#o"��JV�}��2�oD�0'��H����"�b�.P�x�<{������h�v����~q� )� ��_�L�fj7�:slJ��Z����l�p!ص�"�U�ep������4	����L�V
ϰa2����oB�����{���͜t�M�2�̙N�t��Mk�1g��=:z)m+�V.*U���X�qX�~~����x]���,y�ۙn���Q _Ӹ.�D��K2b��x� �����ZK�f�8���3��h��~��c��[�3
��;��u;|Z�[[�y�n�=**e
�B#m��F|��}�1r�jp�
������}�[���Z��b�r��[�W��u�p/A�| i �����R�����ǉ�Jna��R�p�]��6���]'��ed��b��>}O*�x�3�Zpıt�I�6H��z�Â"/3Ð�])���Oi��D�8����xG4��>c�CZ�u�b7�@|�r=�#��ܐ�mxe�o�>W�������S����e�N7Q)V��G>��lQ5�q���s#Gx�)kL!����e6f;L^���7M���V�Ye�h/�lJd
�*�Ϯ���ֳ@SKx5�Ǐ 5W���h��ƹ����-
%fQ�~��L�G�B�<��"��r��3)����m^�-M)9�߹58]�K|Ɔ��@���T��-@�k�=v�x�	�0{ߚq
p=�ֶx�|�)��R�"���9�a�,,���P�e���rd�t�M��6ׁ�⟱(@ba]��~X_���	�QN5��m5���TL���UtU\I���J(�N=pDfp#�h� �Y�D��j9���6�$Ŕ�r�<���m�;n��g���N�0��j]C�E���LIl��t[��EJE�����i*H
e���� ���0J�6����h��C�Ho�gn/ږi����^G�f�'���H��'l
��w�Ф��.���͌���H3�6�l�\^8.���&V�S��l��i��Yt��徙���K��Hr�_¶��+�ؔ�&rWjv<��vk�]{�;r�gJ3��EP~�����g�9����4s}�6������(H��F��A�p����❙�"	0���[
�����>�]l0�E���q�UL\�2�O��񭱾�E���ƙ�x��q�.��c����t}R22)!��K&��Ѭ����������ׁ�>@((�{W(4�o-�Yϡ��0�U���`��s�t�Ji]��K�S
B��4�`�\�)є�nuH�}G��y1����#a��� �'�I���g&��/����Ƙ���>��U;E4��ְH��H٦�����z�p��C��1���S�g�<X��ϴ;���[��"ͱt�}�]�1�p�*�{jh~��1�XQV������<3�,R[�$Sg��� �Gb�,9IF�K�T��PQj�Ť>H��"�a���;�5��nbr�R����5_߸Q���Orklz�)����>�;ʨk�4�K�ȌLʪ�%-PT�4�ǭ�}���S'$�	������WH�y���j�����)eg���x(�,�~�~��([VZb�� s�A�<3=�؏���3�9���+E�(^��mfQ��@r�[Lk)p�1$�sV�n���K��#�N7����׹s��bP�0hHX(�eY@����k?<.H�P[;��BK 1���R ��9?���3���B�5R#+y��U�2�5�0��=@r��&F<4��/�T� �+)� ���|�{H/�}�E�\=&
2�D7�)��|��	Wzχa�Fv*��b���������@˲�y5J��({<%d,UG ���Hʄ|t�8��?j��p���e��K�Vݤ���Q���~Ʋ�-�4�৹ׅ�qA�!/|����!$��}y�$�M?㙹�++Z�]V��N'�(?���tZT(B{6�Cl�R�Sb�x�Ŀ�C����)���9����)��VěY4��	���t;�G��p��'�Hf��eu�MBqrV7H�5-`�=�_���ErdUnV�\�p�ŵ�3!�&���Z(z@��h �.��-i}K����bx1����0W�Cc��دJ��a_Vy��Es�ȜUz��p蝑�03�ǫ�]}M��C��)GE5���VY]��T�cR��-�"U�X���֏#�m_���Y����T!���| �o��?�o��&vP������O7��\�I�����t�$'4.w㔜���P>c�vs�t�$�:���{�0Y��'���!��:�g���)�m�}H���|� �N�R	+�l�"*,�&)N )lU��|7��n�]۟���d����[�r�&�
46>( ��#�� `��h�$B-��J.a��dJ�R���")��K��k�&�(S��d���W���>)S7G-���H�)��vx���,��d썯0�+ܮ"�$��w��^���G�-�(7���v��>��}�e��#�"L
b�\�3�Z	�nO�g8�֕M}�\O�tR���Q�hw��X��_���������m�w�1�0��箰 ���א�1o��f�w��҂9A��v��`��!V��{�k
���`�UՄ
p��Q����x>
gM�0��s���w7q�ة9�WWu��=�$^>����<�%g��s�E��=�Y'�����>x��mf�8qϵ�CS��ź�r�w��X��H[�\�G��|#��,ƀʎ<8f[��Uc
e��j3�ڃ�O�1>s��0 � ��yP��{R�ZdQ�tLԁ.g�sf>�N����h�$����|�MI�S�X|�X:R�:�U���L��r��aM�������ʷ|���)s�t�
��|�����>���ÿ������^}t���ۍ�����R.2�����s.qR�N~ۘ,�������2���d>�w�FG�a	��>�\D|N���_M���y	À��@ �^	�"Wͦ�B���p��Y��L>W�Ń�4�
�rXۃ���v��eO�x�<p� Wq[��VE-���Õ,-�,���o��s�K:;�Ԛ>a<G�!����OE��.���E��R�����EM�7� >�����`�)��� �9l�v{�M�x��k�)#yV.;��t�.��e���<c^�C��޶<HM�̚�塎'�8.��R$�@t�.� 6��f��Vʡ�8E�	�j!�Y��{�T(1a�ج�-W�Ulv@��@�\:��;|������+M>r=CE����l��Kјl���s�(��3�]*��8K�2�.���������w?���~��|���?�����?�U��́���/���?�ӿ�����ٟ��_�Է��*z��J�ʲ���m���GN�§Br<G-�(x� o�R!1�x�ka��?a�@C�=��S���C�B ��hW�H��`8k��G�@0�L��V��!I�~'��fH��A[3!x��� ��v~�nc���,����mHsݤyk3�V�b�� �v�<֔!���DN�� ��j�P��c>�[�²���c��*R�(� �!=!��M)�LeY��-)v�X!�$�7&DN����}䀔��� ���W�a��Ҷh3󘅼N�R&�H�4��p���{�<�X�y{��Һ>
�xB�,�,�+�`MV�b�h0���rș�	O)$�_2-tT��/N���|��<_�,c�P]�iĆ�y-��01d�ɵ&(z����G�L�N/)�,TړrT
���7>�M������~�;���[�����o������֏�Ѝ)H�������~�}�������%^Ɠ@)�#����#�S��2���a�4he �|n�!��Q	�q���l(��_�����q%-{�_�D�t��c� �Ͳp��[/%�>���xq�.S�|���h��`u�3ȼ�</��������+�]X��G��11�6�\�:�w�<9K4���$ ��u�$_6����X��,+l��V*1���(�z%�3Q(R�}נ�����j�,}&���hP�6�e�/xC�2�k�>U�BS;�ؼ"{0����4q�o3 m��� �!���*U�izsD,�<�CɼQ�ч�β���m��3�l��D��֡a��x���1�Ƶ���MHm�o����`♷�48Ȣ�6�xi�3�S����Q�pX��O�����_p��ؿ����{�Է~��}�K���2� }�����?�޿����bn�*�X�����r��,K��Ng:8�"�Cj�����RZdAO��b\�y��H�� ��n�n;�#�O ��%<4V�.���+��5�IcWC>��.��*x��"�gcB�H=�s�l6��_�b�ڬc2<�&e-��0��-xkLY��)�L#Tk�i�{YR����pd7hL��KְOȑH�m��'�� ����F��|{���9rR�����r�vScz�V|��/�)�t��~��#%w��Z�b ��ۧѢ�-V<"t:�[g9"�tڰC��NL.u�k1Y,"r ,�F^�ɪ�zg��
��"������	�)�PĽ�傛j�mL<� �T��(��qqd�c�.Ƚ�c�y�P"*��	�HA��l�=��-!�����o���߷�W���g��{���/��>�=������������?��?���Piٸ�AT��2�Cq+nW�]�J%?T`V\��+��3h_k*h(��'+.�B��p(�ou�݁��3�v@������F�\�7�	��MPR�=�,��L�sDZH�p��n�f�h��{�< ��d�XR��*�uȋN���7�HcJT�T(��y�� I�8�O<D �$�	�A1v��y0���L�0�X�#����nU�{J�(�[��+��2����xCL�a���)�6�xB?����1[T��IT"r^�&�y9�������S�%���P5 �jfgUDF�au1|����ABuI��4:$��w�E7����N	i��FӉ��b(.p�Ğ
�S"
���H� ��Z]8���b�֌�]���������[E�+bL�}Y:Ox�gZDb�;FE�'~�c������~����������Ϳ�K~Q���?����/~�O~����%sD$#��O���R��bw"� K��o��dׇ���Э�~��i�����4���@�s���J�a�n��Z| �g�Bʦ���P�_�ާT��0&�
V	}���8��,�i:�C���?�7 ��O甂@��d�8���ɕ��8�X�Fט"?M�T�c +ˍ`�1HCٮ"c�t��#����� ��fm�Yu�_r�r o���6���
a�!�N�)Z�!���M�E�b�	:LξXR	����<���64���g��g��ղ	T����l�G���ґ���0�t���6Oh����ܻ4�7?7�xb�z��neLi�q�m�AэK�Ue�J��ZUN�?��(TM6�ߖ<�i��9~���Ar�u'�l2*�Be�b�v*�	/�}pi��Et���R7�Xَ�����I���3����`y{�����ȟ���7�������_�s��ὋG��W铟{�˿������>��o4GK�խ<���~?�t?9�1�Q���Ł�ά�h���5t-������I��Q,���<�#.�g�7����t��A\�`��3*����@��ȿ�~���˞�>����Jws�p��y����J� mF�8�w����ͦ�C��RY�����F9�\=��Q�l*��v�"Ŷd�&?�F0<��*w���~���s+]�+�T��AQ�=��7(ޗ����!�_<(_�J}R�M�t��N���0]�PɅ,�u�]q�\^��;�Y��:��aGs=�E^Ȃp�c���u�V�����k4�K7�h��� EkcX�OJK0p��"v�C�]�xǭ�(w���N��k��%DI���)��U~s���z�7�Jc�t�&�+����zs�����|���������?�Mxχ��7���������ѿ���̑C�M�'੕$�����.v�Nq����k`a[&I�P�~B��m~/�����K�&�}�,(��x����,YO�>f�S�O��x��z�I�)C�Vi�����p�`^1��t�#w��C��",��������~��X�j�NE�U�Ӕ<����%Q�H<7r�*R?���.��Ɵwp�+AbP�'P�,�����l�{��v['��9h�<PĺV�AV�Y��z$�[t�S�0�k=�8��	�]�𼥉\�B���������o` L�YZ� 1j1\���Af=�C�����&��[ׇV�d5��/ɑ���Sծ֜�v�CF�2��s4�)��fC�Iօ#�+�T�%U8�Gg}�Ei �;�����G�f�9SK>ӳL�R�����~��w��������?�m�͟���<����~��_~����9����o��V�Su��F�btK��sg�An�;��D�L��ur���ߺb6����;7��:E��:���0;���46k����"��p���� �w=&����4���>�_^(ۑR ��P��?**�~esF�$,xl�;-cfu2�Ԇ�nRԩ7��^�,GlÞK�DK�O�r��8Rc�;r/����(�''k��`�jQ(���'��<f珵��0)�>�|��r�ԚK�qӘT�2�����u�S �~�@ �ۇg3�1e�}���gɦύ%���p�1���FY#u��)���Z#~'W�Pa��5�ϖ�k�MփYy���&La��h���*��3���g�커���_�;?��~������_|���7�e�3;)H��^?�������5֞e����v���XĊ�D����x#�D&�����H�H|"�H�b	��R>�$�qDl�K� ��cl@N�L�#�bl��o��>�={�=�]�U�Տ�5�����;��Z3=�=���U���������;D�Zt�B/����ZHj?�ܨ7��y4|�n�]A��|���fAR}���tSsҕ+���?]'�r4�\����E�.~S
�k���5�la}-� 3 ��Q�0���ߣ�s�R��Ygȕ����m��0څ�wICB�����{����
A"A��F����s�*�[,�`N3~9��9o�p��0�*e�J�R���)�Ƀ�C�K���c����^C�QDq�R���g�Lҁ���g8s�pa-,�q`�G��?��������_��?��_����T+�j�g?��_�O���_������N�[V��#0�Gx1�������s�r��J�ŢV:r=����7%�D�ϒQߨE(��t��\BR�0E����[|��d
�`G�C��J������$��۷��	%��:Rv�&!%�+��,��]}XWiD+;Գ&�ϿkTO�k�K̀<�&�h��`�g�![ ����V�x/RP���s��C)�P�z�'��������O��Rװq#�,Ek��`\+c9M����^���f�?-�7Ooo��am����ѹP�*D�������S]bʅ��9�"����/���_�c��w����[��W)H��F���O������IP;�:Z�:�)�p�P�Q�fs���\���Kn���-b��Kd�OI� ��dI��';����R��a�}���'��T�� C�@�UdK��-=QRMz颦h�o}�?�Y�s�8FAC������_��]��e(\wn����bUu ��DB%ǤV�j�O4*��6T�/�\�Wb}�bD���/ܧߚ�s�Y`��1�[B����K��_���Z�5n���c�D�P#šQ]2��}g�1̿����#�(bQ9嵭���k��i!�qC������_�¯��������/����[����d)�b�����������O��w;�+vL[����b�i�`%�N1�p`l��K��dZ�d��[l<����h	�ɽ�D9fw,�f�D�Q����$�8�M�Y�I儚��$��Z���
'�۽�����ncl��|��f$E$J?o�/���4�ߖ�t�_w�O��$�q�o0DvtAQ�u� ���\�Lڸ]|�4�]��ӵ|Ša�sx]u{�N�����9�Q���"�ݓvD�j����*k ,=�	�y9+x�*�8�vu�x�4�|��Ԯ®3}�nf��b�:���Ub����l(��_����=d}�)��?�o}����������������,R�~�>�7}�7}�_��rdO�7��D�,�kV���yiH��#��<��
�LqF7�L�׹̯���'M�-�ϊ�g��FR�*@��Q���� !�`�[���0o`w��דB��.�E�.DR�c�(��GH[;�6�zY�L���E��3�*��X�JyY�x�R�+�%"6�c"�D�kj)��$��#fkխvHq-{Pj�| k3V�S�柳V�g0Wy����q��ߋ+@V��f��$|[�>��b�Ɛ��YEM�?87�ٟ�����HCҵ�/�O�7Л��.<�� 7��Z�R��������O~�����������F��V�~�_�U��M��������tw�g���E�S�B�����JG�ȺعrdW�]8(��v��;�����B��>R%�&���gY49K	����hpz�����]�3�������y�,YY��{z�)!�C~Ϯ�L��!��-����In��@��E�"�T*��TA ,�S^A�\�z�r9q���}4�,r���K�~���#��F�Z�d�|4|�l�,Qg���4��/�vfa�9��ff�����b��Н�0���:�m���?��&�	���@2X�c�8A.0R�2�Q��M���(L�13^��r$&��gY=�8�l�k���T�;��?��'������������n��C��_�������-%�#uB`>I��,W�A�m���8y��,^�4	���W�^ ��^0+K�������\��8��R7��bsD�	4�Z���4>����_aC��U����iif���*8V�*Q�5[�Rn����{�u���k!�T�t��ҋr�.E
�E
�A��^��Sy�&(M����h{�F)G����)]L�� 2�}=[\P>���K;X��N�[����=H���4���a�ǃ�=���Q�~���T�k�N�DjG��NTe�F�"�M;�Y5������Ky:�-%��-�����zq�����o��?�_~���o��_�#t�KA��������ۏ���T�����M"]�C!�H4n��S�eB�p-���[0�������X�IA��������O����i3�JGqEZK��w�)Ո��1�:U ���'8�n�N�'�@*Y� �y�Nk:J�sk��<~e�Y�.=���u!�27s?�����:��p�w%�H��cR�[�V���]x�o��^f~!'��X��upp� S�g>�ѯ�]������|�����T���_���~���ov1�e�_� �EEi���Z�����|Ɋ�v7��N]���\��PR���fע��b_��<�����ֲ�P��AY���胳�^݈FV����������R�Tq%��`��s�=�u��P�U�0��h��(_����={ɼ@�#��ZE-e�V�&
�.Zӝ��5�V�L���wE,�:�JF{R)�"S>�s\ٌ�hN/]����/TUV��
�W�si�]8�w�I:�#�[�����C$>~�G����}�_�����o�~W�_��G_��~��|�{ �L~��]�82�ЭÖ�7�*�&.0t�Ko�*=%���1P��_GA�,l��F���$|�t-Ʌ!�LPN���U�v�\~��h#�Z[oA�Qn��)I�q_k Ə�A�J���R�s��,^c�7�ML�4��L[��u�Oe�����v���k�=Q�Ղ ������%`u^��$���9r�8�����) �2!�I��};�{�2zˍ,ݘ;kZ�����)�P$��'}���j��Q�Km>`}�b�#���������|՟�{~���
ҿ���o������� �[6b�ohx�e�,y����\��.:O;$+�=X	�R/iZ
I�
���U�˦7:��6l�ԍ�ja��rf���킵������dFsO��<N���RʰD�M��؅4��j̟c�aB9�4RBh�Z��6��\��tk�)�Ma<ҥfp���}�VXʿ��[��.Y׳q�*��<ϔ�ptve��s��[B�v�{bk0�(�>�N���b'�����w����?�{��� �O�����c���{�%Ț�N�|���i��rJPPn%]l� /	��ƽ�U�`S�f9�S�)�h�jі�V)e��KF�v���p���������E�/f�+���|��Q�m�A����E��k��Es%Z�𡐏�_�[IJWAe��h|K ��x�8:,�xw&p�dA��UW.w����Iq=���W/�"�(�Zz<ϋ�KfH~,�_����!|F1�86V�t.���+���Skm漉��<?�w!T�� d�����k+U��&��_�D�낒:F,�&���5V`�i&e�`ܺp.��t%뙾G�L|u��`ί�@�������[�����E�_���u��CJ�׭��%�K�3r+��>��@d�,���-\�Z<jN���e[������U/v��ٞG��)	%�	��sV>��0�����b��F/rqD���b[`;Z����cط�*�۪G�ii�b5�3�4!Ž z�Hm�B2s\"�u�x	ۍc.�s]hP��
P�w-s	���|��QX+\y���  ���!�, ����J߹
ŕ(:H��6�Ҕ��ЯdE e-����hg�����۾����T����������t��U#;�m���)D-����D�������t��`7�m�����Xw@}�ʆ�1���KԨr� �0{��{�c��kjݚ�����o�\U +յC7�ϯlR�6e5A���oR<�歀ի=�\���,�#4���G~�'�+��$�sez�xL�l��v}���o,�4�u^2J�$��6_��*\��6gd3��i�I)Oz3ۅM�PL�����W��A�;�ʄ��!I�o��ŹK1:0�����TQ&�CRO���Ե?-�*A���?)�����؛�ny�����˸�5����>].���w5�o�����Y�����z-w�������a�ԣ�邇�!��*j�x�J�!�qX��]�1���q@��������?�S��p�F*�	�,gV���X�PATp'9�xr��c�������*��cŬ=?�ή�	t��(ʈV���Z(��N�*�����Y�?,�s~��?��X�Rj������������K���`>y�*�<��Q��t�g�/#�Cwl�U��ZS�0&��^Pbҹr����K6��`>y��8���)H��'�����)�Ss����}�7�=���-���W��(d8�q�Gz�4{k�й4��[����z��\��~���S��rĂ�{	���TF���59/�!��Q�z�b9�^���˛��L���N�PN��֬ǆ�hMȄ���,����:귋�}�͕����,-o��ҕ������<��]c��~mL����V�����/kSi�
m�w�=�k����
h���ؖԇB�Q<��s�1�
X���2,a@;C(H��~�>���j�`L�37�����jlv�8-:��=��F��#0�n�-iH@1����@�=�dí��]#���a�^נ����X����C����X�.7����:4�n��UIи��ta�}�܉' :�s$%����y��I����BD��x��P�����������[(��ޡ�hY�V���4�3,Z��20ϗ[�ﵟ�5��e3�d�ڰt=h9�����v�	���P:���2��M�A�"w>��P�c-D��G���B��t���n�?�r������wk�����Ũ���k�{~z���$ǃWOl*_�����?�h.�lK�t��uZ�R�s&�U�#ΜQA���|������~�;��~b�2cK���cɈ
�/�Ch�+��P�.��&��f'�+OI^���+~�+&>/G9�M�B��n9�������Z���O��j����G��
r x� �,��u�[����w���[|�����a��ygK�*e]�0�<�vm��䍙;�l�}Mv��|v�0�k}��� }�������頾�v2���pϙ�:#H��3y�/�x��H��=����aZ�K�EmKaMBzF;X��*�������������8��\�����0��
�z�u�t/�?]������X�o
'��gĊ�y	׶WA�B�>��=7����}�_���@��?�z���!�5$�n&���Nwa-��
I�K�i}��K�{��80z�D,�^���ai�ҽ�U����6;D�c������{I�N��<c�=
F[��ǝ�R�w٥�����̯������Ѣ�,���:l����X,Sue�LZ&dU���}^&�B�St����;��
n'��wA��q*��R�h�� h�rp� Ǯ�{��1Opr��l1K��9n��9=Nׅ����t��]Е|��#b����#�^��p�&�vL����m������h%�������׹� �L Y%@������u�ޘ$�����^�����	Q{f��E�熘l]yL�v�����nx����`O�v��b>�h�����k�~��Q;��v��8d����?,)G���l��x量� %�՗Z�k���o� ��5�D���z.��p��eH�ے���Z=.z� ����"^�
^�TX�H��Sb�̅.���n��Q�c;ɻAI��]>�o������
ҟ��O�wj ��~r��r��^*M+l!����-.�����������H.MF���Ч��O��;��"�v���w�^�A��۴*/w.g��_nv��`�C)�
eG�K����-�)�՘���>?9�1s�ͣ�=��	�}�r��l�"�]�j���Ӈ���������}�;�pE^_�Y��$�|^L��8>�R�y��t�H�*N��b�=���r��\�}X,�=��E��?J��P�VUD�4�A�V��,�b��zD��5KH��{��>���̊ʳ�\���m��[��w�0�4p�j\B*y���N����Jzc_���9�Y_�[0�c�Ї��c?���I1���M���O����X8o��.�ӌ-fȅ¾�X$`w���~
�?16����<87ҍ��+�]��E��a���S���(���R����4e��H�YP�������v��G�"-6�>��>|��?�ݑ�/��#.F]~ ��߰���É琦6�k�M?�.�(0�VpW9.t[SgLw���9մ�'~��ܒx�=�Lό-�*����`��a�k��JB��P��N�J��V��RF�D�jw$Na��.,��Zφ#a5o����4%�F���ed�FK-�]L�=6Ӈ�|�iX
D�Ax��{����8{�����F��uq>ђ����I�=�ӏ@J����� �Kw���4��;ĺ�f��A��@/�3�������b4\��̪�`Ҹ�O�_�d�&@
�D�j�"_n�7�%e���2��iޥ�֚���Fz̾䏃q��Ҹ
:+���؋S���ցɄȮ E��x�-�W�ZFT��7)xG�����=����W-��_�UAԏ���(��t ˟s1~��!)R�	�R�\&�G�o�]�D�M����cH�<26��#�	9;��f�q�4����Z'�t �bV:[��[��9���*ݏ�O��#Y'�?�J�bZ��((�N$��𶆒^}�c妼oc�q;AL+s�d!���V�*]\ �Ud
�A�]XU>X��$�p9��O��/�-�Y��R�O �r���f����592��6 ����bSڼ�.Q�AٗRuy	-��u1��;�y/��=��4/ܡLw�٪��Ud�tu�X��z��}?^z
�?|���rwRhm~-����������t�ьUr �� ���-����F��J'�����鵱RP����ӂ�s�i���Z11V�\<��{6ڻ�r����ư��i0=�W�Lq#�"���GD��j(�cU_���<�������N���p/����E=�i��n@�2�}7Sp��K�TG��5��6������kU1MO*C���[��G^'}d������w�4N���4�YF�S㎴Wk�=���[�{���j�����_���q8m�Z�s4���/}���V�2t�wa�.Fa~���/�»Z:y#�M������сy��`��w@�z�*Ǫ��9n1 m
X�
�}$ܠ<�E�E��y��E;ǆޗ�]��]
����ǯ����L.Ԡ.mh����6X��=�%
�2���_Z\B8�j�A��֊Lɂ��L���; ˹��=��m�+Op��a�Rh3o�X��
L7��qd�,)D��gT��ڍ�c+yk�x��p�l�9��l~��O�RQ��+��\���I�s��{������|i��������T�L9z,l���9wӬW�\��R��Ԋz���b\G���#��}�
�����̯�܌j�H��A6m��ߊ�}H ��؋���ԣ�m��|\1�����",�c]��i��������I��Q�����C����@E�a��:�,�2��Q�z"�J'#����r��5O>-��N��O*?=��d�LXJs�c�a��װG�3�@��hX�l"���L/\(a�aF9&O;��$L��؂:�R��m�"饲������3�B���ц��Y���:گ�	"�	��e=��殺X4�,��T����՛V7O���]�����Գ<�A��5^�[��h���ķ�4�}��{*����m-��4u����#��.�ꂋ+I��7{�R6�GP�y`���{���MsӃ'7,\;s��W��@�ZT�Ϣ�.9ӄ����CQtB3Y+X�;����|2�ǽ�4�����)$:�h�
�F$� �{�Qna�شš{E��Ș��#�/<L���d1�Ƣk文Y��b� �!)I���hW�1�8�ƻ���c@%y �	�(Ckl����s�Hs�{.���v�_���w��� ���r㏂f�wD��������Ln�A�R+H�3C�Kx���N�y��Q�#g��P�׽��<<f�a���O� M��5���a�]��.�q��VHb���V�@�,�ھ�3l�B�[���0zs�X7X�&}�a��Y�`�B�+i���'ȿ�Gk����ظxO��������<�{2
ɺ�*�&w/~���z�"�Mq�vKvv@���(HM���4��%�i�E;^��*2Y:2�Q�qH+��}����%O�����*j{P}�Wd<�v��<GO{n�����5��>��֢11'N.)g��w%Z*�Zˊ��½����e&�xsZ��]�|����@�� �t�}6��Q��0iݷ��	o�z.��8D��@�q5u���D��*$m���E(ua������UFKW \E�x6a��l[.��v< ��Wx4�%�˭�G����j�_˝{��5��y��O� �CT�dnYq�'�5r�b��9Ϝ�s<��Z�J�m.,��
��U���^��ԡ�����|����o�jX�f�I���Ӡ�E��G���d{6^����Y�9v� a�U�y��Y�j�=z�����-խү΃�
�c���x���>�������_뽕=t���<G{J��'��D!!�y�Hw �9>6�^J�{[A|
iP�J��X��Wb�յJ~��짹��,�M��VM+d,t-6QJ�o�T�T�~`��ֈ�.�YVX$&ac�G�a�v���M��6iSAC�P �l)�<��Z!�af��LC.6��K.��r{B�^|X�'�@~��L���,/<%��*��kPv�yE�ށE��Ｆ��#Z���ޝ��(��e��O� 鐖� 	�$�Ȥ�u[]07��B0Z���a�"_q�Μ.�4���ʼ�k��/a�d���ܙfM�ow��k= �D�:P��y���l��##��AM8��ppY�MJ
�6}�j��I�J=Y�k"U�����UE��e��֤�]o�X�I��ҕ3]E�M�MC�Ɲ�����x�8
��.A��[���8�&G�ܜ������ߠ�X,��w�G�4JD^ėX��w|��H�<���}�<�~/���O� ��JC?�������ܹ���R���U��(ˡy��n��W���Y��]�}�U����N\}s�ȷZ�ݼ����V���^��9���	Mam#�f�\^�FX\�庿Y*�45^�a4S	��uw �0�&CC�+S�@s��m��=�$
R�/�	, !�T��ET���F�ݩ<�,B��R���R$f�Yɚ���2�f.q�5j�w7�����y��Ҍ��!p$[��)g/a�Hma������6�B\��N%��P]��T��t���Q������(�w�r?���<qw�m��ZH(�4A�����u���>UZ �Y����jf��HH߳ۏ��yF9�I$��"!-Y���@��{�/����ӕ�@��B}��	�����{��F�YQz2I8��\��C��D�l�p�
�zy�M"������L�/��j��c�U�t�G��
tE2�u�Q��5��\k��́}v��r�n|��jk����5�f���nO��oOy���z���L�|�eoh�.]8zh�~�єsZYQ/�iٸ�6_�4�Co&�@h���y2j��w�.q�����2�T�Q�R.,�����ϫ|�%W��.���Y�B�`�����Ó(H|��6�KA6����[	����q�y�n׷���Q$��T������W�hOD��0NLb��Hv%�
����Q�S��T��j��C�@�pK,�|&�}C��F}�"
���uTE�l�6y��HјJDR��(<�\T�Xl�v?wҎ(��F�6A�R�`��"+tR��5zV��o@�D򑛗�O��U��Fi��uV���1zb�)X�Ȫ�LϪK���$ˇ�A�C��-(������.SSl����\Y7|ᄗHN���-)]M_��;�/�=���4ę`cǎx����5U�TDE�8*�������=�c���?D���˭
y	�w�!��:�'ne���*�'{��t8,S
�Xx?�}S�1�]���ߟ�P2��z��
��2�u���ueV�r_3bE�g�A[@9��}�f̏L����~.�m�V��l�@2�w�%��S+HZX������x dј��3�H���Yj��i�q��H߻��������q�>���ׁǐ����0�-�V.d��TU�-ɺ�姓��y��/,��
�ۼXi�4$׾y%�;�p<��������j�����HSK��Q�N�A�!�1�ޓ�DClY�[��:�zP�ZɗKGb��˳�����������"|J�!j�m�MѶ�5��i`+�rw�B��o��n�q�|�rz`V��n��V[�S�{G�&����ؖ<�AW�1cUZ�	��U
ol���#��Xmt���{ .	:.=����G�y�p�F�t���
���Kv}Qn��&#� �Ϟ�����h>3薖0|'=`��l��k�E�=0���6k˃�kg�h�_����/0��&o[D
�L�3�T�J=U���>��x�>[{�F�c�8�J�~[��W6id�]RQ��Pn$5��P��
�{׀�}w�RA��v�3aVeL׶"�Z䷍Jpe�M?��Q������`�{Ğ)lZ旓��NiNe0몰Z��YE�HW�ԥ�,m��MŦ��=&����d���Ao�s��4��=M�XŢ� �׫�DV����\Z�%���zM\)U?���SƋ�8�OfŖ�Mo���(;]�u��x,�4�Uz�-�S~�્���_s�7h�u �٤�6Չ���>� ����%&���"P����9���ק2��4�x+����_���]`�b=[ ��Nmi�/�ҙH����)�zTmD�pz�p��=��tĆ,a{�(��b� B *�)={�&K�1S��"��d�k�t��\⓻xk9�u��,��C4���&a˱}�%��V��7��V.(l?�P}V�qA���tn3��t�m�D����v���?T���Z�m���XD`	t	��B�X��`8$r�(�8ѫ�ݗ[����ͱ����8d$%,$��<�&��
�T��<���a���I�51�}�����rmӅ�S�����f--���A4|}��v���y7��B;^��h�'�)����������A ��A���P���U+L����?M&�v[��l�D��I�r�L%��BP
�6�ף�0�cE�V�m+�V*隅�h\q�&���z�U��җA�z�j�n�/���y�tYRN�|)Jf[}�l��,-��B�6w��fzZ��}2��B�Iu�آ��W��w���G�Q뚱��#��duѰDE�w�_$uQ�9Ev�������t��s6�A��R��6q�)�%w<|��υO��*��	+��y=:��E�w������߷X�4[E�#��$�V7}��]�j(����CX�;Taz��gYu_h�� �1��~��:��Mk,��U]�=B�fUI|��"0��W����^z���K��)�6�f[�h|��k�����\}f����{���4
�<�A0i��y� %�d� ee#D9'��pr;�Q��ڭd���˂���n�a�����t�E���
���Ki�]�ER�\�@������x[О�m=�� 8�S�>� �;(E��aA=�%8��h��Y+*��4�ƚ��[���h�>��q��'^���R����/p�a3�\�_�v���W����q�7�д4�9	��*؁S��"ʞ��*��(.�_
��������\l�⼏g��#����L/H�Cμ,��W�8�
s6�"1s��J���y�����p��bN� I�_�<U���^(X�"{v0kpC�l��_WL'�8.��A������[��N�՘t^[
%�Y*5f���J�Ւ�a�o(�q�3�![��Y�)ݧ{��ny����D��XA1���I��Do�{�
�=y�0KY�EC�=�߷s�,���:v5��ZA�ջ�PP

���'��8��k������> �a��R��KW`��$<T��/������9��ݜ-ZQ�2=X�uMj�\��������<sHz��u��G�4
Rir��jB�wJ8��>�C��/��F ��Z m�Sy���f,E(���*?�+�a!�Q �"�$$Y�zg�l���.B���b\������m]�&zFkC?�30����/���RT/𨨩�!�'�G��'��֘���a�z|��'$��"�E����g��2���p�}��+�:��@PK�v�=&��H���.j�i�7��Q>�Q�,@�Gop����r�
}�0^������bG�d_���S˓W�L�%�x^ݖt���h(؞c�����1�=��8��-,�?&dk��Ҏ|��/��S(��d�4R�OY�߹`�-��/�[Y�ݢ=L>�.�����{S����cZ�}K�<���ik��ȧ�����ilW�G�~ۭ�Ɲ�Af�G\I�P�Σ �&���U2
�h{�]U����,twj��2�pAO�u+=QMj�	�?��{b�pӍ�y������u7:em��^�>��dJW�[����Mf�9j���2���+���@��Z~�a�ڌe��9��⋸��4���Ů`/h%�\�L�~��$���+�mk���`���L�7�4Y.l��;�O�uɚζub��}v)�!0~/�|-IB�ܽX�?�Œ*��*i�;��nq W$�d�5Z�DII�7�u���{����x.��<
��ۚ:<�}�7�b���M�3_GU��4ڍ�'�]U��Gm!�.0ګ���{���at��DKb�U�4��[$}��V�У�6`s��8���u㱓�����!K-��$-��U*�I��ʠ�ù�9��[��o8���h���с;��9P�3,�.���WF[�ڄ3�,�X���7�����Jm�Ħ0���ؼ��^����z��y�P�d����LOG�h,+HyVw	�C�d�(�� EM��J�
VK4�-{�Ck�m+Z��XOA�i�~�s������3��WW0A�VG�J�77R^�"�+՛��E�Ę�FO�7d��@��B�LJ���J$E�NҌ��<=��l
�0]{>�����kӘ�Ҍ�?`�d1�Oq�
/�4!�C���jV����f.���0׏��I8��G
^Z1^���0��wK���}��yl+~~Q�F����6Q��5�Ω��r���5�5�U�m<��z?���K�@:)ש}н�U�_\hƉʤ�5�����w�/����[i��j7^�t15$��% ��V��c�ԣ�8��ʠ�����K�_&J`Z���6���e�_��G�u��3I��n�؁���B�PA�OŌ.���4e� o���N���w#!F�lC���BH&�����,�2�׷�aj�(�򑼂���c�Rǘ&���f���M��G�ޅ1a�:�V����75(&Ҡْ��q����Sd�䡵��E��Ԁ�%�!U�t���a3.���J��=���.��x����q��Jzdi
��yx���f2�qG��{��O�c�8�	��gFI��Ix�oNb�Mo�>ۘ�>�8��:�"|�MM�ª�'YtS�T��?�R��?"�}'�jJ;�Wh�@�&(F> LN�3�Q�b>����Ok5���[4�_���q�ၞ
�G��kT�@��]i���T	������ ��=��V^�n�0�a���\@S.�]��r�F-� )Œґ
��^G����!�1�W�ƞY�()���S1u���!�Mi�!�T~=:G�8�s,�� ���c7�c��A�"�p���,j�� ���[mvz��kx�D��<N���S�vR����w\!���#)LaU��`�8S%���KG�[_�ﯰ<��c�X� V�eE$�Ӕ�IA
��b����	7<��T6�wY;#���_޴V��k_�
�U��ѯ�0˷�KtP���@����~oZ*W�S�W�tZ��7J�*�r?B��x}���"�W��*��gQB�Q���1��l�-膭3�J��>	�a#�l�`.U^���&E[f��v��2�gnS��]#���B�SՊ��_��ir��d ��]'/����{	c�Ol7;X>�D�h���$w�M�q���z`���1��V?�{��.Wx�}���&w�#I[?����cS=&�Eh��"��A��U�pM����'}� ^��?�0a�es��aK��G��fr��!t� �zf��� ԧ6Q�ʈC�@
���%��G��-���xw;4J(|7�1��}n��7+�X�~;ӕaȦ$�K���J�zV�$`jerٿl��'eJ���ti���i+[q���Bb�ƭ�K���a�K�~x�1����%qn�8��R2����>�%��ϣ)�'kx�\cV��v��{@0�ū�J�'4�&Z>~��~�?�O�K�6�м��n	9˯1~fv��6d_zJt���3L)ΰRݐ�1q���,Z8�$X�ֲ�<�ԧZB�M~�$,�t�B��ۮk�LƮ�@�7�݌^Q__gei��%*Z�2;���eX��|�jcir,��1�� �R��ҶZ��/�6@8����^^��
x7;n�E��{��K��P��z���6('���[I��i/����?��_�����H�/�1P#G!�+��=s1���x�Q���<*ʹDg�~�I9��7�	��x��d��BuΖ9N:��7�B��Q��|O��㚫��+�ngQc\ث����%~�������6��~A�9�G9������0���wrior^��DZXa��9���F5��8��TJ��g�����'�B�x~�^�W�����7|��}����Dw�`9���}�Tue��-�r�����������F�J,�RԪ�DӰe��Ё`��@�	B�"�5���V�&ZAҴ���P铛�$L�Q]���7�#�s@�I���h��Y"��b1�(�Nt3�S�)F�����K͛u_�f���ﮙ�ق�Hcb�0������+$�R� ��3qһ�����T�jB�7������GXI�&��/���˾č_��Y����d²v�I��%h��W�?rԄ��3.	e��~Um|���Mhuo4�:����}x���� ��#k����`�_�Ig潥<1W��:MZ�5KI����*�e���'|k�Ih�����e�p�Fc�����S��wG$2M` ����院�����@I��YL�%	L��������}��^�>��/��4R�H���Oxu^c9 )* pP��Q_�Z�h��}3��#w��b��3�5��
7�ô�{�o�?L��6��_�	o�^���AA'ㅯZ␾UJ���L!�5�����9�o9,�-��%
��[��bLI�$�e�y���r����S�}p<�&��sƀ$,x�p��^ߥa���`,aW7�|k�9�cd�䙮d ��q���-��ͺݙ8gpw��$�p�O�'�0�������/���>�>|�c?�N����3G�c��<\jY�q<�ʱt����	S?_�dd��I�c��=Y��zN�x/þ	a�x��+���v��|�!�	��	CXA��/�R>�M��:���bU�~��f�-��1�н�������q/���lчIpu�H��6�x���`C����j��<�\��y}�%�6
�đR���{kT����e��E����a��ml~�Dc�ҽ��/s���4�SR0*��5Ӟ�*4��S��ӫ��K��m���9�4��<�?G͜�E#템"�M��39��_r��:{&�;ڻIJ�8U,��J���J���畕3YD�q^v���8E��J��xzG����}���M_�ܬ��|ɛ����ƺy������� �3a]��V��v 
w�)�`��r�$����
奞M��Q���#�8i�k ��dH��Ya/h��椱� ]t<ɑeŘ5LnAT�	CۡH�ҫe����=��0�-ބ�Ͻ	����!ĭ�]@��Ӑ��A~cI�l�'�X|s#y6@��vz.���_�2.����}l��5|���W��c��W>�ۥl9;�` /b`��̮��g?z`�菥!t�yWE.��h���X�W�f��l�Q����Q�>�k!����v7L+\���&�N+o�N��n��J+s���]Q4��%��٠D}м��![� �9
L^�yk��om6)៟�dL{���KJހ���$`)JO	�[+�F.�ob.ȟ5VhBP��Xk��]P$��f++~4�)�F9!b�K���X.���d"2 �ҹ����d�^B�
�a�;�{H�D� �|��{Cc�^��_��5�Y���� mq����qB������=f���Y(��3�P��3����F�=A�@�t��d_H)�r�E� ��
���#��e�I���x�F�L CV�s~@酎(Gd�%�he�ʙe�zV�⣼J�ڢrl��U�fڣ5�����J����Xa�{uqE)	{r�7�l��� h*/�x:�N.u�B�9�!�a���w�lm��joJ7|�]��>����")����
��V���TE�5[�,Z�
�V/����fښ�M·[Ç�k�~��ˤc��8��;CPV�����!��*?�ζ�ܣ��R	�D]���	b�l�G�q�t0��/0�s��8�wp�n�m���W��j�k3S��:Q8H���������Y��F�YLޗ����O�������(H`�vo=�Ѐ޽O�S���˥�ެ�noDF��:�1��E����5l�u�pn,��S�(n�&9p��u�Y�;
j�A��|Iu�۟������I��%�7����E˓�;v3�(P�nNXԾ�p�e�'*=cHi�%���?��3{0AZ��mD�&+7�r"\�7�?�w��,UE��'����h�OT�m��/S������;u��IE���
�Ҹ#CD|(������?l�u��Ig���p��Ѩ�!xL�k �k�G�ioJZ�IM����J"�ýq��!tHS��!ǟ��H���W��2Z9��pH��eq�W%�Vp�Ҝ�J�Rc*�KnZ��7̠%�z�C�>r�8��d�ru��a�@�pg�:g�(�7��j	�Y$���Z�#��yq!7���щHIo�O�_!��4N~�o��22�|�	*�ʳ�Zy�Wh�ji��� Jʓ�b��H���usv�*��W���<�a(GQɦ=0@Q�VCHIB��Cl�(o-Fi��l)��D�Y���`ԘS�!�`n���_pz~�0\G����ʾKtJ0TEU&�H��k��j�(	��-�����g���>�y?���1f��g��;EP�>�9K�X#6�2*q��-��])c���s�1������.���p��YCk?D�:%ؼ��J&N�i�Z�ݫe��N+���)�,$k�]Y+�w;�����D�+HS��:�Lk-C�X|ZT����mr=�!��cSd8���}!�rk�o9�pmH��J`stU%�o7���L��!����v����C�s ���!�зY�|�j�Q�v]�o�	I�����SJ��1 �a8��8$��:��W�1Ȓ� �����e�q	q_S:���f�+4��T�ͬ��P�9ӻєM��Zus�g��n�;�؋��lA�j�����a���kj�Vd�T�%=e�w�;\�e:�$R|�.�Or�|a�1z�\KkG����+�61��|�7��������R=��j���pa� �C�N��g����L�p��n��Y{���@I� �,MgKmSX�����0�k���о����0�L$$Y*܍�=!l�L��x��!�=YHL'+Ԝi�
@�(O��3�L��R���>^��m���u:�e��xn�֚/$8��0Z2��!6?��/.��Ե�¶�3{� 6M�۟� ���Z>�ڐV�<�q�3��u��[��� ��R��J4@�S�D��{�������b"s?"!��Yn���6p2U*%�g5^k1�~�l,Jf�ܺƸ�*V+�E�@U^�v>�蟙��������CRc�Q�`�-*��Y%�&�j��|��:������0��k�4�l-
k.��:7���t��F2�R�)�5?N��y_�S8��9�TB��=uh�}Jن�9�7�b�,8���ED��`
K�q���?�/�G"��Yf��Џ���Kr�u�D�^_�6!}�ճ�&E�ҡ��xb��_�X�!A�
Sz>��J��$�#�kJ�2�������̜����Z�AݙZ��{���6�*dZa�K-�O_�a#��CM�&
�h��2܊GR1��2<"]���ZF*@\OJ��
�B)�ZU�az?�&�D�߈� S�vLcsI=�r�R��ޫ�ig���U�dRVq�Y,�^ɑ��=H1��̣@]8�t���� C�.�Cy�/�@@�y~�$��:����#38��1Q:��P���*�%�t�|%�xX�+����>�ȭ����j X`4���yGP�����j,�Bb�y��Wg�O���Cj:;iQ�
���n.`o�^v�m�����O���U�M�`wˣ���"�T!��|QSJ�����2&#�� �TVr�d� y1`Ng�&��bV}�;�g �;�G�6�	�P��a%�<
��@W7^�l'�Y��V��)�^<�+ /�9��1�j3���qS��I�2��O��M��x:Ϋ� s��C��/����^��;���OM�s�|�=��KJ@����	�8����r�s�Ajv�B�&jM
��̝t=@|�z���c��gY������1͏�VG��.<�߹$	Q6�d7i���.z��0�W�ԋLeG�G��O&���U��2f0�X7d?��?ޥX
.�.�v냅f�iI�t������^CG��x��.�.��(ڡ�5ƿJ�22���w��O]t(��X�d�x����U�fI2�{-_��0��߻�+�;�hp����0Y��(v�RENB�вڇ�R��e$;e�}��Ţ:�l��H�k��B���n�hC=Dy�����'�&rBc	A�b��g���lV���9a'Mh��|(-!�Tڪu,�X&��BI�%t�!���	-sF�V��%p��&�nb����線j0��S�%�!����2N�I���[F��t�=C�ք�q_~ih��s�ju-�3l�ҧ�\�5ï �x(G��>�����~�5�����wn��?/��IP��ϋ�*H}���j���L&���� 4,,/<;��AJ��.xuRJV;��V��υ�%���QӴ^[�M+ё�%��3���\�^�z��8Y�!����,!{�,ǧ~Yo��GM[e�?�{�зYk�=ԕ��i]���Q�mNJq�Ӑ��"�C���"���m�٭�eٰqQ�c(\_�Ъ���*#
�B������#$�U��J+R/�"�,4\xR�ZA���U3�'c�� ����I'��
�(�������&�x��Ʉ�9������	�B�hSdD��1�+o�-O��V[���8SVB�e+$0�2�1]}�!�~�կ ���Ng���W"������(�f�<��U�l���U�WV^݀>�_\%.>��h�6����$��ќ%�b�=nA���Nc	����?k&�\#�NÓ�|��Kt�����j�X�|���o[?@bUUc1�� �����;7^����2�����ϱ��}4���ȺIg
O�n�&9�3��������Al3�]�V�,�k\'�C~^��z�|�t�����:�� �ʇF���U*����V��s>�����;b8)/W�e�I�M�a�'��1��N��8D�	���x�߼�Cz���n|b��@��9>�4y� M�yh^��|F|gM�1��8�y�5��N%v-��� !�d��'5*	*Oq���J!C��
�;�J���C�SŬ�
��>�3)r
fA��~
]�HI�ԧȆ3T[�.��#Y�+OAzF!�j�d�H�A�P�n�H�m�O6��)��)��o���/���c��{R�������7Y�&����J�>�@��ء��� �dTP�?3�-T,*���]V�{�()g� M�\�(+�y�|�@V��r�3z�7��2M-���¥}KI��⃪:(�Q/ԁ�C�>f�����
�r��aF\�[Od��-,��6�(`�"�}plg�[���\��b�~"�u2�.��&�[�s�����?�1�f�gL�4�F������ыK%�-��j�&!*BKDz�8F�K��x�a�*6j��ұi��1S�Q�a��U��o厝J�����H���ܴ��B'��Ҷ�rjGB��4Y��x�H9|�=����y�K�r����t�W�w�>}uyK7���7��k��(u�>L�t#\l��e{>�`�l ~(ξ�.�ܰ�\x
I�?+4m�zή�0A�eݑ看�a�%z/�s��喹h��>���W��T��B�g{5���>[����q�4���]!8�' ���`4��J�����ۀLSH5�x:~f�t�`}�44n��j�LdW|L�Kտ��\P��
�i�)�ٳ�A
�Rc�/��ҲjL��Ⱦ벁=�Y�8�� $�@�����U����B����ǅ;"3��Ps.<��$xW=_�k&ӕ�p'(m�g�wC^ȕ�� ������˼���8�0#2E����t[q�\@ɂYd�e��L�k]�$�`�2}6�$>�1�A)��%0�4UꚂ,�r&��lC�e�M�Ի�����d/���4��G���ڽ�l�ׁ�cXi�����\S��%9ڪ��A���� �mF�]�)��{���;1��-3Vu=(у��*���8�F�C��p$<����?�1�\������ �@�d=;��4�-|�[m��E��G]3$'��5�K
FFO9`�"S�v��{YJ]�`��E�y|�D��lک����!\�2�N���=p��7��2��[�>����oe����N�V�U:�Ǌk�:������)�s&����$6��Hcd#%.�ɑSZL�0@)����"����}@�_��ZX�4)^M���?�ܢ%�G��>���1-�w!hJ7G�yӪ^�@Pc���vmB�YE}2?;KWkC�Б�F�PW��}	���=7�8dr��c(A�!�N|��[a����vt�jaE��o4m��N��9��C�@G��l�o:[��/�p�W�{K����j5P�ѽ�|��������,���y��I�@�s�|���,�,a8��2�iKaV��t�oC��s�����Qδ��6漆p�5�x�x�1����fQ�x��������J.��2�훔�
������*��\h���9�x�n|K?������$���+K��?�K�|'�:h����Ȩ�S��>�\,�����fȽ�P
?�u��������KRU�-��۠��K��(��;�O"+l��]��y�&~����4be�:�c�w9����9�������Z�n6�8��1qGY�dX w:�F�f�o)����|k��y���̿����U	�&�j:�r�W�~'��W�ǢR^ܭ��{����=�y�v����M�Q�zdˊ֍Y@�
�1��[��iV�.�{�j�l��Q�O3}���VD����&�����x�r�#L�r����ym��{pNl¿�_�z4���O��,�ulH�;Ҳ���D�Wđ`!�Px�P~����-4a�vZk
�7VE�.��kPz���b�۳��6u�.)X��z_nHWLW���$Ś��C����}VQ�$ &����+�ݡ��Ѧԍ�u���Fg
o���}��6?���O�pga����ot���)�T�SZ�p��Ë�`~=&v� ���=�J0�U��^�wD�4� ���oer_��z�����5�($X`�X�������cY�=�C�s�Hi;V��Ā=��<��zI��0X���eiM�����4��O�|�R��D���,y@+�0w�"	rׄ��5�� Z�J
b�)r?�!D�ҫI�Q/����(s�����1����+3�L$?��F=gp�=I9�Tcp��L��	�16Q��k��2Ť���L�S6��K�v�}դJm6Z�.��o�'3��J��q�/��>kV�z	W&)�2��[ ��3/<  ����^�g���FAj�5k�u��f`���Տ&?f۶�E�.��J"�p���B���>$Z�}^!�\��ߥ{��U�t7�wx% ��Y�')�)�1�=�?Wr�����Ŷ�ڰ�@J�tg��$�@��o�}%�H�u�2�
�h|�P}�r?��=n`�{��Ǒ��^�G/#��Q��2�~�)?rގ�����
)o�G���Uⷬ�������F-?���t-�ʃ T�\����7̆�m�_?�4y�� !Ec�c���"��"�x�/ո��p`^�}���\&��7�G�_z��^�Q�)41�^\�c-�(�+U�B,ң��ֽ��E;��VJ=Q�`��i� Ѹp.�,����d�2���Ĵ>�]�>�3}�0K��[��|�ֽ�
(��RNF�"�`�nf���!�i;���%X�=[�D871��r���U�u�i�%;G,
B
���T�\і�F��#Pf����ܤ�|��aX)��o�G��-x��ZQ�ZF��<퓜��H���ƹ߹HQ��dO��,0��r�����/ۦ5]����j�P�H���D�dPD�P�k��$*Z+������QE��2҅��i��Ɉ3�"���W�LV�ʽU�k[�K���+R˹��>�Jj8��䪴Y�^m��;ƿ�G(,{�|�P�+��4ߩ�c5�R��e��4�d�g��0�eo��}O��1Qs�M�t���g���lO*�"B:�8]_�c�����y�.��Za$`�ؔ��F�:Yl��Bv!A�f�Av{a&$?�!�����X���x��8�p+Y��D���l����]QҎ�~W����٦�l�D����C�
3D������oQrK��M�%�!��+.=�\�cHm�E XH�P��W���l2��*�΋�� �Z�y��,>�BA��� ��-.��@ ��3/���n�D� k���	�z��3��u���� BM*��4�,�;���|�ޫ�Y�J�<->���k����s�����sT���<�۴RP�M6�e�yL�p,��ŗ��
d�'�S(H��ޅg��7�4A�I�5��cR:�D3��q�<��<n���Geo��y���P�Hg[`{O����y���ƌ��\�v�liC(QB��
�K��URJ�p��+��w!F�]�ͩ��r�P��d�Ts^t�B�����յ�&���L��֌@�(u6ݢ��d8�i�G��+J��TH�~��$�O�����kC,D�C�g�g������L}�
�*�Mf{�4���GϺt��Al������墍��Eh?��bl	v~0+��@�-w�����I�`l!�)	O�_��"�G�z���ʴ�]�
�e(!��=۲[1_]�jՃ��N+��b���0�
��k�W�l׉��|���,8��l ��_�|8E*�_6w#���01�/�e���3��R�i��T��# c��E4���b��C��Q ����O��dQN��m�X��
���\��񷞟��㘢4��4�7�8��H��?'G���a�{�Rfc4$B�ӽ�����A(s;(�@�~Ғ�j5�2:�;�3ʸ'P�^�92Z"��H\K�ɯ��֜��QWŞ�������[�F����9K��]�x��з�4n��-��޴z�˥�[+��V�|�4<lq�F���R�(_�dR§oy���5��f�h��$FLZq
�\_�!E�S��\�eQ�P� "�7����s����Wv�E��*H
-��C-��8G-��ʨ~t	&L�{4�V[.P��JQ���A��8Tߞ�a��]_���S�t�WrZY�~L/ߌ��;�V������w�=<ƨ�N���D�U�E9[�U�&�a"qk^��S|���jd��yG�U>W(%��d��s(H���ݟ��7V-�#�u���C��l.WO�(��r��� �ܞza����q�:�5#B���J�V�!/���������?���役\�OI��t��9W�D�a5����d���'u�p�)�k�/��&]o/���i]�� 
�0�ͦ�C��7�Q:A�z��+p�8/<�CAҨ2���W��f!�rQ�Ҁ�e�|��b>�����ے7[r�^�!W���磰DI��ٺ�Ľ�K�QXa�.��lȭ=yr�m�j�w'��&�a]s��&{i��֤�E�Kˀ����#���i�@)a��� 7s�o��s��L- L隸��{�^��2��S���+K�K�3�U4����셜䒌Iy��Lz�X8���օ��iAqj���
=]GB4;D�t�O �e����C}G�䍕`h+I�ϯx�;9�����V�,�k]�{�vɑ�\����RP��#�sc���k6Λ� !������ڷd��#�Լ����sυ��S(H�����J}Ұ�YϺ��H��^��c��� ���K�}jl��kth�U{<_��Ap9�a�����,�� 3��<����睄K�O�"����$ ��$� �t�EZi�Ar��'�Z_��تv{b��h_ZR
Z?2�6��%e�}�a����~�
�p^�}wfx|	�2~d�=C	=����\�U�\q�u�ZХ�~~�ւ�8�s
Z�P=���g�3��ż���(E{b��{p������2G5�S�a���{s���?4ܣ���
����9��~�-�S����Nu*��ޛ���-���{ڀ�i����B P* ']|qK`�E�}m-��}��,�;ԭ�.�y��T����D��tc��D&ڐ2�G�܍
i ��Y(��5�'��M[s���ҍ��TV�א�e���� ��"�1��/*P��'�[��� ���.�`9���{BM^=��i�W�&D@�#���DI;���^qs�X+'ZA��m�x�?RF��6�a\{+�k6����e^��/hO�b��xWj��2�.'ѽ�T:�Q��g�#�N�{��-@���xҦ�ؓ��0L�_��i��˰�����P��<��	��Qq
)n�/0g�	��xn{�9D���M���	}f��_"g�C�H�I�r��؃�n��~c��[��Ͱ�FD[#�MC���N�Ԡ�Z_r][�Ӷr�쁰Kl��*bV	⟓�+�E=����4��!����w �p�Z�)��Yx��Y&��|Bi���M:3�H,a2���@�C��^U*��g�\�g���KM:6Ju�������)�tcC�����m�>q�w��L2�����`B����rG߂�I�Yp�=ݳG��ytd�T\a�����{l�����M5��gVW�E5��q�}�ԡ��C���(L�W�/T�+�5�z��)��/) ����T
�&�c��7 �'�_b�c��֪����K
Z�h�R�nw����G"���nR3h��.�Չ&I��o��ͩ~	+��E�+z�=l���%��F=�F3V��ɔ�[���@:vS�n�����U��R[h(����/8F�̐�� �Q�8����]��ھ����r�:dn~��-���xA�Qh����ݣ%�s�����o�E����R;&:��As��o��BW�i���cu�Z�#��ް2��L=�����%�y�z78p�<���i��W�7�������n>%��?�
�4���H�O?&�DqJ�g�(`crw�e�qA`�Ĥ�:�|m�3���v���<�����̙@���FU�3�HƯ�Q��&��
�k<rk�䈰֊ZK��`�{B��yÂ�1�������;M��¯����6���I<��އ� ����'t ���`�������w��sBc���4����j��/��ѿ0{�e/�T9���0>6��
�}�vS�ïM�����s��|#��B���C�i�u��|1�㼇�mԬsUu��$OiD/csp��)�4�M��S�T�-
��Ի�"�8��ղ~�=/r!�Ų(�C�w:��g���i ��\xv�5ƠA:��4�r���ި<����AϕW�.����t|�Б-��P�4,��T�p���G�mG�hL��YS�x�?wN���@�R��;���4Q)�
ׄ�.%a�5�4G���i��.�l����4^�u�D����&���DR�Zd\_kd��W
>=��016���{&�t���h�S���ʵ��@y���z,%bJ��a�M���~t��|�����o}�0*�`dK\��2LR�g>��Ę���.�4?��cU҃�y��pJ)G��y��|�p&��#�G�p�x����쬆Sr�3�9!�%9����GoX��(Ya	Ǣ��:KM���=��P�D⌤V�.��2�Qʖ&��7.!R˒�_~VCn�^҆Q�#�6�}j:���6V�r�x�*����̏D[{�G�P���$��mhaǵc+P�Y��@�E.�<!�y/�Q~��Br&<���bZ*��dy "�K��A���t]��􎈃�k]8=�_!�J��Q�q#S�Aܳ�?�k��jY|P�$�����l 6�����gFYf�+˖�h �G��pV��v�J�����M��[O� �Hd���.F|��t;+R(?��]��#�.5Z������pT�խ5���|=���ݨe*މ��e�yf�\A��փv<Yk�+9(�6�sӦ��]8(fR���+6zI���>3U_E�s-υ�8��y'��-����|�RAZ�Z2����W��l?)F�����K�5����d�Ĝ�:8g��&��@J�3�U}Ƿăxő�q�=H�������ù��)F��bɻ51��P�t��~�X��-�u�Rxjs�?�[���G��?A1a��`�������' ����ѭ�9O����Վ���ԾE��"���Ρ�{i����/4=����4
�7n/`s�:�y+?I�D���B@&݋7xf��1�6�)W
��۸�6Ov7�������l��6E���� ��[��qLF����-st�v1�V���}��s��V��R?�q�F�np�\�� 3�_���m�%|q�aY5������U�^�91~Yh*m4XH�hpē�GR�E�-�+��s�y	C(EzdG鴀4�̜�+1�*�T��{��M1�ك0ع�qi�.�}�IML,i���lRv2J�����J /�{p��a�
����<=堟;��r"�L�
�����.��ڪ�L�;# 7tx���ͫ�+��v���Z^B�:�ɪ)���$H�����q�f?�ÌH�rɒ�"���ଣ��y�����5_1p��i�=�Ӧ�U/q���/���C�B�]�n�?�_D!Z���T�=z��qE��~�
�V٫�N���w�K��%�A��<�(�|W��2s�т8Mh����g\0"H�ŵb�dPD�JV���׃���(H6�+CN�
I+ͅ�@������r{MJ�S[�V��ͨw�͹��~���Ko��.�2��<G�8��{��t�R����W���a���6R���r(���-����{Ay��kY���'W�JK5�o��~��y��(;/5�)�|I�ZE�3��N��'�!m�Y*�w�/Zb�;�2%�ͷ!���D��ЫΗ+�2�y�e��,��~���z[=z�Rk���p�I��
�/��d�GnW�o&9���x0��k��_�nN ���ң৹�]$�3�K3��@�7�1�x��|�*u��z&������ �!Ji􈮗�S���-������+��h܋@.݅<n���Ъ/,��`Ύ&�) ��j�Z/��ɷ�
'�-�ut��H�I$�j#���?��8~����W2^4[��"������H�$���� n;���W����)$`�1%5:�f1����v��P�d1'a]���`s�f��h./3A��w�v2��,C�J�~/��R�G1*�܌��3��<��ܓ|@_�aϘ":&�P��OS�ѥ����
5��@��M7����h���OTCMG{ubn�)+EG���9�0��2�}k�F���<N�*�����un� ��c Z_����n
�A�P��P}<��}�=�H����*��	���� ��(8yD�a�t��;_Ȁ�јԖ̙�L�3�r �����Xa�`;���y��-���&1�®Nb���T�����4�����o���$S��&LI;σS(Hτ�/�\�P��K2�<���Y��C|�sK���y�p�1-��o�v)E���!�J���J��K$x<��
�Oic~_=��F�����QO<-�KL���^�Z���m��(��_�/ȈS��Ip,���*HP��S�h5��0q)݅um�[�쐝���l�Z_a4G����U,���� ���E��D�&�o��cA�\:r�����=��lcm.}`�ۆ��n��b�)2tw�}*M
�r��V>�����i^��0� S�*�����&=��z ��[��w� �%Υ�Ɨ~��ũ�[���wi�~�p���Ǚ\�o"�U�'���!�����[�`�9��P��]��4?��01���W���A(�#��}j�	��^Q;%�4܈����]���V���G��A(�&Kxɽq�b�0�H�d	=u�n�I���Z�g�׼Vׅa�i-��d	��Vr.У<�x�q�%C�ݟ��i����O� �K�:����wq��t�i�@�}���s�E��vΠ$���Y��)I����`��NT�{A1���Y��F����8ƣ:�F���'�#���	t�LA����O~u	�H��Ԫ�>��G7�[)�4��n;���T��o4�pV������X�YST~_��AK��{"l\���B�FA:
NϷ/�H� N���DI��p4�1��Bl��O�ʥ(´ԥIȫB��
]+2�h5��lu��\�cRۏ���x�̠�*�Y�}�󲽊�"�wX��z���U5+�]6n��.��g��F�9�/�4�폕ۏ�)���g)�Fjl1��Q8Ԧ�zFXw� E��5��b���23	HY  .��|+FQ�����Ŋ�]&�^��C�ue�����BnJ�:����p��2T��o�}���B{�}Oh��O{`�(Ik����k�a��k�5	krٙ#T��{4�W5g�JEK��}��S^��W*K�: B�Ƿ�{�4��~����s�Wp��߻�Y[�l"��_L^r7d����@��XX�d�����%{=�LC�N���E��j.)�}>`p�ss����o�9�۽Wf.҄�evYY�%L�����
�p�+K{�x��d����(�"c�c��m����l��{N� �{ؚο�a����Z��=���m���Б��g�=������f���dU�l.i'����~�H���W	�R�Hԗ�sBk�9R#�F�g�MQh78�����+��R1�o�^����Q��\I�p��b��t�
�B��^��QI�>���y��y����&�'A�hI,�Q9A�Y!:7mIQ�,��kY��y�X��vRF�Z*Fk��vQi���鬜D@�1�ȻS�>~�M���+�U�O#�a�ˀ����6�x��B���\�J�
�j���rzρW,��|.�� �F��h�4����ʗ����:�k�ڌ�,.�~f�R��s��Y�=�p��Ie��ϫ e��O�f$��H��<�.��p�
s�9($N�/r�,�H�zB��Y�D���2[�^+��J�l%��z�V���Hh�J�d�2E�#$O�܅)F�2J+}����w��n1�#���6�e�bQadL�t��Y]�}+1E��9��P���  �?�~���A�]v#7N��\��{�e��su�d��眻�4�B����-f�A�`���K�����̼�	�4ݾ�c�?0� Pl�$�>��Kd�]kE�_F悸��\n��X.@�h-�1�����~�p��ò(������숭�*>�5�G���%X���i���釳*(�R�*v*�+V<���Ia~a7�I�n��7׎͠����1�ߍ�dw��\�av�/�>���H�F����X* ��{�6���QrkVCN==�tBt��;~�_y�6H�s�χ��V�ߗ-5��/R0�v������#N���WA�=���ÿ�C  >��L3s-���VK�=�=C�^�B�E[���%u�=
�FA�!'��R� ��GY�v)��jtmd�3��j�ҵ�Y!���������M�s1�7��ꄼ�q��h�_gi*�r�+l�j`���#�9���f$��WgV"BĶ4�V�j�|�%OB���@Cs����&?<{������0"���S_y)TT�[�Ke��-�t��Z�鄻�c��}NS�ܠ��`h���ǰ-	�
���|���ʤ/��҆J�� b����i�1��|�L<�}������>I+R\�:�����y̭�����ˈ�����H�Ĺ���b8���2&�f��mE�QtA�$��Gd+\��	��)��rN46Ϸ���`<��фw� �E��;�/H!�R��%Z�t� �R�_�ok2Hyhܥ{��a*b�0��슾kulm�_�~�����V4�1bW�]TY>o߇7�o���kO�w�ʚ�+��'Gя;� -Q�󴩰�v��o�4R6^a�H���X�u���i+����G@��ؘ)��M�c
|Q0 �k1ȅ���Jϒ � RL�̄�-}?� �A^�Z'���(�2h]�.Һ� ����[�$�K���$+f�1d���ۏ�VA�,�IM`����A��_�.�94�#F�2�!#r�bN��YLZ�,j�j��c)l�'4:'��Vw֔J�Y"��<ں�@f�2�"8�jur�(ղ��D�{-�U�9�QP�?Ŋ@!g2vt�?(��^4G��g�S�u�U��g���ϱ�ƙm�}}��\Z��Xt�d�O�N��|�l��\���B2_��NR��p`tO���~Z��-��[q���Dj�\ۄv�_:�11-��
������m1�o��4���T�]��a7ii�#���&�u��WR'#)I�
�\3�������[�n�0^�U��B�#D�G������AW�!w띪�uN��.dF`HM���`�����cr(�*ʤ~3R���el��y)Q�E6�Ƹ1�ʮS81��*��o�)#�ce{}��6�QWȖ��8F]�B>#�C|��V�w�=���<��U�9ߐk ��>�;�B)4���Y��ڊO�T���z�>ܨ=��R�mqJF!�+2�D����O�AnC�By]Zu��a���Dc��0���=C�>@�G��1d���F�~/����_�,�)=�_� �e��&����D"*�4C�n��6e�t.��S�;�P�uŧ�����V���G!W�dV�߳7�L���n��!0����a��"pE��J��6"U)I���
;И�Ѐ�/8x�OAֹpi��ܕ|G��+n��Y��h�*��wt�?'~���'.��p�-.4$�R���9����v���׏\<l?�����z��z�7���&TQ�L�r�q*ܡ�sr��]dpB�������'L�e4{ۇwn�ci[�AZ��H���A�re��i#��o4D�n��0�FwRύTYX�+�S=�o2z��tN/�L�|�ʹ�$�������0����\R��ּU{�b>z���>�����v�<HY�$�a�I��%P#9(RS��?�HJ����$�V�Zο��0K���W�.��A��GR�� ��&�U��d����֫ �Wf��(�uԲ�������V�:y��6�y;-A�PDQւP1N�&�o������b�om9�"��&���?)kK,{�=�kײ�Ds����R���=G1�ڄ�1a��6��GJ;��@�[o�s�A⬷�?���콉�庎 F(뾥���/��y����{y�R�I� P�Φ�J�[y$�;Al$�Q�Նq��ζ"t�W\ّ��M Z��B	��-B*V���K��)��)��"B}eeC>vV�k��,��mص���k�
��M#����q��s��m�J-T�,9��f���,_c������[%|��h�DW��򾭈�W��AK��jBU�Y�^#\�mV>؉G|���(�f��<�J�\!9�%T�<|`�sX5��ٹ"�a�u�|T�ժ���PJ�\�����/�miJҞ�`M����7�F#����x��V�Boϟ����۲��K����F���$�����o��ˇ�^��*�P#"�f8��n���W��Ŏ�7Կ{�vo=��ܱ��&Y9nf��rؕѷ �S����A�*�8�[521�n�S�!����e �F#Iq�0�/���k��
�-u�a������[߭���%Uf�K=@��NBHR����UÊGJP���y�0SR��m^,.���"W�"<�Ȭ�P\[��C���W�����W|0�d5q@k�ߺ���J�j�2�
�Q�,����d$[x� ��X�F��y�B�C<
I
�����"��:R��'���v�z,�n�A}w�U4q
���F�X�l=�4��r�6yT��rS}�.�k�e$Ɨ���
⯥���=%�˭���}�B�}��2<!��v �(����	?���{���TCMb��|�u6{�S�� ��@��=�;������j6KX[/Գ`Y�+B3[���_ OA?vMA�2ۄ�^ߖ���:�t���t�Ϛ� Q�- <��d���qd�p������dh�AE\�@d7ǘ�2A^�Jd'�k����=m{�x�A�=��$��埼��m2RH���;��u��=.��SG3wv��"N+9�*7l�`;{jJ��W��P�rU��*pa�@?�:=�O񄇢���D�=)�U��d������3��/� ���01i9�1$g���R�ÿ���W��#$#/v�I����%���
����x����$F��ʨ]+�lt�LH�:�d�PbU��<G�j"��/����U���q��s�З��|��-��M��\Ŗ���Z�O3V�XoŦ����K��Jǉ޶������ќ�Z��->�I��Z� �^�tΨ����|p�j�~�|�R֢ �̺��P(*�b[�K�:�Џ�����x%����>�6:���M�ߛ9�Uqٔq����G��x�H�>>Ɨ`�t�%�s?0��+hwB�n�9�{4`��@���￠l��/� u�-�B�&3���`�O�����hvJ}��c�j���m��j��_�� ��/�$e��|�hE>��\�&b����
�r�몒�ҧ�pٺ��^H0]w�2���������T�T��92;��5*�lD/�P�^�Ψ@[\Ɍ<v� �<�M%�	�?��n;9�r|M(�<��JL�� p�~[zE%�Ƈ��I����4�X�$wӉ���E�R��V���Y�FO��v{�369{^����N�\t��7�n(��}���W�X����A+ם�X���Q�W*w��݀V�k��/M)�ND�y�-Y#/C��y%~���R(��e��h�Z(Ӵhʪ�x�ݢ睵��-mA��/Z悮R��r�F���ſD����z��=�5�$#*�3A�c."s&%bK�;����6L�5�˃0`g���BL���g� '����y�&޷^������V�`S=�Y��rjŎ�4`��^��G�nW�Y  ��IDATsP!r�����2��a�#�9C��bYZ����?���$-�iyZ��E��d����h�yW�U���I�^�|n+A>����Y��-��h�6LY�q�}1+d�ݬ�A��97�C��5�G��ʃ�[,9�}֮)+eP��^c[j���۷���RX��]�W��U���7�O{k@X�+T��5���\WN�w�Fq$(!��n��[G�Ϻ�1�XH�1�h�1�k]Q$UB��W��� ��N��0�:;���U���8(������AvFa�1�|�\�]�Y���R��6�������3�(g��/T��:���=pޠ$�~ZWaH
>��_E����W��x�#����|��)����|��||Q���ǯEE|�WG�V�(��'}Ba>�������͉�&���u����5�о��8�+U�s�0K�+����	Ώ+�A�����Za%������B��mYo=�ǭ������d7Y�����G�U��E��&g�����P&����|룛���Ǐ��oI?��g������^���憏m\�Vo��CsHP+�+�)%�KI����:I�i���VKj���^�aح�4#��KVh6����~����3���߿�:��@ј�:R!�3{s�Q�`����;E�CS�m*~��bõ���}wxW,����V�WA�W����s�ˤw�0R�1�V��k��Ĕb�Be�O�����n�����e��\�Pޥ�/�9�g�{å7��Gՠ
~uW�c�	�5�%�P��ҝ;Ŭ��_MR0�M����"��˥��~%���4��{�/_�ߴ��*�*6���i[=Z�ǿ���#��76���n�7a�6i����e�'̮���������}s������]�qCmyr�݄����Q��M��	a��	]�>P�5����Q3L�`mi��v[	���3�_!���/i���ݔ��&�J�������:6�+#�J�8��߶���24U4&Iݫ�V���U���P���MX�4���ۗ�ߔ�:�?�X�(���/#[����ߪ4�/ى�?�%����5}���,X5[@)r�
�	�LW}���>"/��s�� �}{^Ȩ�ۢ��H��Ť�'�Jٜ����O�S����ˏ���v,8=�����z���:��M�v���{Dr�w�|���K+H<���i���{u�'�_@
8�pf����ȱ1ܛP���&��\�9���Y�7�/�he��c{��4V}:ϳBt'P��;kKٮ�2���>ѿt>k��~`i��m����(�d�/	��(����Z1�
���W�-,�z��X�����ǿ�-}�?o8���>e�
Њ��a��g�&�ƣs���Z�+<�u����Ú��g$+K�'P�"歭Y/����ͫ��f�H�Gk^�4o5֢�����.���K�?��-k��������R����/e��!�2\��W�h�W\R�{<���m��Y�.�ո�&l�Pe���Xu��hB:�)���1q�_����/�iTa<�x�,�9�}5��{�k�}O��4u��q�y���~�K(HV���+ �L��J�%����. �`!{NN&���B�[���c[9�Q/�@ޏ�.���� }6� �ަ�%��޷�,m���J�]j}��U���������D��(�S?�o��d1�n��'٠�G�h�ᖈ`Z$Q�G> �Y�ܶ������*�*�Y-�k�U��
���&�P6���� E؄g���qAl@t	T)U����-cKv���5�g��d'cM��i�p�(Gݘ� r�pgi5[Z�Ǚ��b��V���_�~@��2Xˊ	�[�-�N!��.m%ڭ@! �^����]wD8շ���+�����B+��@m��Y�z+Y^e��,�3~��Mn�+�c%m /�k~�5�@iR<�ТX��n$��j%k�$_�����o�<cB�x�fN�v��_.� ��ݍ��WQ��5��u���=����v��zĲX�c��[Z��t�M��w��oSA� �jX�@L���T�.��T=�8�b�y�BP?�znm^�r�m����]Ekr�-�g++� ���4�+�����xW�~"
���+ڬ���C't���5�g\Rr�\�V��~d��x��l�A��#!W+�E�����e������K1d��5�۸j�2P��V|;�g84��W������,Fܣo����أ�:�E��
N�lɠ�!)�I�}�X�w��MC��O���^exg���J�l�ؗ;JK��2�h���:�y��3}f/17=�V�I�ڢ�tJ�V��֞�4��۬l<���˴���;�<9	v�����*�����QP�]TԽ��d�R���zH)�~hn����+0�<,6�,t��GRK/�����PJ� c=�'+ɷ(��J��A5���n��S�g6��
�Ϫ�Y���R۫ϫ@)�B�����zU>%w��b%�]EY���jH[�JA���:4|Ъ(��G��y8N��n٩��6���i�)3-y�q���뻧�ᮄs�Jܼ5���eg�2�`e�j*wcj%:+����4�5,��`cZ,�~]C�ƙ� Y]څ���G���?��$��p��M��!�=��d%N��f�'_��޷'4�I��S�6 {�*$�߃#����'��O��1�U��M�_ N@��Ȉxʑr]��2]��%�/�����NǱf���^�#z~1�ޏ�H��~��$�/�M#��z%d�Lb)��^�Sv����
�KM�"�H�/���b*^,��`�i��\�7f��-�*s��uui�{[,G4=$ɸ_���"ׯ0��	�Q(?˦�(.">�Re@w��/��J� 	A�����JW�T�^���Ɠ�_��sD@�k�m�l�n�,N�=����:w�xd��"��!�$x�%ZI�s��^��1�C<1�G�B?�&~���mML�XF��˖�?+�K�^<T+S��cR���u`t��7ݡy��4s���!��Tn�⭞k�?oUYɲh��{�j����\RA��o�� ]N�Xۑ�Y�QF�En�Wd�sI���l�6a���g.�3h־�1��X��P��[��׺t[	b��n�|'��Y�	�����	F�q��J{5�4RP-�eP3�?tQ�8�$��;l F@��E�l>R�j��V11m�~�)��,N8O/�B�V�HE��F7���X�8Vçn!��!��B��]�QSZ)>���W��[Az�0F�&Q��5u��w�ox-<R�z���ݴ�,��L��	��5����c1�E�K��]7�S���Go�`�z��lυ"(:�V��v��^��E�G�EK-t�����֋���!�c3=�W�:�uN�˷���^΁a��C�L<��T�R})�_ĶZ)&�)e
����̠mc�V`�҉��#]���&|��=�Km�Kh������i)�Y�[5����ޡ3��O�`E|�?��ǖ�s(7�N��Z�Z}NC�:Π)��b�/� Y+�gWU�	j��Ni��/291�(x|�<u�`�ؠB�p�������?���AI�c��V	:zA��]��br��X�����)Eɭ�\Z�pU㊬�~Q3��^kgu�(�N���&�
��+�~��ːF�� ��hE�ս7��Q�i5USw��r'9}�hB�e��y�4�N�����ı���uGwLn|OY�c����Et'�c�,bq�W��Ƥ+���}9�[��5#�6z<
���
���ͫ��Y]_A:���|�����w�:�5��a�)��	��u�Si��Կ�J�+��Tc�ԇ]������:Gu=��q	Ș�����wQ�(�����?Aq���ώ��w����ӥFcJ����L�sê��v�D�>9��Z������)�F�=\%Rj�_[��l}����	N��A�n)G3J���W!�%���t�3mtQ�Q����^U�'�2���?��U��
}�0�	�������W�������L�u��w�{F�1kcj�����^�=C�]@z3�2�$�BO(r�p�]��*ꘃK3�A����>��) k&}>�M���@g,��D#�]�+�E+���y@|+��䫀�����W�W*�A�
��#����ѱ�T�����=�(�R�vo�;+N��v�#�#,���P� U�v��l8`7~uqn����z��ߓ5<���\PA�>��w�n����F"D�(jhN�5���į���N��Ȼ
F"����V�����AC�v�܄QLi��}����Hk��a�)IHkq$�(���<���F'��6xTD�!;i���sy�j,W`�q�;�l8ԉ�.�����F��\�Z~������LĂm�S:/��\�a�C�}�ݛ�K(K*oM�f�է�����Q'����O��30hp�>z]2V���
���P|��dX�kp��9)�n��@�;�Zc-�D����Pُ���N�:�)w#ό��O��&1�J��V�=NVZ�ls{�n�ڮGn�lF�̎ˣ=i�ÔԊC��"N<�k�<�%Uvя}��s�Z���>��s�L�S���0��S���b��$N����f��O��Nk/6��Ėڸ`E��Z��݊�eX�����[\�@ծ��l�\��2)<H�>���'I�E�v��m�����{ ��� �s+CU'a148�lX�7膽��3�dm2Ro�� u����D�Q=��r�\9�µ�����|��W�J'M�n �?����.�_��4��y]e[v1;Z�}�S`�vI�ky�L�*�Vr>^7�v���n�k@j�u}G�.��w��4��i��?�o�W�*�lP|?����S�f`�Y}�X��)�rQ�B��ǚ&-���@֏��3 �#�I�7d�K�-�����@^�mͩ&.p���%_ �2���Iaܻ�J�/��&9����;x���>�o���ƹ �6�>Mw�^],��E�\�J�N�.?�a}�rn��}��:�Vݵ��v�;\�F�����O9��)W1��C����s�(@
d�:���J����5�9[�(&�UQ��WQ:�Z]�-�@���$�p�4�)*��մ��� w�I��hO����,�����kMB�p���+F#bw��d�~�t����iueP%�LimL�
�p��j*]�3������R�k��Ȉ�@V7Q7��Tm��Uy�<��S��1�x^?�d*�^`�&6�ЪI���8��#�B�B�J$�7QfapȯR���!�(S�?Eգ��:m���.�0�G�b�:�#��p3!��^�m����	vS���-��-�p��T���y\h���DV�Ҕ���I4��)��w���{�mh&<�c>T*��2����^]���	�U�c[$�|�0��.���DƑ�_A��R]!���o� �����*�C
qy�*�a�g��8xd
=e���
�9��THHrk�=��~ǀθ3p�}~gAwc����a���j�*z3[?<f��n?�(��&�џle�UپL��K��y��;C���iN�_n�)�ĸ�M�CʐI>���׏��Ya��Z7���PJݼ7�â��)3�OӁ3v�T+.�宩�#������*�;V�C}C�++G��	Z�U��y9�:+Zb\�!�
`��H���a���'�r
R&� v��x���PwޭpHq�&1�� ��yd�!�|��sI�s�YB��`���v��=G�R�ЋN�z�������O�؅[�m�Mz*���L̉�Í5��d�����P�i۹9�j����J��K<|��.�T��r�x�{��8�����쎺���jV@z�]�3c�uE�A`i(�@|���H0Vr��S�-JU��:3]9��-ܿ�rD�"��_���3�ߩ_^PA*�iC�Oq6H�Y����{�pQw�����l�3����7�<�ݝ�P8&?�DKf@��Y3��ɳN���̄�߳�x�9�JMi�=bJj�|�������R~��-S�̛Ή���L!d��a�Q��;���^�0%�?�VgB[� �CFBeS�(O��)�Atq�Lᔟ�DV�uu�d	2��e	<U��7 a]ϯr,����R�$��:Fu�`?Ms��0�(�K3��6��K�p��-U���ڕ9Z�?�j�wDY|KMං�K}kU�۠Z�I��7J%r��;�2�̓�B�r���Xo�9oo��C����LP�ʱ�q�yE�8R_��Yy��Ӎ3�߷����㷀�K*H�B.����g���ʂ�O�`X�Q�A�U�o���8���X�T���-ɸJe⅚��j���$�̬�j����)
�n۝��p�����Kٟ�$T�����]}� ,��LC`e�� X�WJ=��W���k;�5��V���};xG'	�����[�D��&�E������H~G�����v��c��v"
~S����N(��7���F�
;���iH�_��1�|T�wd�n�*w�R�G�(3 �G�`�^0?^�vuII�$u�n=>I^���G.�y��6��"��|�P"%�M�x���*L-O֓�Y�u��L��Q�p��%�SR�K��av�>�v��Å�� }��ǧ
v_�:��G���C7��0��%f���6 �(ߏ�Y�e��pY��F
fn��J��oD=\�����aNw�#uJ��(y )Q��ty��v�@h0��mO��^++5�GQ�#���k:&� .� i���p���x����>�@�\����a�ﲵ~�� ��>����Y�|Qro����7qx:������:��}��-�4922��`�����|i���W"<46&�[h8�H����7�ɚ��9�~��21Ƿ�|x<�{+�.����i��b���/��һڞ9��]c�k�
�pa^}���Pa^[{Р�Qd���{�F+�:!h�Lyg�4b=*��W<���:*T��m��[����+0G�8�ҺW��M���J`=+��2ե���<�,a~%��}�����D�������c�rNh�zow�,K���Έ�^)(���KO��?o7��l��y�<$f����]��0��t}Уp��`J��~|����\RA�>����R"6���
9H7Lc��t�����
����+M���c�]�Ԭ�����|_��w��@��,�o&�#16h�������`�X�Qق �`ܙ��e� ��{j��`�Y��Voi�����x��![�� -=�-��[Y�w���@���D�O(�D[Ϝ�2�n��&���Q��O�85�r��W�X�*dݬ�k������. ��;u�O ÞC��s���T>A�\,��}��Z@�B��ֶhe/?�����K�[���U9�<���
�>*1�wkv�b��u:�+������0���X��I��-xG��
vF�)��t��(��w���xM���g �����,����f�Cb6�i:���pW������9��T���Be��'C	�%�"��w�ڌbv�< ~���g���P��d�'�]yMI�'��V"Z���gm���XJ#g��`�o{F�ਏt�X����/��h�O����O�H����o�iI|e�uE��=��1�\�{8���
}��9<�>ڙ@E�_ ��j�^P�Ŷ�6�w�����$[M���&�����qL�:st �g�J ��IH�ƥц�#+w��*H��>�O��%�ԃ�Y����L��Cw{�^Z�G�x��r`��gΎ���_7W]oc��p )��h����wMa��-�~c�aWF��]�I���%�0�!#��
�	�ޞG��׺�g��Mr�,�O����/��SZ���k�7&<��.� ���^�e)J�s�ov��!���o���Q.j�z�B����7��#�f�خ�ʕ�}7\zvJLH첫��_�d�a�hi��*i'w0`��u iؐ�����d����G��Y������5.)Oͨ.m�����#D���bh5>v)�����qlCf�$NT;<ЏɀtE���2��j������!o��2��3�N��l!L߸3�[e���N��o��� � ���3��[!O�$6������w<�Z�_��E
� au>&�5GJRS���!	���o�ܣ�4�(%�xt�>6�P�dh=�ٙ�a��?;^�rx��̨������� ��X���U9��$$k���*�͝]y�K��k�g���t��o�0_H������0�2_�R��r����l�me%���ϊ�G܃�,�e%��	̏�Br��	�������R�4X�P����X~�ǁ������z��5T%_1��l��ߗ8�%es�8��o�(�oJZs�Sۻ~~=8NA@h�Ia�g���W������yR;ʺd��Nd^�YZ1*T�������1ϰ&����s�p�'��P����|�Y�1���+��0Zz�)[���7�턻�ܠ/h�^?1�C{-<R�#uJ#Ԅ�0�UN(�Ic�Z���]d44.����	�)�E��̋ո�(J#m #�ZA�6#����]..��:�(���Ŗ�*�eAA�w��S���b��t����	�(/����h�߫G�p�%��bR�գ�:dz'{����W�穋0U�ȗ�paP�� 	d�s��a�}#-�
�{�*|	В�08%���n�u՟X�ǻ�>�@���&��5Ḷ�⽭(U[�0��@`/�����*ִ�zUtL�Jgo���%���g�<{������@0��P�^OA��w\}v��f���� le�K]�q��߅J҅���vi4��R؂_
��E����-�阹�Fy�t��}/ �$~�V0�:/��|�g�#�ps_ʸ���w�%#;�Ԭ��N��)���N�����U���D�*�mx,��s$��7)�����c�ڴ4�P����'�ʈ�����o�!�L�H��ׯ���m,�����UR�[�I�m�$J��޽�tY���;k��Kp��"�2ʛ|���0����	�=���X��J$��]U;�����	.�.=�q%�%���p�7kro�����V�
�7�+m^���������o+-�B�2V/��>z�/z�OtY�A���,h��x�C�!�Z�(2�V�<�M"�ZjK��Ot2�U�@��Y��j4c����L�)@*�0*[��+�\�A��YBNH��"L	~?
)��� ���{����H����;��Bo^OA"bS��X�9��H����� ��RS�S�1.'~�b;_~(H�wmЋ��9���@�����<A4���\�����.Lw$�#��������#�w"�,�����pk$v+5cE�Ke�-�<DJ�RP�AfKs}O�&��ʬ&�n�e�!���5�ʑ��� �N=���kK�S�2��~(�������|�(ג�{pVq�g���Z<
��d"�挭����/� ���k
���W���Am1yJ��F�#�����
x){w�����Ж�ԾuZ�$:�K�#f`�Y�j�t��m����T�c8W"�=h}�_�׽h�ɢD�=�|/iG������:ɭ�uZ3oN���!ၤ�)���Ld ]Z2-�cY�ږe���^����-�|^kݱx�l��r���j�}�1�^�xmۋ-�9��IW�����NA %x W6�1���
3������c�v�Ft'�;K[xU���kzd\pn5p�g���#H\B���T������3�V���L���9�V���MT�fܘ�<��&�SW���Y\�n�{�ajH6�����o�[��nůAwP�E�Cñ���$��NfA�t��@�ܧ�"0�c[Z�֘9��/<`/����,AW�$��s�%<Tg��].J��N�*G^��ⳇ�)��D� c�a�ю��ݫ���@3��V�!eL�N������ȩ}?�y�m�#����p���Τ�������;���X����,�5Ѭ)K����2�[�!��o%�i�]�˶@W�V��&��;Oq:�3�ݓ�-'���� \NA"<f����@�t��s��.���}2�hrhi���y��J�+w�C"wڥ=�q�wa8�s徬ͱ��Þr������U1�=_�T�s�~<�ʵw�٣�֣�8���U����xە"-��$[C�
ņ��k�e:�x'�F�HRu
��U%a|�0�r0_S��K����5�%=L�y \NA"��0N\ğ*�P|�.�wx� �� ���o�N�&Z)ĄכkZ{�R�Ҍ�t�9�d�1��e���P���"�f�D=�f���J���ߊ�{3�{�H=���%��k ��#�g��!9�xn��j��W��J�Ұk�ƞ����b̶�݅˸���I���bR.D��T����U�S��Ä�����*H.��#�\�y�O����dxl��;$D�mK����ƾ��^I�!�χR&#\t�Y��l��Us��k����MU���t��	V��=Y4@������] �����+���!�"5H)N�'c���P�":�,��5ɝ��Քo\{~/��WW>e0n˚��iYᑶ���y����X�?�4�|���䣽��>�d_J�t>�7�Z��o{�h/N{?�����H��C���o�������+�� ��Wb�0��>X3���|u2��JC����Ԧ%�ؑ��K������3��hT�]4%j���}ë@�
^F�p=��ө9G���e�:��zQUX����z�EZ�G..��6����e�喝���RT�]jש�5�fD������lڮ�9��H�m����V�b]s~���r��
��0���Ey��Gh ��M+׿�X·%��g�>	z�&]��H-I9�m�6L-Q���;p.v�tz�;��,AIy�dκ�Uu���mݲۺ�]�ܼ�9up�q;21wV��|�Ҡ�:��Uj�ׇ����d8u�X��E�B ��������\�����V�!8^9ߋ�g��܃Q=�DЧ������Dy��v9�dA��[+'��ځr��.�-0۹�m|����d�"��Y���g�= �t�4��x�HT5������B�I���7g;zp/��!�����-�=&�}j>\��_SA��Ȕ]E��y��/������<���.��.,M��.
�ݑCc؃���_`*
�����K��4���R�f��3+�3�e����_q�"61���Vq��8�MN�_�w�����r�-�D�����I*��!��<��б��2��lź���VAII��:A�9�g���lh_Ѻ�� �;"�hn�~D��9��t�]Ɩ.q�U���3�m/��yk_0�?��P�}��?���dCz��^(��2Z��ִ���tW�1���1	�)�sdH_��?vX��p�ʠl,S :�}ζ�� טoYc1*�^:�q�*�H�D�@pE�4҈��v��w]6{����P*�q��
z������-T�RhXx�@�ë�
Rs=yHIB#P=f2�� t�u���Z��_I�d˧-�HA���}q�Z�+�)��=x��nƚ��r�0����)G�^(_V��ߞЫ#G�����z����O��fw��C�d��1p߳���i��(�z!�^��3l��1�9�������?S��{ٙ��-��m��V��۶I�I��(���ڑE��Dq�<���xKCЇ:��\���6V��;���$�J�s,�Y��G@zv*K��`�jN?V�(�P	Q���g�==�;�%L����_�N.����c����7�X\�l������Hس���oz!�i���r�	-�:�ڥ��h	+�>�}�[A��RS�H�;5�@�ձ�E�81���ߜq��L�@�Q���%%����"ȝ"����s��5;d�@Yuڑ����>^�DH���}��C*� D���{��1��-�膬���ekXw|P}��@o �JN~��yin�x}Ok��l�,�V��.����< W�^9�ghP�zJ�#B1	�9�_�?���k5�U��2�-�R�$Y:N����z
�;�ę�kd��eׯʘ��ï�x�����΍�=��4T)>��__΃�͞ȫGmN(vi�KM�ϧ	(�9�zoDig*=Ů�X���ǿ"&��$Փv�U�ӕ��$.��shx�T�{J/��ݺ��<\�"�HG`�Ǧr{�I�ۓ���ઽ�Y#�����#F��h�Mm�K%0�.� ����`���o��=��`�N��������1���I(�g�5ge`X���h��c�[� �?`��W���"��}�pr��� o�滰m���}��l��UQ��la�.�N���=\����Amdp/�Է���r���K�ɝ�&JO�Q��(4�@���&��:�h�b��7�8��c*��3iğ�y7���=u��ml���o5�>��=/������ԍF��qJ<6� ���5q�=U��xB��Ů�l�HQ�M9�D��7�09L<� 8��N��ǀ�̃K��(��҄���n�vvq���W�n���Tv�]\�)r�xD��Y���r�׎F���N����qI�e!���������v)�UY{����\=�䞶��"��ţ����,�3N����#z�����ᚂ��1rJ(?�[/L,/� 5(�HC~ r�\��=[����us�|��v=pb��-vQ}L;�[�f���W�V���[�V;U���|Si&Q��Â:�((Yt}�^�q�'��8�ab����b���3����K�_ۀM�;�(gS�]<�Kls��r�\�iN^�^�x���^�/��x�O�V�E\�:S�4/����zgArZy��&/��6@�ޭM𦌞�y��P��WI��s�M�F���מ�c@�W�d2��n�jW�޽k��
R��>��8+�3�lЍ��ϳ�sBTd��-�r���&j�eT��,��xg�9�j��g�z�XAۿ��a�\fp�#^�0��"�i�X*j�u���c�}e��֩*O}��,e�����s8{/���6�nw�?���:3�Ǡ�5+ƪ��5�M0	�{\�+	f8�x��sܾ��Ǡ�d���qM�e�4����������<�̶���9b�ސ�	g�GeQ^�.$^9�V�����,ߞ+��l��~�uXy�`�~��]���$aݣ%�-
@�h�Od$���2��P@�����ʑ��|�Z�!^��=}��"P���P��嶝C���Mg�Q�E��BJ����b#� ���FE.A~Qa2���r\v�Jm_QP]	���!�dV���>�[YO��6(�%��3U�#�H/��t����1J\�*���&2�\��
�@+�Ra���d�휊Kk���mj6����潂�1�ψ�x�*���Nϫ������x��g�HT����h��Y�qR������A-��w��᠂Z{��|�76��^�Sv����=���PXf۩q����8:��ײ�V��A�]�F�}�$rT�
������!�Oo�FE��l8�V=��w`x�'��f�4���(y�=��9��ɰ��V�M���Vx_���ڽ�%E�#����"����5N���e����(0?Ɲ�p�{��Ӝ!��6IX7�a�~tt�z�k�ُ� YΕ�%�e;y�@0o���x$Eq�$��S�����f7��U��@�XO�7I œgҪ�'S6G�<������^����/�R+8)Y���|�d�|�����=����
ĭ0��2�nZ7�֢b*H��L�s����-+������+����V�U���/%�V���b`pi�h��	z�%�ͩ��/	�V�+1���i���"�5�"��p[��k�ѡh[��]�sC���y[�䊖{7�$���(d�����;E���R<�ǟw���*��X4\HWd��*H0�b�7F� �*W!/L��{`x@��#B� ���� x����6����X"�{
j$	=E�p:�%�ʌȩ9�F���ZZ��w��CXO�ĩ(q�x�6R�S5��1\ ѐy��d�In����w���bw��x�ޡ�%hqfk7��.��e��$���o�a����x�
�+��ؠpJ�������?/��*�|	�uAo������iyK���d�1���ʷH�Y��lNDNO^k@Է��P]���6Y��~���
s��	p�Ph�U��=��R��$7�;�����ǁ��$q�g��Q�L�(���/� 5`K�
���1�h���
�P�RJ�i��˅�
� d�Y��\��>�&��'�e'�E���q���T��$���ě�{P�,uG(�3Ì
N�Iܷ�E�7pDV��H��vL���c�=GϹ�zOa>��C��!4aeD���%�
�a�e��J��V��q�Z��+|GE�B��p1!�S�X_0:~W�al@��6!Ȱ�n+���:�И��{��z����-Ч��%��W����W�b:"�r�v�+�2"s� ���*]&dw%�:�Ӭy�b��.9@_3`����T<N?R>�"�9��>j���?�4^<F_��ٗV�vaG�{V9`^2%}>�a��z�^���?*b��>O��;0�5�� ��ݐ�����>o5�x��1�%jھ^�A�����xVp���Q�nXHrBz��SU�6�5	��4� * ݃�ߗ�S�olx����X�t���qxa�2�qQk���n��:5a|t�*���pˌ
���2V=��| �GO���;z��bʽpQIX12�[��-����b�eV	G���X�^]xUs:�����˴\�'؅h���;0�8�8s�AP��4[Ѻ*U�{�D��),�H��~�W�X�`���ꮪ���Վ�0���B#�RǌU�	��<��X��BwX��G��ytq���̢����^�����7s{��T>AX8	�S�@Y�=�o�$��d��L#�S<�*�P��G�C[�E���z�*D��D���zPB\�V׵=O���2�g��:�Cۢ�X�h47;�@������4h��#?&���*�o���N�<	4m̨5�TV�)rE�����涡G.ivA���������+"zX=����X^*[�Z����^��
����T?Ѥԁ��ܧz��l������	�jOx�l��O�Y����oBXH_'q����	�8��`�>�q���q�`a�:�U���s��\Kk_~XӬ�^<��ц�o�E�%�F�~k]�e��ASF�|z�ƩyU�9���/UT�Hc���`�l�4����J�ì�	��<�?\!��Ϯ�t����6�uҁ�w����m������=$���ǥ�y+���n߹�~_��[�{T�6Sf�+	�0�r���^��k��
��c�\��*cq��^pB@!�i���s��\1
�/giD��������zt�~�jd��OA��#���@σӀ�{�c����:�1{�K*Pi���E�=d���=�wp����O;�V�B�)����d�.`N's7�P`U�x�x4�N���f�˕�U�ik
MD9���ފ��:�v �
��sL��8G�l"p��*�u�Y�∉��Os��=@ـ�TɃgpc��� ��K��^)�髢��:�-���,������p|��#�ݎ} �9q��ߋ���멠i<�t��U>ܥǌ
��L�5=4�r��im��-�[�3!|\RA�gO�(��.v��9+�<��{�mŎk���֍���啄0+7__N3*��ɩ$&ɏ�gĝ��Ŭ�@"6��,C�����Mv������)��$G�R�G^��H����
��IM� =L��8��/'H$��q�u�ʢF3ފ�}<>|N��s�
�Og;±Q���6e�K?�o~�|���|2�ޝ*��U91#�*�nz��3�[�T�8a�U%��z��y��~K� l4�X_@�L�����9䎘�?	����>����v��3\RA:$�=j����k�捒��hj�y�����|weC�_Q�}V�N�����M.���\�����@�����r��K
}�PGW��#�ˣ?�J���6%鬴,���#pMq������^y��nF����*� +x��V\����5�)���ڕ���й�G[��H����`\xX��ڛb2�����.�\Opq��:	�5�1�L�"�"�$������o��'�� R�i�A8��O����(�����w�[�zZ2!��e��z�Y�T��mÃ�f�#cG��o6��
��#�B�r���X.����E�0��7��mi�<޼����6F�9��P� f�V.���X6����l��j�[�跹(|��fPrdq�����ҍY���L�&�� ��}��WZ�$�Z)�7��<�3��9ʳ�k�ݍa��
JI��i��3�[�(wk��l8�T>����R�B9W�@)=L�I���5�8�4*y
�.E�9E�k��M2���p徛�C��2}�����L5F�S_�1�H�ް��[V{�A���+����ȢQ��WL~�+�bW�������-pM�8O�{[?�]��F,v��?��`�?�Y�^�q~�	������d3A���ɏdЦ��U�H�YӜ�C�q^
�f�X�i�:��!��50ٵ�q}����K Yyu}�ez3���.�}1K Y&���31>D�`�iմN?G��3B�{\�8��$8�kV�ųc��Z��0�<���o�����iM\���2:[�*e�(A���\��TX�M�(���Z���p�	F'�e��%�d4%x���C��)��ؽ�X�OwB㌄�ڦ�b%x��}M��I�9! �	���Jy�� ����u��ǩ .�H����$���xV���{�t1���m�����J�Yʜv���5��t�U%���7����ΗT�8�����)�"�͢��KcC_Z:5�N���@�{<i�'�(�]��#��.
�U9ef�mp���])��p'N��Fj�/ox���Š��o�jtX�240T:-�p-�� �qB�ӌAf#�u�
R��/,�"-[O]#���J���ʎ)�S�Z�h6������N��������J�ϛ:�n����������v1�x�4N���H.	ܠOSO�t�^�Y�$z�]r5���_<��]�G������LK�:�A_t��/��~l���[��B>wK�����
מLؾ�b�K%y��x�Q`��w�7{j�9P�.�S��&�G�5$$6�����H� �X<�М����x �m�[��M �UX�C�U&��{�c��d	B# R�}���
���s��3,�2d�X�e��K�7���+�� �6 ��#!�i�ϭ]�dI��$�v̌1(�C��e~��+m���bs�JyMC�?v�$o�t�s��M�|"�`�S�Lr���ҭ��)Xa!����4;��}�M��EH]��y9�x(Wb�]FB=I��'|�]� a�u�.���AU��;�Y�Z�ѝ����KP~��̏���5�j��QT��)r�%�o�3���;�G�"
v�L���pII�T��%�(?i�I���0�I
��q�7U�}5�.��y\x�@�E?�	�m��)�%a�"��(N����T6�V0 '���� &���Ê�T��y�j��r��8*4E�=#̰�]�a�}��3�k�*<h ��4�9eR��*l�'0���۰##IR��Ƙ 2tF�c�]�9Ϋ%�ꝑ7:|�9�Zݫ����o�mW7�����b���z�tx�^��Xu�N8p�$z�����W/���>u��C<W�$�y�U�d��Rz]��
RCj0��m �=IZ+��~E�u�8bHG๨�PM1Y�w���MV֒�����<p=q�������ZM��~C��L*F�!oC�זA2v�s�N3�H5&Av��_؛���^�
�q���e�mà묾��S�틕��`{���_�I�S
��=r�����#E0i^4�s9XA�zwǴ��[7��m�I�ֲ�Ɍf�"Ep%������ [�J�G|>�8�#O�,?��6hË^v&OoŲ�.:����J׽=[2�A��]�~�Kˑ~Y���膙�Ȯ 35T��E8R���'�cX-O�<�u9�x�"	�D�d'���O�� @r�¬B⛎�70�9���=X8@w���F�G��I�8R�W[�9|�w��P�9�c�~�&�#�cY��aq����L�S�� ���0�)�3�d�p;uX��֥��:�|V�	��a�}k��^� ��n)jt,����t��ZMe��Q׏ae*���@��c:5�΄�]R"!�)�+���k��ø���S���z�*� � �0��X��+��D"V�����FD�8� ��.X-R���y㳗�r�J$b[�ה�e�}�������G�сJ�Ŋ�|��kS���/��.� e����	#H���?;T�&�����D[�(<P����x���#7��MD<W��b&>�ϼ�W0��g�@X(U14����Ԅ�@([雱�d�{}^�1!d�,�{|��k��M��nYs0y�~�w�=�>*˸ۿ\�>�7I˼��QHߒU���JŠ^���|��U���n}#��N]����/u��䲤}le`�eu4��~"��}�Dq$OP(c�ah�T��QZ(�	�r��UsA�����bզd�}�����,�_5���`>p�W�ࡤ�PW���ќ��,˒ֵ]�L��e˼:K��K�7�L�N���j�!H��?y�r�!#X����쐎<��e~L�F�E*��9�7�[���^��xx��c"r�g�)��)lm�XZV �z�]���K���]�E�;�fjS ؽ�{�����x�?�r�bj���e��y��؀����)H4��_C���»��fp�d�;���� ��~jL
�P;��1��!������4C���Q���db����/u��f���W�<�0���5����Yq��l,{xEbĭo�	�C%�Q}�ey���<~;u��'N��H���RPwxq�)9�e��؉��U�Ⱥ��I`q�,P-�> -`�8a{��8��9=vQ�]!��-20=!��TbO@A'T�������$�ҙ�Q��z�p�m� �9��D���y?\}����z��@�r#�]�!T4_���gK{��Q�4�o���3ؗ�f՚ap�[)KR�G�{�'����}/�\� �IN�x:<cD	��ak�V�kf^�L�]E(wo��}N�/� m��@mY�ӱ1��� ��0����:l���W�rQ��5����C!Z�
�����Mq=q�:��mWyFl��FN��"���k�������d�>�K�0|u?lM��&δ@��$�3�{��n%C���s9�QX��Xo��|���_�L��2 ��$?�6]Oh�|�P׶� O��DO[��*�D:
[��od�����!G�d�9�S�܊u����k�:��0:a����Q`�i$����)b�¯��sB���W�b�`�u��ܻ|�{JM9��H͔߃:���:��������l� y_�Iz���l���F�W}��$���͈`�|nM���d�e|iat��4���q*�f��%���~��
J�fZ8AbF�)C/�u�:ȐNX��y����T��%����%(� �m�1�3�t��Xv����"�X����e�&���;�������m�g�-N,��(����f���H��L����[�gW	��@�[_���%P]��C�� ��I��k"��qsJ!�&�y��b���	�wX�e�i�<�4.]ͪT�	��9Z���ҽ;�*g���p�Y!-h��#����ŏx�zP�-M��Ȑ� ����hۘ�5�����m �T��1\�g��i��>������f*�;a9?A�x��T���Zݢ�����5��]�D�j#Y�L����������D[�]�%���5,+ ��*�A�,7)sE�E8\DH���'�pW��ף}e@~F��®r��K,��P��Ī��D�%N�W�E7�u��2�}"�;1��Z|l�F+�=��^^�"����a��S�c=*b���]^m���K*H�ㇸ<L p�ԥ�TԜ���!�L�Q ��Q�{	��G�^@�-�(i/�'i�108��*
K٧�(/�bL�r[ދ����!j� �2
HS݄v�ё�fۺ,�JMkj�X�ߡƔ]�y Z����)1�dm��M�$Le�R	�������M&�I�h�|�>��U���CY^m�k4���_r>��d,���)�LJ֕*���C�1�3�Lc�L��
LC���~jtJ�7R^�g��.�"^�8@}����IH���}��	����Q!�=�W�Tn�f������H	�³��c)E�r�ў}r�ۿ�]]ς�@@n���7w�Z��8������[���s���wj�U(��ؑCN5d�d��j�k}�V��֮��#�"խ�W��̸���#������	��"(�i�g��I9ד9*�.ࠕ���u�5)�5eo�/x{y5���,?Rb�0�*o��)HB�)��O��,�wzUU������LhL4�lp���1���.HO՚ݚ����x�����&t. I��z�C���������3�|$gIl:"��=��]McG|��	���w���m��!�V&J3N��,yO�g҇�IP[���`�hj�C{�L0�!�:�L��{1�����1��7ՙ�6�=�$�Wsi���*V��?�[m��a�Oi�F!�>�M��	�e<�;TD�K}d�4O��"����<vk��O��������*�tH��rf�Ҽ����caU)�L��˫Kb%qe�5GO��8�ಮ��@'�Ml���:p#ۜ��4��\�(��
�*�k����֗aċ!�K�_Ϡ���Xx6V���Z�����O���``���%i�rݙj���( ����m�5y�8��f%���b���mV;�u�~Q�O*#�P�4$��d*-WO�'r_��Y����-O�Mc�;n���dC���ް�����}b�u�������d����l�2�o���I�}�9gg�`�f���/�~�h/���x�"�|�C4x�Je��%Q�Mp9is�����������X$BK�(�L�K�4��J�0�~ ��UL�M�����S�]@�7�+x)Ȳ��Xb���K�v����#)�������k��uT�k%I�G�
s���r2�HHL���XWE��������Y��gf&?�)V	�f=�ɪCޓ�_l�E�=�+s�T�9��8C]��Vޠ �b�&Qpwb!�P�ń?~ܦ�G.�l#����11�&�Tn�-ʞP��S=(
@�b�����V����g�������s�mf��q���l�H��Buk� ��(,Hâ��>�|'���ۡ�!�7o�fЖ�5O��[~Y8Y�g�����Q�u�rME�싍�,�N;�fy�OKJKd)��6	U����2j���NZq�t�2�����SԆ[��,Є/K۵A���+�Cn��������$pփc���s�k��D��\"�Vn��.�E�y�Y>n��Аm���4�Uq*꘬ N�Q������ӶK6��m�T������6lxԭ ��S2_�Zʕ
~f��ǭ/��ٵλU��>2.�y�ZG�+�ͪ��@P_`�I�	����=�1P��>L@c�^�E[:�(�#�8�q�|cg�o�h\������.����~�����2��#��	Up�N�!u$c�/��1���SMf��$ك���q�Zh-�G����.�3)�[��m�a��2��?%���Ҧ�"V�DV�m,\�/)&��H�������9h�����'��L��g9�dq)^��l� ����3�� pq�="[,�Vj+�A"R��C!��_��.�E�g)e������f��	�ví���i��_���,cԾh,�n���C� �-G �C�-Y�+:�Y��M��y�׍���g���&|l^��%��_��>H}����{5����!�����#x�+�4f5>�H@�+ �Ig�pݖ����uɟ˟i������{��qb,Y���3@��L�9 h$w'�t���dn�G�xN	ſlo�+�������n�V��
x+Jn!+�M��ʖ7�@;�+�ᦪx�c�cO%�H�h�)����ꅕ�m�n���r��G����ֿ��M��P�{=Jo�ț0z�6�S<sR�x�F�B�j��Tn
����GJ��3+H�� ���yHIL4��e6>���H�y����`h�zUI��Z��)�Z��2j���N��1���NM��G%�ZV<�J<o����k�L�n��_�=��� mց��խDY[�����YC!rѡ4�3�����U��?���������p7�]�-�^?� �,<��l�ӟ�7Fpc ?n�����e)��|���+���]�W��鎑���8E����dh����E+
��,?�L?oL`����~���eə�Q�UqQ�x� )+�}. �74��!��H �|.��Y��c�f��U��MF��s��gV��������O��������uIf��`�˼�t�CA(���䠙2�n��*{�$��MЂ�G�����)��?*�Z��`+aM��Z����� ��P��ͩ�:Mn�S+p
�y��N�}�ʜ+}"�:ou�T$�y���y�aU��_�K�7�ƫ��ʲ_t�^��o�io���$�=�C�r�6򰧌{���U?	{���V�'�ɛ0���O���%��f��|$r�XbU�k� )��]�w�#�+�0>Hl���D��"R�*�BX��s��m��#��x��H���O7i�_R�[]ݭ�ubӶ�R�i�d�DB���~&�K�e��eueH����H�R  o�[n]�Ͽ����ۭ�>*���l�Jc��Ea\K�o"c)���ܟ~�[#\�&��W�1���#g�K�L�Lp��'�@���)a���h���g�Gz\OAڬ?�Xo�~���ۑi#��"��_��x'XK"��/A#T:�7C�m�$��+H,�Iwpu�}3��7��&�Jy��������L��m�����	�:�������*�g��G�Gj8ԗf�[��jF-��;�ޔ����L�o7��?P�1$�ͳ�^h��&��v�ǂ�y��w�r�n0D�C2_Ȋ�����JHY�@�h?s�kb����L��ςO����h��нm�xn�F8��`��¼��u�����v�{�;��	�y��ϱ�=�[w���5�xQ�iE[�O>^��NJ �~PK�L$�������|X�Te<+H���mm߶�݄������_�W��ˢ&��Nb;t���TPqxڟ\�,���U^� �$A�A�$H�,&��g?���y��}��g.��̐c�,Ou˵%�����T~���U$����N�E�y�"�u�|s��q\�٤�?�\�z�i���&�7a��0xg�ǰ�!xW��Fi��N>��.���N<r��V�or����z�$�֌���ھ��	{�*֢���z�Q�O_={Tg���i@ �N�(&�Q��)�	`Σ��t��q-�*��S�n}���ָ��ǖ�?Rw��m��H��1?BX�_�+4��Թ?���G5�hؕU�V�4}�E�VJ�}J���'�q����������p4m��(�G�"~�ʑSZ��Z]��k�Z�?u�����-O*��ⳎW�6����ے�1�J4
�,c��q�;ԵM@��zpe�!Nq;�	A��#j��ό������L��ِ����6Z÷���:�Mő]1;�ă]av.����Z�GAh�.J�mu�`��e)g6��c�H���>�2��!��0�<y�9S[r��Pz���ܭ����n|ES�Tψe��Bj�O�9
���b�*����ٜ����6�׵�L�-RV(e��փV����֫�5h�$M	ss���#t֑m����/[�����Gں�s�9!�6����y�]���~]�>+o�����*Id�+!^�p�]]!c
E*AKm?�kZJY�ضQ�M����䡍7|n��F�ȓo"�:_,��Qm��By�/�����lZ[I�[���,%���R>�#���g�e������-�!�#��%�V�B��
�E�}�LG�RAgID	��pD��~�ա�*�|D�-�Q^��TD�ϲ�V���܇Q�N���m��C�KY<��1�ڷ|�@J����H|��U�`�{|���a��A�R)�@�;o�a�k�~$'ܦC�����8	�y�>�	3!M�>�[	��-�UC�#��yz;�m���ʪ�;�� Rh�&5�%��Mx gXW��B��mh�l-�Ǫ�c��Wn���:�X��������YP�'G����ϓ��:n���Aͤ�߄�"��s1��Z�R��}������v���s3_;�E5x"���+������got����1:G#.�z��^�	c�u�a��M�kS��	�}R�[�:��I�����̤v�;�բ�J��*B����EЕ70�C';'�pc�d;��N�L�`��m����۶R�I[��N!u+/���$�n��V�<.R�*h���.-�`�Q��Ip,#6��.kV�6��)UsY�g�V�'�Ħ�A'���K�(����U���NeG� �̕7k.���aʹu�\l�����D��̨�I�X��[��ru'Q����J]!�/�	<�ˈ���B�LMY;�B���$��$�TQe��X�;���G�� !�Tw�wKl#��Y��������wF��6�S
N\��Cqb�]̒������C/w�W�W��5.��-�Nd�@��,@�.nB�BRW�_��R"(�`����,��+M��Ll={(����(�sT��<��u���BW^9]+s�v��sJĈA��QSb���
!5�����u)t39e|�zV��C8T�9 lg��>�	ե�Z�C��.
F�bu'N�&� �����i <�z���vH���R�j�5��Ua4���T]���e.RDs.��4��<K(�4q����b�� UW���.�>��L�_o�?R�hn�6s�mq?Ws찗R1�U�G�em^`���;�cR�!A��6=t��J��E,�p�r�.�q������9��bƛO�� �DyH��&�&�da��4���X��ve����D�B�%������H�Bg��"��Yr�
��<G��b��}bx�5�m�HNp�R~K?=�2��t�f��JS�p��X�'�3G�+��QG&m� k�,�� ��6��y&V���t���Ox�����4^Jb
�Fe������\dQl�76��w�%$���/����P�8�I1�+�c@��;fG�����g��@�$��GO�0i�,�0R��!��w�@�@��spXLk�&
mDߑv�PhBWG�'��QЌ�;!�D�}P�ɑ�CUD�@RI�L�Ax0J�%$�]
�І�aZY6��[�-ͰA�,���l���
V�K&XW���k�����0���I�G���d8fr���� �`�]�H�ܓ|f��s�����$bq	EM\X1l>Ƒ�U*�t.�&�m;p��٫��r�>M�r�R��
��A9G�!��_�H���k�LΖ�^�A�ʳ=�1I�)T�]҅���5�� y2��jۢ˽�m�o�Z���[ɡw����({E�2fP�={(�&a������N��xP���+E�����s�'�Z�K�8�;���|�5k�����3��$��R3�I�<#,��FxjJOxyo�iM6D*lM�5"�׫�����jp8E,�U�k��,a����S%5f�����������Fy�Y�&:�4N	�}5�4�ɞ�$ɡB`��<��ш��/�T��~K�)8��5��υ�u�x����e�.��|��w���PJ!��%���ף� ��P�k��Q?��	�P�1���z��n��*��0W�s8K-�V��= �֞��{�<F�٬)��ڧ/�����?ʎ�Z���I��Iq�����x��!��sk��eA�B��rƃ��xiB���l+�+mt��VV�%>xN��U_��+����(�j�NT��{�S�,u]ywH�/0Q?B�#9/�~%��W�Z����A��x4k�3��h	�+N�\9�������a��	.� !!xY�nV_A����p�^�NJ���0����y�'�Ǉ���T���v���)��HB�dU���+�F���F򚰬�6��y��ј�ԍ�Z&g2߸c*,�` R@H�b�,�U��@���Y ?r:xl|e:��7�ST�c_�<2ݝ�
G���֠e��t�ka��|l�U+��s�W�>B�x=�W��.Ȃ;����3%A
�(�~g9U�x����LW��qFr�nv�p�����l�6-�KKs/��.ˀ��Կ���'څ��b�]b�
g��1i��6�A|��;[׾�05Hz����s�e�ٱ����i��L�-�R;P:��;�O���;�z(�r���7�G���9����K�g'IKGdZ�8�T���mR��j�dY�x����{��n��k�ks���k۔\�xHp����[1I�;�!a6�	1�E.ؔ��*�;
HIR5�Q*,h�! �_G����v>r;�rj��Zk&ˡ�]�XճkWY9�T��X��i�WM�J_�x~c]Hg�w���KN��皀�g�>��BmG�b2�u\R�3ӭU��<�P�QL�l7Ga&DyO���18����*%���b"�wҨ�E3=����p�(��U�ag�<�ǂ��S�i�I%����R�ߪ�wh2�l>�ڑ�~�)�T�p�犷F'��^FТ����<������\"����qf���+��-pI���q����,�'����; �LG�i[�8U"�+{t�}[��]�`9e�������I�F�~ �<���Y?�s ޶K�����E5���@FI{��@S4�qósh��Wm[��C��C�ذ�i���A���"�XbWJe{N�@�Z�� ��\��I�W�n�Mt���0{X��9[
��U�g�xO�P�}��.��ĩi{���$;bqi�����ЯmE"e��5��.���Z�S���h��C�*��:^�8�IzeŤ(�li�:�ծ~x�������E��yY�E,�h�j�z��k �6U�����Y6�x8�F�|I��lԽ�Z��UC�yL���ʁ��܍�I�ep|����֮��.�`J�e+vb�%t;0C}G�%��mİr�j�����&
&ڒ�jML��Z��\jxs҇m����
���FŹ����5m6���e����D���Ue��U�Y��Q_g}���v�&S<l
�:�IBA�ܸ4�k����9��D���P��r�ȑtu��r$�cޢG�Q����U��Gb�<��V�ٵ:H=M�F��s�x�@�R���@�P?R���Z��m|&���زZ������!q@7W�7���c�hi��u��(�|[��tZ?��֘8���W����Zh�+B��j�v
V���qU��w���nO�����t�?%V��-g?gG,oc]�~u_S�	:s�d��X�[&�fMh%� 9��K�!�h\�)d�c���%�H���"��Ѣ4S(8m�J���.������[[q?Qmt�7]�||d��r��n/<�hD�gq�ɳ:��ʮ�Vwvv������
�N��	�S ?���ɟJ;PjҡNK��"�_���� ���0�����%��^����\!�P&��̈́��E# V�@�	m��
R���(=��O�^�ء&�cûNk���4KRc�^N*��#��0�5 ���⅜��'ޭR��O�ɂ$ �R9 V�t����8��]$��N�x�Sa�<Zu�B�x��a
o��U����I|�-��]���=گ,�؄��]���Eq*�I�
p��Ą��`�QQ�"����xk�F�Iۇ$N��3��z��J�ؗqӵiu*
.=�*d�(������g]�<XS:���I �8��~�I��bAɑ��a(�Do��8�pL�r�1��KS?�&`���Z&�%L|#F~0c���nOg(wI+J�/;�9��� �^�e��6v�tܩY$��t����h��J�Dʷ�E$MP��1Y����<��-A��Q����`}�ϙD�����Y�JJ�B����=a����>��{��J�����rAW�̸�K�h��eu�Y������_��ME�Kf-�yO�U�l���*I��j�|(W���DY@�ִ���A\���ЕO������#��=I��n{��(}�����iq-C�ʶ��gU�����Ww��R�I��NT�X	\˂��PH�<��R�$�ʓ35��bu�� \������*�P�-�hT��''��Dt���#�����YRB��@��t튑[����G�_.m�e�ve%�B�p8N�z���jswA�32ґ:�{��&����G���&OC���"��r�E$�D|H�;H����Yl�حCo}d6V��¢&�q�B3���ATy,��J����Rh��['�.@R[��Pz"�'"OS�w�4sy{��G'=�&�`���eYM_|c	����R,�&��2��ZA���AG4o�AG�S
�/�6��V�!��C' �G�=[G����w���}6���i�3���L
l�׹��4��wnd��*U(�CF@gT�:�ZO��5��%�C��[V5�1�!ˮC܌#���2L�7k�@�˚�>��~�\p&��n�j����\a��#�k(H�d�u�R�w�V�fK8�R��^RZهr4cn��`�K��8��fIh�*(��=��A$�	�F�jV#�G����(^�$��O�r}�?��g@�?c��{�E�P�қkt���ȱ9�p����id��������'̉�0�W��,�N7~+k��� ���kW�;HQKW�EGN0`�{��x)+䭝ԗZ�ը�G�|I����u�����`o~4���ڔˀ�]N���I%�.������Ao����]�mĶm�-��?'��g��OoW 6H��`���-vN���x<R�ɧgi�6̉���..��t�{�&�6�E�H.���-���m�� tV��h{�LQ_��㈰�}|G�-ur�ߕ���A�"D�^d.�c�}_ o����mJӸ:&���)�-.��ll�A�"Άā]#�Q�X��� �m���\��l��dm{'7�x>
�}��j�;����;�0I�)Z�͔$��i)a��^�{�R��[�&����^Q���ѽt;�l��Ѱ�틖jw�1�i�ah<A���T�:��Kۿ#�~�
׏dx�ow4��@��>.{�[e�]/GǓ��W�u��#G��>�k@;�s4>?%xQ���C�K*HP�K��Y�Ao�*�7�z�M�6p�j�X?t��d��gu���O�J�Ӌ-��{+�	
��o�޻�遾���,���J� �y�Z�E1�,aVNYc�����եi3��X�Q��ڹ�Yk���+���JAdy=��{ϸp{���=���z#�V�U;���5\A����z�S���uD�`����|E����R�����n��t�ֶu�����R]9��z�*\�#aD���{[�c|�LӐ"�m�z:t�L��S7�I�&�G��M![>{\�߷�$���3С��~}<�u�z�,�8��s�Ī�?@J�
Rs����,J(d��6f7b����1��3H�)�������qS���R۷�k�I��]!cd����O᝟��.UI/��iD�+��2V��ӝBy�5�F�=��T�f�kr�>5���{�
��ڈ�gc��b��C��>M��a�^��1n����#|���M;�fd̗�H�BV��٘���[@!9X�J��
����<xpά@Y���"3m#�����\&A
-�#�����2�R!��o�	ϙe3U;��0>�CF�:��+���o~��b���Zʇɬ(�1Ž2^>~T�!��aCz� ��L���GкQ�~Y��G��@!W�YC@�O:'����rlp"N1B���+O��͎�w��1h���L� �����\�����9�������,�w~u�j�%U�P'e1���W�&�;s���5��K����f�zh��k���}9�K������p�p��vV��l=���L��a���D%G�1Q����g+Gn��oyE���r3��u��ּۏ� ��$ע$љ�Yk�^�=Vڹ���C���Ug�O;��g�M�d�q�@BY���=������s�0)� ࢐"y�uSAQ\Al���������v;�@�qS@kZ{�s�2
�x�?i�|�s%�E�	��4j�Af��ɸ
���±)uO7v�+C������!�5������O��Hķ<�������
T쫽�����#"x/�a� �{e�'���Z��A��q�EN�[z�z��kJcM�<tzߋ�z��;˯-��y��t[I�s�Y�|��}Bx��ϣ�I���B�Y�*}�u$o�eF�W��[q�3mbG�k^���*�_.����sf9z�cf
\�r�ټߦ�J��پ��-�vߓ�t�A�o-��Q��)V34�ʙ۱RB��0x��,F��a�o��a�����J����#;�.��kZ(���-�j��ף�5b�ׇJ$�G�aW����3qo=�����ӴG�Ytna�=�^��S�ņ��m�Ā�}�xцj@��ӄ$��0�LO���;\�욀x�gi��)���Eq~��a���ϙ���}\��qsb7O�)6�p���3&�n� q<@��*����m�c����ʾ2g��P���.)�1�$t��M�,�Ytj�\���Z�a�	��wZ!"|�(~�qF`���eg�4{p]OK`춵!؎�0x�j́W�ʙ/�(Y���O�Ȍс��R��Y�M��iӀ�v�!S�	G�=S��,���� �H4���x��tK)"x9pW6x������3���,&N��up�1[ �r���K\��Y�ݢ���t*c�ڗ%�/����Tw��(�pm
W$�WiX�#�����/糮5J�$i����MM�/T��=7��ͨ��w��0c��G��ѹg��N&��c�f��&�=�+���c?R��)vY4H���SvO�C�[��d!\!��9��vZ�
��r��;�ߵ��ַ��F�k�`�<�_&j���XPį����;(鬴��� ��"7�B�DH�X��߂�܇�4b����#ޔH����ɒ�����<7����Й�wOt���l��$;�CZ��Ft�W���m�Y�BN�v�B8����:��s��k�o�c��;��;{����L\�(_)g�z�ϵV�hk�wRy~ ���W�(�������Y��yl�y9'F����r�D��E�"�X��Lѳ��f��)es
�	_��/�$B�5J�X3���"� Fe\.I���?c�,�2כţg���ݞu��-�ݺdy��Ϯ���������g�D���6-�N�����Vz/D�ʏzP����
���?4)NQ�`�I���u�*���ߥ�4]�mȩV�C핑o7��rIL�!���߀�g�j_Y	�J`a9�e�e�Y-�;�G����RsgU�F��ȳȑN5
~e��dg��]������
(���YG�,�9�X_�"�NA�CM�o��68� ����3o���a��6��Ev���8�9d���H<��?`��@�]���Z�Q����ׅ([4�w\�?R/�o, ���������5ytW�8\K�x_�*�σ:�\9�w������WY��̐₦ѣ4�F5,�����K���/ *B֋�c��q0v����f���twҺ���O)me����W���B::�q�P��d3W���Z���E^�$�|���qy�5�QW�GA�oT�}���*�����܉0�n��l��M.g�M�G����z�b�mPVSN�FO;M�oG0efbY�@�0yЮ��)�yg�c��g�czUZ*���>hlRj5�g��=�!����i���u���*?	�Q�bJ/S��( �E[����[+H�pW�Ђ��l�S�Q�����D���@��xS+K,����{exCŧ���ÙH;���+�\�[��upW��8��\IsGC܎�n�� ������23]u`����s�u���5����.է��^�9�*g��)�B���j�;�#<�KT�r۪nh�u`�'����,�<��x���|���T��#�B�ߢaY�\� _��ζt�z{���#ְ�rF�T������:I���Ax/��	w�Jkޡ�t�\mC<q�Ze���L��q���y0W!g�5��ѥk0b�?�>桶����l�cT6w�N%�PaWW:m"�oeb�}���Ub��|�`#]?�4�a��n�M�!=��˽\����� ��N��Ή���M��#Eɞ�Q-K�X���(A�a�gAk�,�=C�l�gG~�F�W�Kl���@�{_m��-�����]�V��E(�G�� |)5
!�%_�x΂���'���瘀���	 ΙC{\o���`t�����twx$��{��Am��*����,������{̵Ƀ}�v�ρ��h�)Ե��+�wd\�PLP=1a<	,� n����U�b��\;ĈrD�W��e'%�2�d���F��%�o� M!����_#�t=O�ǄIYFf¡�-���1k�g�aM�����]����l���I�k�Zh�E%�޹�1|8��3;C{t8���c^��9�H"E��D9鮢]��]���	��aTX2g�V�+5���s����1E��㎩���1�����.ׂ�� �nг��_�`��Wq�G�`�v��P�4{��l������\�V6��>?�4�Mnr���^����;X��>�6���C�m�u�C� ��6��£t�IQ�XJ�
S��ޮ�l�}�hS�H����nܠ�{Y��И��̌��Rh~��i�O�Wuh�4"��X mn��O]w��sjH����J��}�Z�<#�=�ȫ[��ݘ���;W=R�ǡ�F@g���
ҹ����>]��K����%0�	�d!R�'�n�\���ϫpj�L]߆ą���xB�6�G�uI�ႎv��F����#�pŷ�X���1�/u��_�}I!�\}+{I�V�x:�v��{8@��t`�"�@��i�����z@���ݿ����v���~%�م�U(�"�^K3�XJ��#+�	��qJ��^"^X�]���W���[�0��~�yD���n���ݜV��|�mT�U�MPL�wY.h��q>6�nO����1[�n�TmŵF0 ]�Sq����q�Q ì�*��eW�1$���,g�iAi��^_҃�#I[�v�m!��g`*D����=�d���jW"���܉��:ԋ�_�=�%����>F��g�����,����r�g�Z���ٳ�2�3n[
��ټV�gBo-��ﭕ�;����
ҙcB��hT4��eQr�$�Ћ��u�r�j���ͷ�ML� �?Av���ar�~o^-�3�`�V]ͦw3sS)�#�2�!�P�R��w��t����$mID=:&��6
�y���A%<�Je�!Òv>����'�Y�������M��֭!��n�|-4@Qo�HӭQ㍟:��r,�Y��i�	t�T��<��ި���h�=W5�z��W{x���Y;U�EnV�kɕ�:�u� Yp�y娟�+ʽ����������3������8@�ߊ�!.r�Q��o�|�|hG���7Z\Ҏ��?`�
��۲��O���ɠ���s��ƪY�kw����(���k5����׹��w����O[�n� M��fo��X[�=��<O�\���h�x�͟\j�[G�K?t���A�6[5�>pOl�S�F�mO������Ʋ��]G����I��{n��c�:�G�h|֨�]A���W�H���)�8�?w.wP���	�������Rx��F1T�qPܪY�l@�\\����x�ȏ��ʹm��`�'���X�[(HՏ�w��k8c�tԭ���=�R9�NQG����O���cL��2$�n�)�ֆ������,�CD�e��NXZ{Be����}�z�%��i<��@%���/{'�!� `�\���R{�$UĪ�/�����r^�%8z���y�:���Y�M�)����	R(�-t��4�=^<"G��&��	+r�.��R�e]�rF���{SYt�(��������k��&��J1��sow!����z5!ҷ�^C�|�հ���M6~�.@VL��E�̷X��s����f�qk��ΕX�T��㒾����q���ӇD0�R��x����������x92���~�o���"3��:����6�C��,���񷿳�9��]�]��}cm;-5lg��I�˳H��yw)Z��Y��.v�q��H��f��������� ���z8��S'+k���ׯ��D���7��W���)���e�V
R��%���K���p�^�4J�s^�`/p���^%
"Y]���)D�7�ȃ;�u�_�t���Z�E��I�����pSXA������?��l�e#@��D����x�#�\�P��w�G�1m��JK�[5��G�5��Bn�q�}�+8���Ű��2W�^��ص��)���>��]Wpdo� E8F4����z����xɿiwB�$�	��~a:$��� �ݖ��B��$bOJ~�B@�`�9lES6�o�x&�Jo�o�a�}D:Sz6��Y��A���2�H����,o� �[�Fb��\H�E���J `�;��h! <���7:ϭ�Vz�� 6��"~�$�v'x�=K9����|�e�Bt�9�mZp�l��!��N��w�:�|�=/��t/x+��*Fx@ړ�s �d�w!X9C��mf�X�����W��7�"�=���iȯ�q}��t�=YH����Z�ܭ����?�����������RR,��3���4z>��4���G�*�ց�w�-�[���;���1~���Ƕ׿�����8lqs��U��KX��WH��V�g�u���XtV�g��2b�7;<x�f��|i+��u;��j��D�9�ra�+��7�hLn\��_Yn�\>����j o#�� ���M�|��~{%�c��t�j�^>�Vr�ci݄�����J���nǿ��	�G���?c�.{@D�oKX2�G��꬙�d�Q�1��*g�M�6�A�Q{�� )b�0�H�Kz�w�k�J�TE���kI�Y��x�l �(GO���fb����,�j{X	���P�������χ�i�6��}g�½��)������^H��`yf}�z�g4w ��ZV���yeR�e�dߒ8]��S�u 
��*r�`��+���$>6�`�� �TQ��q�{4���pc>�&
R�|>J�S��(�`�}��<3�����6-=5��u#Y9�͈��;gS=��J��)r'�,� �8ە��(xhx��Ρ�դR�Mq�S�F��)t\�>��s�R�n�c�CA�M��E�Z��N��cP펄��C�^	�5�S��.Z��5`rl��+��[=�n��]m�`Il�����0�����t���7cI�T�9��J��Bt ��q"������=Mo�!�����փ�S�ӟ�e���QW4�>P���X��d�Ÿ��gT�F�[�S�L�`�Ϥq�Pzn�O�PzB[5�c4���f�p���� )���1n^�]����b�ܔ�_� � u	�
Y�i�1hpB���� G�c8/�Da�ԗ��9`������i�n��E�L��B������N�����[AbĽ4���~%�4<>6��dy��� KI��T`��utS(͒E�yh9���S��j���T����MY0|�̟H,Bq�Cyx>��H".�+o�pa��V�H[��"��"��ɁD ű���:�G���M�� }�Yx�
��"C���4~�7��e���/1�ĘE�E@�5G��#,a���Ŧ����d(� [�U������Ck���<[cڲlȾ^q���,
�F��@��6E܃�$:!v���+Zᗈ�8TG4�pY�%�2�0�;�Z���b��P@f�CA�7?�_?K��{��.֜��O�����n�=�����N�����k��]b���D8~-�3��VTw{��RA*������o��=��w p �?�^�1r�G:+5 Q	c֮��P�<�!!������o`��Ĝ�1��>;�>���� �?�ii���6��}�m?￦>�{��z�n� 5��O>nv��2��^�4����ƣ
��S�uA�oݯh,���{�{.�ZD��wa��֝�
�j
��_��2�,�>xւ<:j��)�kG��'vg�NA;��<��O�pq^��
3F�;"�+NZ����㬇�\�<*A������w��N(w�ϛ������p������	���xֳ�p�E% q��`��� /�^��7���v_����H�:�M\���n� YF54���t�ⷀ�3m"7C��"�`�j�&L�E�4t���N�F���yh�s��N��?q��Q����&$�V��3f��,Z˥�!�R�)��cZ�̕p��lA� s�!�]�C���4���r-����v����r���³���ȇ�U[O��+HD�g��#��E��&��������J��L��߆/GA�Qmd��	��Jm� �OCN�Ư[� ��� чY�aE��C�n��)$w�S�?3(��F��BU`Q���e�V�L�V��x*X���Ľ�R�^Aڑ~e˸
'��!������[��H���^)d�t�A6��Ĭ�>�������'ī)����l���Ӗ�a�YN,2р�j��d�p���𐻭��w��q׉D���)��_����k�1@�SPsH��aM1bFw���9c&��K��$����W`#hy�<�������Ͷn�|����h��Z[�9�l�Bh�n����������g�@�B	\er��W��|����u�jGt?���:�؅�N��-�۾0��]�Jih����]���)����'��RS*kI��L4�He��,"����Ш녤�'���n�r����
�.�	�S�� �rd>�T������v�J��I:6�?���CE�v��<$�j�<���
t�:V졹;Q`�EZ�T��0�yG���V��t��(K��6yB-��B�2� +1$8�O�_b�#m~0vx-�	`�GƇ�c4����e�p���"�n4e�V���R��gZ,?P2�͙sJ�@��%xg�F��ot�{gx0��B��B��-c� @�9~�Ţ�Vf���4]�)��L:��`�a�`�l(w
�1��W�����\O��wͺ��k��k������P�8�Kc�eA)I��f>tX���uٲ�vG|;�{=���=��Yo&�u �}v��Q���ڭN+O�e���ل!�� @���*�1�
9W�%�r��m����=G+�����u�K������q�)P�Z��{/!Ԝ�?�Ÿ�"T�ͅRr1�r�o��w��0?��E�s�ulr  �Ħ���}Y�����H���-$��,|wKI������?���ƭd�0˙`��P�N5Z�YZ�}�ȓ�@�!�s������H���P7l���J)��1�~=�Ũ~O�������6���9H8bu�@�ɦdeO�Z6$��]��v�<\�҂��HY��P�#�l7��Tv������� �L]�	���..�0���>�`�ٙ����[�*��E
2!R?8�`h��2TL��ݮN�~3�3OZ���}l^P�h/�_#� 3��m��nm��!�`oH�,xh�����T<а@Nݑ�
<+�^��z�cQG>p�)���Dqq��dt�"��-�_��`���]��n���,ǴMI�B�|-��A��
6մB�j;-W�B����Q�����L��T�R>��"%w� ��u�.x�����SX��Հ`Ҫ7|Zv��Z��
�_\����w�-w�>�%��<�����k����@�J�(sz��d]e$3�\���^HK��z"z��?��}�㱍�l�����E1�
E�8�RA���^m����	1��O���*L��i!E��'!���8-����-�w����Ϊ�Xr����#�/C��쨮�������l�� �jW3�2�;\���
�����+�~
R�Ybύ���}�$|�@2�5�bg�T_I�8��g��=	��c������AUjf⏘��-K���"����Sޓ��h�OH�;*!$xC䇝G+���+�?�X�W���^�[��U�G(�q?�3����>�.��)�%�cڮT�d�	g��9p?�cM(<����Y6�dI��9LoAz��VM��M�����,X:�[��P�|��W��9o)M�k���N>�dY-�&d��%����: �2ULߖ�?~0p ��m���~����j���!(�z���ZG���@�'����|'P��u:��]�/@�k�R��!ò�����zgi,|�|������ܟ�r��|��͈��$�����Bl�'/�V��&毼���q(9���0�D���5�nKx9�7���h����B�w�z��
Mn�����Ȕ�Ao�����\QVG0�
���K+W��v\4N�qo�OB�D���Fn��?�2��v�@����^���e�RIѼ�z`��0�b���S�W�O*�D?W����@����^_a���O���e��-�D����!R�ƮQ��!#�۬�ă���~�7OƷ����V@��2"���>�QijA����	�����<On}24l�SKp�΋�難��_ ��U^�ȣ]�W�w>� �4�hA|��f����l	���η{ �ؑK� �����\A�!����h��x.XW��_�M���r_i���
<2����> "��\~�U�1�[����P�����Y�b�?Gi����7*V`��~�a��"�Ve;��X��T���a��T(�d�	U�Po[}��g�k��QvU\�0���J�{J��g�`Xƈ� ͟͠�co/���*H-l�Hg���v�4ӳ�3�Yp�`,�ZvM��Y&n�FL��(�f��G$c��V]�1A����h3�~F-��	1��Ӯ�ӽ�%�z�|�iۙ��	�+]D����.0��xd�eYķq]�I���R�a�-�X8~ra��sծ��`�!|�$���[�~m��Z��������ݾ{)I-���BJ/�d6zP�@wX¾n����H �{ѮQ�QE��JV�x�h�	��q,�p�8k�l������m;�ϋnt���ݾ𱈪x��eB�g��,������9�}�v���;����a'E����4]��?1+G|w������O�����e���Kl�!GF���݀&�v�2
��q��T�7���K�{*H��E8ꕱu��?��vo��ߝ�[�U�e����=J���Hĉ<O���`�-�T)�v��i��~��I.�m��J2݈-��E��Ɣ���L"3����[��<��Jd�G�.���7��-�,r��f��E8�s��^��-�6~�:�1࿡o&6l͆"��j�S.od8m�1��.�Y��
-�<�j��v��4�)K�:�Ў)�b�ׂU����H5s=�X���ɹ�T2�TBFQ�8^��nB�~1x)S~���9�~5�SA*f����h�=�Ty������;����2��������* $�ǲ��,+O�ƛ�����4�-v|���Q
�K8�hYW(��?srZ;�N�fXI?�X�F"�q�o}�הl�Jw�HAL�)^��������k頥��4�nr;t��=���e�3�C�WbKZ�\�AI�Bx6�,a�LEJ�2�[�nk���n��	�!�W�6��,� hF/e��>t��Ꮂ��
:Dd��t�'\�r�{5����~r�A�ĪM���'��i�~������8ZC	{]}x+8w![�I\�;ͯ�4�2�����
�j:0aT`�h��uN+��*B-�;���J�.��SDAh���ը�B�L+4��� \E17��� خ����m`�-��oL����;ͳ�yo�OGW8�+��
�������gɞ	�T��?�'g��ڕrv�΄�9���},�x=?9����YwvAG?��g�c�k�7]q�P�44~j��)!}tm�F�� 3�r���{T�f��J����R��VDʛ��y:�Ĕ� ����\��ZI.��c�v0
aZ�j-�jr�_\�9�������y�D������ZnE���7�/BƳ��P>GwZ�g����{]�Gd<ɭ�N#�{�+�t�o� ��"�̾'$�*��*oԵ�@���8����s�@E�!�W���� �|�d�#(.n���
�����_���ayO�D\S<	�^m��k�<�Pр�^_F�\'g�9���i/����?�0}���4h�q����9B��4rR���$y����d�d��I�I��o���0�k��u)��
��9WAO0�;��8�i�1 ���oK*k�v��ff�52�4�,Yn@�%��P?
����x�t��v
�&~��X�~�[�{��R^�(��.�D,Z��ql�K/��W1��z�ҳE��	�o���6_�N�oY���;H��Q��~�7!n���Ǖ�<���{�����?Bú��/kbl�Feqe��ߢ�l�(c���9Zx
��-���}:��W&�ƴ�D_����}�ϭ�?�ǘ�����۟�a+�m���YiXޔ��Y�.�;��������i��m��m��H㱄/���e�ʡ���706==nf���:�yV~v��Ϻ/�!k69�r�������W�`2�Pce�4��Y���r<�hMQ��a�|�*G�D���?]�7Hk/e��Rh��\���w/�k3`!*�C\�+)61�F˶Ȝ{T�]i��LɸEt��8� pV��g�4��d�r7�;ݻ,�߄�{�P��$S$:�|��W<��s#����}�$�@k\xpC����#�W�f�����@sS��;�j�-/��)H�㳄����=��'��J+%����֔�y������H,4F�3��u5�q~T�}
$A_�xX~bu���Ԡp�BxO ��w8��]����|��WjPg����sa����AaZz��<z`X��Z�Q������1Hf�����&hhL�H/�8'�u��?�&�A���T-�xVO��	��ā�4�s(J�TX�09�"W�y�4�̟H1�۱ H�~">``��/HC~�U�r>�5�)�!��1y�bDpK�iM�����b/�"������D�C^+�K1������b�8�Yإ]�b��)�ӻ#�/���63
�Y 2����i�EZH�\��GX���-н0�r�Y	X���Ҋ�U~��������~����
*-�����ؗ���D%���T�Z��8\����k��,ݲw�883d ��­�\����K��af��)��?�y��,%T��%N����.��uU��qʮ|>Ȱa�
��E��m!����b�-el%���.Zwd>�U�H}�}C�����ְҹ�d���u��2�Z�?����]{��=x�Y���B�O�뤢?r�Q#ʋ���
R�6-!�KD�^b�s�;Z�%���M�_Ыx�n��;W�RD%
R�*��ڲ���+�I����ѧ���A��+�������&��`q=Qv���l���bm}B�t��@����A�Q�a��@�U����szn�������uB� *�:�rp+�"�M�uPxdDR�6�1������ͦ=����ot��z*�r�}���D%	����pF
����X����ݘ�����0�45Cv�{��sVmGF1(+S�W����7��ٳ���G���M��DV��%�oW���j��ҋY�=$6	�i�-ʒ��a�j�Ma�}�<Öu�ڊB��=s!D�c��S�\Ƹ�"�e[8��2(p"�kK���p?� ��_#�|QqO��:mC�	�"�D%i;G����z�Bg���n9-�x�J3�<�,��#�k�v�����,�}R�=&�ƕ�R�?dl`g��?q�(�'�k��"P*�"[���<�c��5`�u�q��O�ux]1�j�	!�p���=dI��������m��I��Wu �1l��F�3������7cūb�wa�2�t�5��������ݕ<	�%���<n��fV�;6�D��%�퀽�Ǐ��Ih���%��f|倾ׁ1�ݧ���ƠI���M.+��z�so��O�%�����W~#���G��=��50��e����_�,O�̤�rDs�&�15֢�~��6s�,U��@�����6	$�4��u�T*u�M�d���,5�k�%�3��w���)"G͢���, �g��r�`������1\�#xȕ���щP	b)o�
�� �Xo�hL�$J	��m�_h�I��&b��5���������S�(g��l!�a,� ��`1�d�N2{k�@k`
G2=�ZX�����X�G���Q$�ۼS�g,��qr(��\���?v���W�vJ�@��p�i�ŊbmŨFu0+egF_9�F�OZoܭW�8m�ή�3�&�/L�?E�1�)~�K�&���n�f���5�W{�_(�Y�&����]ѧBQ&u�g7���� e�Yu��=[�(���8FH�~�a�Y��%��fI��/^�9ӂa	��+�*�V(�JPQ��:b�Ĕ/]t�p��t@���5�9Ft�s ���ӖT*z�	2�T�*��C�P�ڭ�fä$����F�'
b�����������kr��5�`�(f6��`����A-쁑NL�;2�WX�/��+)?E���r���^�-�?��&��P��t�!�/.L�A=G[���l ��*a�[�gAԡ>Pe���Z�0����fڹE����'�8i[d�U��N3�qM��ָ��Y�����C�z�ĨX�m�����qL6��,�����ks_�\&UC;��|%�3�z��0���p�� .]�B�����;���|�д�W���{�F���6���u�.#��%�?�muoudDF*GY���XT^� �3z��X��e
Қ�7���!l;���39)2\�����s���Zf���G8��gqqt�D�9Obv��525������ǭK^?��^��5�W$�ew-�i�a�w��9�k��k�G��.��в��F������H�Af�� �����N����D�䐋!	�ug �9D�Dt��[�vТ��0��G�Pjcb��V�Lh��q�!3��� �_`
͍�|mF�u��-�p����Gxx�Gꬁ	���
A�����������`�pf7 z,,���Ϫ��t����VB\yWw���}��B-d�H#^r?66$\����m��R�S��c�k:�(1���T����]�~����W����.�n��?�����#+�T��	y��O��^�����s�E !�7���{���e/b��wV���d�#�Zp�R8@YQ<��N� �	֝�ű��ԝ/���楄r"d��o�PcR�j.i�sR���`<�y��Wr����q�k+�|��(�&�l��w�v�.K��I�3�U����2�/��%&Yo�������73�W:%��`!�l��w����\��A�R����#�!gB#4Ι�ݠj�w
�x���K�� ����S�v�Ms)6�׺V��i:iad��.؄BsBڡEpo7C�G'+*n���_� v�@w�%��(LR�v�5�:2z�!���!d�釕lB�f#ޱ���I[3#����+.���(�@���o�	1�����*9@���׾S�K4ly�w��*�w:��{18���V���I�嘍9r��,��Y�b��]C�?C���4!�ܗb�k���+�e ]0� o!���W�B�귇��Yra��̖�,�.$�U�-͑>}m�]"��no���v��+�>�Q$��b�*P�������o���Y��������� �3EH��������)�_?b��_IX���N�T4�B��x4T.j�f;Ir-UKACև�3Vѐ���������nt^�)����]�8�$׺,�2_���u.#��R�8ީR�a���@��r�<C�1��-ߛR�W��]��w1��[���e�mys�<[sܚ�
$fs��zhD#,��=�C9��s��+|o��#���Kg��nQ���Ȁ��GH#�i�ȗ}��N�'8('2�T>gT�_,��5�/�z*xU����`�G�clg)�g)Æ����&�&.��u�O�)�2|�KB`I��R
1�ǔ��Vx>fFax.*�ǋ�J�i�9�tk;�������e�:_��3���y��_�Hl�YG�-�!0A��5pz� @�Y ���mɲ��ba��e�#��@�k���*nc���_�&�M����1ɐ\W�҅�񲻿�h;�!�ш�0���SPΔ����tsd<�F�ߑ	�t���δY��+S6fS�����~�����ߏP�{��]ެ}��^�4Ğb��Z*}�XxZ�h]8��5�[z��ƿ�ٯ�����?����Z��M��� �̕)�YfE6�)/Yikn�ndM�����d�4�\2F�~`1�Qv&��n���7D�'��݌���!��_ѝi��T�70�85�\���H�N���&Tϝ�$=�
)�s�]zo�W�為<
)�������ϟ��������=�ܬ�	��K��"�2�<:��Q9y�r2Nj�ĝ�/����/�ݜ�/�m@�ya�\���}���7}��_?���}�b
Z�D��ej���R�`�c6�L[��Y��o�>:4�*��D]F1��]����f�͂��+��_���&/.��|R��i���yTEX X�0P3�\�{7�rA'"�-뫭�h�ߨ�Y�uC�۩����g$|N��H9������$ج������������\y�� ~1�<�Z��D��9K�y��Z��x���@�ʹ���4��)й���p�L�_\gat�B�n�?����__{J\0�ŝ�dqS�2�
=	r3q.i��M��+Y�����0į������-	'7A��J��eg��:&8�>�9@�.�������J��2/�ٟ$���P��"�m��Tً��~����û\1�zr�ʮ��1�K��!�5�D3&��^/\nۇ��|�|��������?��?�c�y\�,G�Ҿ�ϻr6�ͥ@�}��f�R�@{�5s��E֌d*�Q��m�S%�5
��������!���g!��i�F5�93;P,��h����J�w����G�3��!Hۙ"�������
�?���	�-�s`��n��ٛE���Ab.� R��U^����ҡp�#�K�4��}�g������m���3��HT�X[��=� ?��De� ��H�!{��ؾD��|;���������Yw��iw�kH�Kt
�:\��HC�+H^T���aiY;�����`,�.\Ϫ���>�-����L�R̶�A�èEҏ��'�
n� m����������I�9<2eg1rr44Z�"A+�I$��@���'��I~�`�JVE�Tg��\�3���Z���1kq~��?�o�<9c!W���Ve���(��_��'UYA��}�7�B�W�R��y���Ͽw6l�u������1sJ�A��+{�"Tf��+�Ԃr^ԋ���|������\Z��&!~��~����|��:�h<f�C`�*��8���qbT�寿�_?��W���KD��Vq�^ˠ��v�Ҹ��Wa%���3�E��:�v����f��l�$���w�4�l�����uDM`Yx�녞B��)�˿7��������-y)'�C��GS���͉/v,L�R���dZ�ϝuT6*^����Y���\�K�ZC��@�=��{?��k��w�h<�a*��"��0��_�a'/V�뛜�?���_��H}���.'�Z�\*B�62�QW���=����\0�"�}<%˜E�<r����0SB���o0�7�|>��/�:����������3p?i;��o���K�-���5�ܪ��F��j�'���xr����eWj���φkI^	l�r����Tx�^$Q��V4�ҿ��$bm=@���]�"���6@�YӢjCnF�J'v�RD7S��d��/l��хʉ=?;���3����F��{����СDc�1ځ�G�������.v�2�����b%���idK_q��=[�$cbh�K���\�s�L�?y$��DXG1������y�4Μ���sG�B�@��H�n��_{������V��
���1���1����x�V��b'$Xl���LarI(݌<ٚGJ�(��4��+�1OZi��
l�;}����B>Q��1u�P�OS���S
	[1�Q@i�Rh�����{
�aa�����o��Z�X�~�ە�zE{�5ݱ�GQ������g�y/"��ݗl����Sh9b̷ю�Ӛ\��fl0�qUb�n�z7+��#��A;ү�cb[�K
ڳ	��E��r�W�ɝ��h��3Z�,��L/e�r��]�����?V�Ef3��d�~��L�^B\'�*�9g!�I雯�2����	����A��oeIYm �}O ېx-�e^�Z}`�&�^��-�Vay��2HgF^8���o"1��b۰�I�O�h�%�����n���@��*���g�,r�-��J�p0�S�.kq�ךW�1ܻ���g֭�L���m�Q�H���{&����w�X�D+��]b��h�VV�3�Z��Y.�l����<^>�{G��w�Zt{��������i�	��v�������>N��6��� =��~p�����q��|�5�8�n�e�Wh6��^ֳE����:�����p�H`����n	9ȍ2!P�JJ�¦&������E��Y��*�@��X����B��4�C� /ӑn� ��x�����4C�FeEy	�Ć�u=��Nߓ57B ��r��A^��:Z���I�X�&"�m�����������V��RP��Ufb�'�#b�0d�[ͅ��z��u�cN��� h�j�}>��Ԥ�0�tےXv��ʐ�]�~�b���{��ne���y�d�����a�R`w ��R�2`)�.�gmA��߾�ܬ:8ك,/�Z�[SZ1�&��9}�<��[��?|��*�Hn�)�c�q���r��ъ	y�r�!�'ڗ�`r�<����+j`�H�x��m�4���;p?���Y��AbM͈���&%�K�Sʠ�JrJ�xZ(:�x��,���!�w��g�p���a+�n^�
)��Z	D���Kg�·�d�se��bd̃Vv@S�u��vm/��̡����5��I�����t��T+4s������rw �zeM� Sql��W|$[h˨�D&�_�򐐥�ZjM�!q�@��+
]�C'��|�]��ago<^��C�Jg}b�Gg-�31���NO~�/����Go2�W��� �v<�2��6s��,x���[�}�9A���U�/���,h���:����ȱ�>�;�j�DN����]Um=[�	�$x ��5���P�H��YW>�lR����q%A���5�X��a�����u]B�9zZ��ʰ_Թ��)b��!���t%�B��!M-�ּ:@M}P�Λ�&��,W����p�R7���i{��Vj�m��'���P�i[�~PZ�pe����C�΅ʌ?I�Hc��tGP�b)����n�-+�Ţ\�"��]9hR�� M�d��t�鏴�~��H��'�u�-��ë�W��G&�'�Ѳ���)��$,�@�g�VJ,��^"h���3�GP��(�>"iS{
<x��3&@!
��U>��rr$OBP��%����B���sID��Z�[e<�|3ȶk՘:��X��ڍ	I8�4�|�Y�;C��_P聴��[ �����f{�'�1e	��^��0��5��^�M������ ��"3_W��	٨�{v.�\>�gꆍIcc)l�]����k��/e�҃3���d�i6-�5�)%����X0�2Ϻ���hebT\���I`�(�ή����R�T����l=����|
��ݞu-F2����c^��ʉ�4��n�/g.���Vn� E�+Or�q�������@�Z� qVV�m���N5��������e��)R��.����pe��
�L�\Uª� +NLc�㉫��)הN�v-��Q��ǀC�ӆqY��;�� ��JCQ�l+�t��Q'A�⑃� h����v�`�9�Y|�4cp��Z��1�^���+��N8� ��Ra�I8��p�+��F`n[��f�܆���38�l���}�n:�Xm��v	�d��""Ж�;���4�Yi-�=Ŧ7�T�܍�~�w�j�;3cSs�2m���wN�A���JQ}Np2>�!Q����ց��ί�&-K�m�_�bzQ�s��NTzJ�e,���!S�O.?c+3xp��L�B	�M�UW��NA"A,����@��JFfGYC����M��"J��'>Y����ɄE�^}�Z��B!pܒi�~4��@#���^L�]k���J�\���ԏ��9�2���u~6�F�(��c�1n�2Zp���T�myC����~C�d7@:T�~��!٬�i�k)f^�z	��*�ҽ�]8�5`1�T���ئ� ^�������`bZ8Y�9I��pM�	��nKtϐ�r�IO��k%Nh>�����.����c�1�`pwi̪/v.��D�2)D�p��c�<��٣xBK&�����o��v���\ϱVy��VF�$��9��@�Ĳ<���t��~��k}�#��W¿W�\_��o��>	����s�G�C��ܯTcZ�Җ�!��A9���ma8�(Y˗zo�,b�G���XNۭ�J�[M�-r��X~M�8�;�)8���7�'4J!�l��M&��Ӽ5F�]c�U�����n� I E��*�5z��DS�UY��"���LX�u�T\{� kp~��8�=| v�f|�,lu����k)^Ē��s ��,S��^��[���CD�S|Vl%�,E����	�$����,p!_�]T��زrx�a�Ā#�3�J�рm��#X0��P�����iA�����59�<ES�Z<�$M1eD��P�|OF
&�^�m�ÃB��4�;����I(��8�t�^,�J��_��d=yV�HSQ�G �N���:C82<<�p5c�V9D�J���Ɩ4�\0�um�)k��$1w!A�!�/���5m�j�+�C����g����ɐ�
`�E��>g�sb����1o>��J�k���/lY�DPc]��uj�E�#�4���T�#h�ͨ����!��\����T,0�WM�0l��������->X��w,�Q-\�F)�2������T;����&��3R_!���>�o��I��)rUOAh�A�&s3�c�M_S��Z��85r'�[8t�ZXkf������T6¿���_E�����Nb�$��q���PC��k�AY�U���o��aG{�F�֒/�2�ۤ����y��^�>���/����d24�}l�qč���M���>~��v�@o��P�g�ŝ����
O�w���(�+�8��i�4�a`ef-�o�=��[��F�:���D��f�X����3Eb��]�^3��L�"׮k4��a���k�Ȳ���لJ��Y���� G�"kS�����-`����V�	�Y8�'f�����GS�X5�Y@��ޱ��\W��mȋ`�?��TYN�õ2�:��P�!�Y�Y0���t1bs!�ڱ�mΙ7e��L�Q�\�B!��I�I�-!� ж��?��3��Y<c?��M1�幹���/C��A'�[Y�1�yh�c>
���Dm@�/���5���M Vo�X�ݻf�+�ۖLBh��WK�O�3;�V���v
��*�m%������---�K�ؽm����]��鷵�A����qve��+�)|T��b���74��\�5��ʑ*3�5qB�߳���Q\�ra�;zd����A�wa�2S0��	y�r�#�7N�a_�w�6]Zo�	�zi~\��Eijd��pM�et]@'	ϷZ~���|��:ˉ�I)M�[Z��M���f�+|�)96�+E���6�Љ�iۄa�*C#�v��K����X��}ֹ�V-�}�7�ؐ]B\ ��2��Ha��*�UC<��65�hQ��.d�����ժ���5��@��c<�d5����[*H��f�#cK��s�,(So1TK0$zX����j��`���_[ػ-q ��K���s�6s5��@��?�N�f���Va�-��k*�Bh
+U����?�ĩ"��z���ZߞH��5V$V��t�ÅHp�9��Z��m[��-�ٟ2��D�
(���(h�UY�s���H����&_}�P:&�RݲZ��|V7��#f�c��f}���e2T}�Hp:ȍ��P�	�y�Jg�a�i;	���.#;u�X�6��i����)k�k�{o8����=$�hɢ`���|w���veI��H#	�Z����,����<Df�s����S����,?	m����g_sϖ"��|�e����>���ۛ� G�ˇjSɲ
Lo4hT�n=��+1òج�I��-�0-��G��c�(a��h��ںv�#B1�|�s2\L�ޅ�����v�ܒ1f{�Cg9��P��3ݨs�)������ǃGz��8�iݤn��^8�H�`\�9C��  R�ҩZػ�r:�j��P]��I�_��F���q�]`�;�u-ް��Ь�=`�Y^��˸)v�곶Q��[X�꛹V�o��3�����s��l�D��Ǖ��H����0sza��=Cy�R{�P��z�ʅ��=Ç]B�x��h���G��A.��mz�@��eģ�������]"�ū��'&M�sF���W���5��G�N��+�
�&ΨF-���1��z��x.�
����c��J<+2���weѹtZDy*���Z�E5�����K�Wj8��=0�Ǧ"	�+5�zE(>]�-	�x�q��ƣ�|���Q
-_��W2i^�8Ny-�_N|�}=�e��yנ���l?��?�C�o)�?�37�|n�;�g"b��� `T^��}k��T��J�w�
q:�����i��6�p�����$)�yH��/����Qӫf��b��9����wb,�٩�b#�e%*@/0�4��ʽ��_��e��,�8p�����J7�ʇ�B��P�mN�|���ġ�P�C��Ԗx��E~ �ɚ��X�o��T�Oz�rLC�?�ƙz�?�mi����J֘�����w�]�W��í V(H�S���w��t`�[w�a<�����d�nyρq�k�� �J})�,�.���p[SJ�B�/�JPE��uԏ�g)|��U�!�9 C�{��<��M�B�������a1��n�M4�۸P�BI�AH4�������0��Q�A��i0s�S���]��-�<���`/l�Ba��D�������ZRr���S��{�8n��B��Dp�bn9 ��N?���Jy�\�=�=��+��"x��
:�lt��*<0�̠�\��@fI���Ϻ���M��m��d�,
�i��I�����Q�% 3`��}��1?<
.���6����|F���#gLᵌ�
�Rf��=)����KZ13���Z�1bT;��W��ּ
�Pނn�?��]����%V!�#�$��� ��FK�� ��T�j�o�n,c�ի�p�8���n�:�����/�"�M�t�;�,��j���$�0Y�N�q�{wl �8�Q�|
z�%ѹ�t��ʛƗGe���]�*�k>��$|�,��"��U�s�`�� �ƀ�����?&�/ҝNA ��X�.��Ck��e�������6�d?����
�8!5Od�F�9nl}ڐv*�7pQ�&k�jOq��_d_���r;�~ǺSצ9��֜�qI��\���es�a�lM��\��K����͓Ç�.Y:��]Be�i��8�VA�[R�__Q*�)�(��^i9m�)�Dph]��Ԋ���,bnPcz�Nj)��ŪP<o�캮����9��_/Ө�%�\p���R�����,���Hcd�Z�1M�����w��4NJS��I+g��"���Б�ՆO�޽���(�>��$(�5�(#�m�]��Y.�P�\��v���5��E��|��xU��o	���������;����i�|G�Ƶ�����������Q��O��u.�4
Kx�o�S̿u�K���*Z%ѓa��B�wp@.�2Ɗ�V������\N(���z�����y4~-`ckS{�RA�B����w;,����/�x����-��b��/FZ����N��,e�ǨE[4�o��!E�n7������Tv��ʰꝃԝ��=2����&7+�p�����DDta¦:9�'┨���ۼտ0No�������/v��B�'�g%�n�m��k@�҉��Y��5ź��'���_�Թ���웝	��@|�(��[�� s8ڞg�-�x;#�tx7/��4/ג��ƅ�Ɵ<�ǃ�1z��T��>f���G��6d����rt��6X���@H`)3��'*�j�B�A'��n� �{�����A4N+�j`<]vc��6Y�M6�m^�8$�m��%@�+�	�05�H<�j�Sy�0����ѹ88�L�ߟPߨR7&���Ya0ٳt�:R.p�Zp�e�Qx:.��iѯ���qh��r
��gҌ+�_y�3?��4�>_ˣς[+HY�|�p	��gN���}�0����*ȮO�=s����x������2^�Ɉ�}E�s�i�����vf��3VK�k�ӫ�ׁ"�[^�<���=qT!qݲ9�IN*�&�u�m���e�y:�p�����j�a�b�	d
�|�/0�	N ��X����;�e=��P���y&��J��l]aѯ�E��Ĭ6.��b�"��^K{�v����y��$���w���
��v�����q$$����	F�{�=�}�{�  �E�le� �ߏ��+�) r��?W@M.ז{KR���Q��d]�7�Ұ�?��k���{�n�~ǝo=ܯ��DoM� ��"+$�,_��y��Fg���<5���R�,�)��*��B�쀓�{�lٸy��ےxJ�&{g��jh�w^��-��T�n�8��w(��S��W��r}9����hh�08s;H�C���N���
��4��,�"5���u�(.�-q�e�~˂= G�-�y��P|��co��a)*����8�g��g�ir�H𧠟�k2�����f�ϟLg�MgT�Ɨ7��-��w���
ꯡ�[7��\9F������h����&h��#���P��c�P�87U�p�F;�fw�4�GW�q���J��[ &G�L����ͨ��ʩL���!��wa� �>-��I���~�b�y#�� �߿pg���=Vv`�e�Y4=X�;�IK4�^�0�T��b��aw�?+#��qD��|Q-��m}��jW\*جk�������"��}Gܕ�|��4�+��i/%Գy�AnmT$���>SѦ5�#o4��A	h���@��L�w����'/�l���p�#�vKa��G�;�����g�Ⱦ���)���M;K���e@����o�Y.���)x�q6�L�Y�y�<��8��X�A|д��N�[*H�������-��L�b(�*;b�1�%m헊ޟ=}���b8��O���[)�
��v=<h6�rg��!
�RQ��}�r�߁S�G����^A�ƴ��4�}_u����QQl"�1$4T�Q��]{��)ǋ ���4vy�ߏ+Uh�wo��WX�h9����7� ���#�}�j�e�˭]�{���&SD5����w^�|�E��8?|��*x���ν�\����od�ԃ��9
L�{�(3�6<8�,�go� e�6MUNׄ����Z�[`
}]�q{�I��[��Y��d�_F.�R�H{��=�����à%����y2��S�}+���7O�A//��MH��;*�j�:�����1��֙˗��&յl��|��s�9[P/�+���Ľ�J���WhyT����#-��M���W�60������o�2d� ���O��ai qb"m�-Bh�i�FAOU=I���#�>l�8�n�Q:Ey~=~q�����Hhƕ�;My��E�jPr	�n��@[��G�!��	�È�� �Tk/� .Y�z (Y��׿�;�C���=��
��_�� ԗ�=
�Т����O��J�ƫ�˗����7˱��YB>���д�=bTحʟ:��K���I�=Z�@���!7ctJ,��]����}�zd�s�[�+(��_�Y�l��r�&.�U���j� ��<���t�ؽ&dSNۑ?iK�֗�.[� ~p�?�y�2�L2��݈�����a�z;iWod	��@�hW!2�PTL͸�܃�nO�BncqVm���_������`��<�]�^A���W��.B��e�Ѵ��ӿ���:��!zA`����KG�e� �H��mծgɀa��t�~N|#��d���6�̊a���H���������%��/^O�U�Z@���,hk����J�)	�Lǭ�������҄��M�r�������C#��6��&4o���A$^�݇Ja����b�Mʤ���F�ZK�����|Γ��W���y4���;H��n����F�H���h�7�����L;%����o��a���(��%�]��n��Cvo���&w�|�U)F�t.?H��xAY�P��:xC�4ʂ�������#�d}�}�qC)[gLhH��~�l��Sy�#mѿ� D����7n����0��x���V3B��n)�
�ZT�Wut�#�Ln������!�:D����2b$z���̝"�����(h-���e��C$dʋ�m��%��)��*A~_�a�=����,ů�BAB6C���C���Ar����Ms�g��j9Sf��Co@��ߠ�~�bФ�31'2e{�	�5]D�o��:�XS�Gd.�%l
n���b�/�(�)�p~������o2���w\v���d��z �BAj�f�X!$(T;L�$PiZW�!���}��X�����j������ �(㋷[=
�e�����?x�{A�굥�t ��v�?=*O�Kwԛ�Q���O����G/f�;۷_J�tX��}pEe[����.+�
R�+k��K#�"��Ů��f��Ǡ���lb�2"s�1�>����J����o�^-כ�
�� ��C#i@�-+�|y��j�0���a9T��oo;���k�&Ísy�������x�π�[����E�ub��X��ߑ��Ĺ����X�STկ�AZxi�R�%���N�/�A���[��6t�>��E{O����m����J}��?���*:H�\(*�$5q���) ��-
:xC��n�'��Q�C�X�^�3�1��F=��y/�0�ߕF��㐅+H� ʺ���7�4֜j�.��\U����DռY�t�G]� oDX�g|���RA�092bG'����|�C�)�t��ݮG��)����X>p	\?�5�[�>p-�KC��?"�`��]��?,��S�u�Ȏ^S2~g�J.Lbi-Y����.מ�h��?�6&L)M�"~	3�
ņ�G�(��Ɋ�V�gK��� ��n�W��b�!o��0��ٺx���G��[T~'�0���b�x��9�����rA°T�W��>�~ShX�=��`���.�-x���1�{�Iց�c���N R�e�k~
tw��@���֓VTF�	^�=��ʾ�5H� ��+@[��7~�ܙOe�p��k�o�J��;�����l�]�	���&��h9��)f�|>o'iƫ���k�v_�m�hF��u@*� ����92�My��M�54�	rd�;�X�j�7Y�=��[+Hڽ���b�[0Bh ���4�̽�:��':�F��H��(t�\z��N����c)�
���7���\�(�K���%��m\1ۛv2�����0$����pX
��o;I��²���S&�/�Z-��Ui�
����o��{C�˕�N�ޙ�Yu��׳�
�� �hǓ;Dp�z�P�N���J�1�ϫb{����F��a��-��#T��`���v&�xL�"*�r&��M� �����3aX6q��׈���]D�w�r$���A�������D���Y1����9��w�(�JƂr֡q��R��(g��KѬ��qQ8�3�P���k(c�D(��ǝ=�p<-:̲���<�n� a�^��a�*]Tk�Q�E��y�� p��fZt�U��0}�J����	z#��Xz*�jm� wC��� �īQm���X���D�1���j�g�p�� SV.���ڄ�\��]�7�r0�������@���nk�n���NA�0���F�4	'�+n	c�H�i�l���玾e�E+���:<�������s�����a�G�@u���UB��kl��H}���s��#��,_����ȑC��}��zT�hHہ)�����<R��3��W���5tZ�`%��:���d�BZ��?�B�s�ܹ��AxC���#(\	�;�oii��e�r_��!��� ��7GF&�}F�Ѯ��CX�FJ�{[0\��Ȅ�=v/�s��/ ��p�)�#H;�]��ޤ��wΣkH@��v[�txI�-�H�����v�ܾ����i˖g�r⏗�&��t������n<���Oy�����R&�4[�vL���bXg�-��M��ӧ�7���sp��e�O�s�������˦c
����z�<�����KnX���3��e�B�m˺��k�M�X=�;T�]��`�_��T�\����u�#௤V��6�N������|�U̧S�_'�����-�vdN��02���AcGY[+3��6�Gt�/��6�UtЪ��ͫG��p�������>��!�X��Jx�tr�F

���ￋ�"�@�rvy�߱�h��k*���0����ڙqw�T��$��x��TCI2>�2�!���#�
RL��ty��by�I�z��d�@}�&�|1s��~h���9�I;P�U�m_1�є[C��d�T�U��A�1<'v;�1��GX��pPՕ��qT2:%�|��c��&h��::�k3��ww��V���_��<~c�.�G�SKW�TP����p��89HP�tc�9�:����ok���C��5��,p��#�
2}1�wT�|��x�n�P��y6�b;���g8��m�J�NA�7���^"6�
ѧƛs����@�$�b���BT���=���}����T�G��i��ʏ�`M�ˀ|0�1_\�s�a�Ls�{ V7����BR懚qKH�_��o30���:VS.��9��b�%n1֭�� �x�(��4r�-��9W���S���ڢ
A�g5��o��NA��y��Ѓ����*���M8fA�y��<v4�����`�z�b�w���<2�sA��`Y����0�342?$�gI]U�7ffO��X�����+��48��/�bp��C��3`d܍)��p9�VDH��rߐ}��^Sn��q�@�;j��^)I)/�]�{و�������L��iϣ����@�=�L�{���)H�d�T���-W��������T,!1�D2���(��u�o��cs{���!˗d���e��V����l����M.e��-e)��,��5جK�l�2㣝�$�e����r*\�s��)��m�M奄g�+�#o�P�w4%�(�p�w6��t���`���0��k:�^��O�:���!K�~ɝ�
��U��e)y�sM�n2)K ��R�ʧ?���Wv�r��wI���n�l�����;fg�*N�&�dSb�~)�9�}.��x�����{ц˝P�o�S�v_D��с��O��sq�xbr�[�]�iV�ɻ�� @��D�(�c`�T�*_�ǩq4�����占��g��T�n��A�Ԕ�G�d��O�,���1�0���Pl}�2��R7r<�)c�YX��$��#��W�sV���:��i��@56����A��z�'�b� b}Hk}[�י��=�˨�r�+w|i�[�]�=�'t���65Ux��ŉܚ�Ҽr'ں?�PT]��8=����<i�G|�������(��=/�}�r�I����w�t�b�8=�*�P*jWg����TW�m-s�W�Ao���z$c�ЋT>[�Mb���-j&�8OwF�p
M�q�/�A�r�˲i�y9e��w����i9�$<��M����#��dPZ�R�%��a.����	��_G�7^;��*VIsE ��d�Wh��ަT����}4dP���GZ�����4��9-i/�M�������qA1���'�.�a��^+o���'�Y|��5�a;?�O�}�`���.>���w�>�Y���542���J߶��$n�	ٲ�����ٝ/�[����yT��^��.?��]���j��ϗ�G7��n���z��lXt4.y�B���q�;�};ͅ,$���"!!!�ȡ���Ȟt�AT��g��"���;3d�|W�������@{[�����p8��aW�b�,QG��G�/!r�@�$U�/O��(�,g>��g�a���k"��+ �Sab`�X%�Rc�>��s�����,4$lf��S�*�߿?��p��� �Y�6��*F�#��!m�8�"Nڪ�w�S#m�d�I[�r�LBN�gȀ��h4u{�U��{��y<�����eB{��iF7�5Qg�ZE>G�r�~
��k�y`��fyBr�q'�,�mٯ?������3}��M|�:۰E���"(=?$�4�=3�HPV0��������HuЅs��Z�߾�D��H����LO|pK�����)k�Z5t��$�*z����Cf���M�R!E��b�=e%���B�v�d�ko%/cXtI���$��`��hq�����w{��Q��Z|z��U���͏�p�Fb?6:��$�}�v�ݕs)仃˴�{H|*nU{ښ���;y�Z� M��N�u�Gt���������א�݈��.|.K2
�� å�JCy6��l%��l�e��uԿtV�Om��c�y�ߚ��G������^Y���HY���p���r���72/����s#6�p?�`p�����-`����b
�R�vG@g���3�[���l���jq�7O3r��P>������#.P���,\�T��u��g���������t�>�go�'�>W�r���Gv,>W����`�5����[��+�;��-��h�0���������/B�o������D�&=P���t#(Q�K�Z��.��hco������_ڹh��'���V��&��ĉ�X{	��[5��$1���Pp̭Y��m��6?��Q���C���ټ�O ����7�&JD*o�$י{����y�Q��t_i ����SӁ+�Iy���f��V�����j牷�N��Y�X�S4���-�{b������E	��I����-�Bs�pe�����Ox6oK��'G�a64��p3��ehf<y��!hވ�;cf��쏚0�M-���p�O%���J�bĨ������.{ �L�F�2��2���J�/#d����ǖ�ԁ�~�>�!"15r�%���l����Y���jio`�lu�[F߄|�}8	���V���7��-41m�ބ`�E�|��%������d[�'���u�0%i�Z�qv��[��!R�l�ļyn4�(-a�\};ܚP��$�V����P���	�V�9��xY���
kj���Aj}�$����(�h�TcP�l��`���{A��~_�Piخ�1�x���0���5\r�j��	��P)�#����w�\s�B7Gw0�3|y��-߫h�Rp����G�9�"�ց�Q�9��^i	(�2�>�Bk���k�K�T�V���8+�nQ��Y�;$�3z�n�E�w����v�Z�'	1�k�K&��%Ary�+F̠���adV{��_`?�&Q�?g��L5|��ҍ�2�Z�Ƈq�ԊUj��
������:D������L�!��{�v��UVl\���&׊�o��#YF����*3_��w�X�v�c��|"5����+����s*���t6�^��7�����5=�#Y]����	�j�n2�eQ��O�����DO[�ֿ�t�_ U$�﫨�lF����0\�/��$��Z-�{d�+��tJ~��r�o��c���b��uGg� 3� 
�6�Ad�+��0�+���S�0�߃���4{�����q�a8�A�m��/�D��ӷ�T%�	<��O��sf|/�{*H��K��[���[���M02^]C�+�<���q�^�)Da�s`�%q�z�7�
��N�fG�t�`HL����Q o�`���C;�Wz֐1%;��ε�쩂�7���S���h2F���+��%K��z���*~Z�i��R�s�L���#HBlU���j����2 ��И�� �Ta���I���]|:�?���s���+���Z{&�5u��yC#�� A�u�p)�ii2�-��&
{ƌ��ş�Z>@�J�4��[�vs�ć��@y y��������K4wU��->C� ��O	z����bޠ~GI�1�kN��S���\�����Q��5f_����2��ꮬ<�&�rq�Q��|\�|6�㍓銎-ti/,�����w�j�?S��q-�]��<�D��j�v�	�cl�%��WG���"��z�5�����O�Az �L�y@�.���dYG��V�̞F�G�8����W���y������^dZ�=��t�F�w*h\���k*��u��ݠK���g�a?���8�y���Ss��8��rͦ3�J�yMV�����-�4�B�ڦ�'�|4�b�e����m�NA�+����@Y�v����i�g�Vʝ��P+�E�]U���Wéuq"v
�Z�cg�F?��TM�-;\ը��-�l�#Y�l�?���S�&R�
���ӿ��;0���p(%;|y>���Q\���I��6޵(EȲ�(R�N��r��d��JM�6�l��cJi�!hkJ�-|�1�PJ��<b��e�����p�����}%
oƩ]	Yۆ�RqϳcJ��Ɂ=p��F<t��t?�Z>�V�}_�F��}J|�n� ʙK�8*J���y�o�t����;0P�sp���lGG�<���B�@��l�՟�2gr{�Aͷ�0p�)��G��zY�c�
O�+����'0�a��X�m ؿ�`	�E�M�y�s��apHs�c�*&��]S��')Z�@������!��0.�	���ٝ�=��u,Ͳ�����oZ{3�P(�~����T}��m�,b�VxDa�ʇ�_?%�x9 �̴"o'�J�룵�[+SQ�{H�$�������D:|���<�!�C�Цu{��Y$g]�ux'g���c4�(ݐ�M,�y�+������
��h �0��+)��弚�U�����$t��G���aJ`�<,����>���'�e?�rp��"�΃��yQ���x�ܐ���)�Lݣ��kU��\�c�r�?��.w���4�\�:��p���@�P�8�9f(D8��[M��q7��yt�.����{M��Z�=��p�8\%��D��vN�ߐ�o�T�.��)Hy�NZ�ia�$�o͂6�L7���)�=�35����fDx��0��-���w��@����Y����?�޴`���GZ7�zL���7��3p�Hcj�Ӥ��r�rg�� ���� yhꞰs���D��<G~��[J�`%�>n�:E��ѾB���ɟ�y�x�(�*Y�tf#7[1���ע;YZM���4Y�AMe ��D�����2�7j����H����Y�y5:Z����}6:��s4��-m�ؙf(��z-;�輋b��H[q �Ƞ�|Й��~
Rƿ8b�����+�O�[d
Z�e�מ���
��a��E:#0�o������˦`���`�����!L/��J(FyH��� d 'z�~��l�9b_T������P�2��
�`8Mjo�m."]�5�|�LP���U��E��	X������h���:�c�%k��Z�X}��xV����M��i\��
G.sO�Y9����z���l	�s�.�.���;��5@gyi,�2��;Z������7��gy,x;�%~�4��1����/+�y�0��ZQr�߲�D�#�&�c��yؔsG�)����tQ���gM����N�a{��-�M���m|����l�%Jd¹�(d85"O�ﭝ�Y�-�qRi8o昼��4َ�Ⱦ���3�~
�`��n�W�q,i۟��T��GV�5o��Y�U��g�Ͷ%�u1B��գ�����5?�k��ꪛ�C$1��PDh��8'wH��Dچӕ��|��o��K����=�z�W��C�J�:~�TsZx6^����?F����k������;|	��=
?+�h|�s��Y�Ӄ���C߹�vtL}�=y@?
��@��]��gW��]o���s�)�^m���o�B4:}o9Ϸ'����{ʉ��+�y"Tt�:��)(de�~yU�D�vͯJ�y
�L>����<��d�AU��sh�0���[\��#�E4A��s���� %Y�+�ҊN4�3/K!.X$yBj�l� ?t��̷�l�ڌ����6e4�#Hv�
�S�Vb~,����E2l�j�֨<)���k}p{ˌ��+z<ےb��Q�ه˛J��{ʋ�=�!3I�Ѣ��=�<��Wpm+��p�~�_yQ�ٱ'�/�W�y:'c�nj1�n7+nH�3�v�l����}OI}�s�7?��i3C�jr����St�)7�J܂�ɭO�@�W`�cw�����V(zq>)k;�m�dq�ݩ��6f�qw��N����T�x�p�,?������#H
��S�a?��:¥�Y*r�-Wd1��nW�X ǝ�r<J�����6�����ZK�sr�p<�W�Qܹ�ul��fC�MKz�AA����[�X�τ�����a��}��ן�zW9Z)n%?���n�wN�~\��9�����7���S�6U�&έ�)�Jh�����1��.&�'�6�Y6��&�ff�o�`L ���E��Qjǀ���֚F85~o�0�]�#��w*����Е�Q A��+�%$���ww
�kJH���Җ<g�0;�����gp-vۺ-��6�bh�vt��o�smK[�����:#�FG�-ѧ�_#��NXS�"�����~��!�l��1�荩��3�$Ų`��*},�>��ڋ�ҩ������ku��:� ٹ��Ǳ2Ti����d.�"kYX)3Zh������5m�5����g��O���<.d/.�:K��A��n���b`��~����OuW�x���:�'��=/��7��g]�!"�6�Z�������ꐆ�Wީ��~~\���(@O IAݾ|X@���T�D
���4���A�g���mꚇҧ ����/��A,YZ�v�E���,U=k,��R�>� ���8*m@?�X-�[���z���u����~��~?�hͻJh-
Dp�e{�x��M�GLM���+��GP��9��
��ڃ�>E�9x �v|���xTݒ����;�!�)���N&8��^\��{=V�5N����ߑ��-h�U�UpNI9��h���q$��=�������]>,o>0�}�*�uI'�&�jH���g��n��s�˯�ԻWF�d�Z��F�+ʡ��eH�pX2�W�τK*HQXh~f,8�/@��2���A�(�ӗŷ|���^��3c�1�H��rS�%�n��rF���
t�(?�L>�Y�~s0��\En5~���k���1�yіH �a�T^�4]!! ~�6��/l�:?H-����W*!@!���Z4PO  ��IDAT4��b��>�,ה0�4"��������%ݟߣj��J~��5���򹉤Ƙ3���t�_�\��{#�!$e�f3�ȳ�V�x�N���mD;���ڃ��n��{_Gz�H�Ih�UŴ$�I17y��_��^i"AԞ������$�jw�B
��t���w�Gf\z:�ب����q(�6~m޿$-�z��{;����Ԏ���$���MdD-���8�j����u��e��e-Z���orH�C����;�J�3Bl�-Y�%����˘QΐM l�)İ�^|T�۶�J-i{�F�W��gu7}'����6D�lJ(ҭ�ʁ�a��@Əz7)f��X]�����q�ŕJ�5���w���f�r^Z�F�B�8˕Ʃ���B���qJ1���l�"�][wVq�����q:�D���S�V��6�ҩ��yu��6D��@}	Ê�(M��ae'Fa��h� �B0F��6jQ��(A��^�}�ot x.|���w����~�>`���\�;� �>�j�?,Y�$)��Y�pQ	ՠ-1�g��-�j+�XF��$���1C�V��}AUC��
4щk�t�\����Д�;��������G
�!�`_Ȕ�ǿb��氊�#nj(��Y��׿w !�CW���+ia�X�k+q?ʿ�b*��T�;~(�¬-w�)J�;�N
#=זRϰ9�7��n�����X �4�l�ou3l>W���v�z�̶������׬������#�BhY�W|@����(���m���Z�~�#�y���o�9�&�6W:��:{�� ����u.���ߐ�k6�7S4I�c�&[ �P0�'�v$�,�Q=���`?p�>�S��^�͛����A���)���Q�A9)8b
��/� ���ܹs}����h��沏�#��z��g����-�b���ܗ�a�i}�+6W���&5h#Ӛ ��XW엷<�"F�)^��9���Kbw�g`o{Š|8�[��n*z��b�>T�k�¥<&LĕpAQ�9�u8���&cxBŉ�.�kM������^]N��k}�����Q3�S��:i��I�W�B(�����-nm\�Ͻ5~mw�U��(JA���u�^+�{ �!%D�S��tj��.�me;�74�L�9FY�k;��uxC�~�A�+E��-/��r�X�W�C
^W�
�T�.Jz]|+H }�/�?U��l8[p�b:D_S+��Sb��{���&��Ը<���˿FJؔ���!�����ƦV�b�ez:}pg
,�e
�(���*���NS�SU~9����e�w��s梱�����̵�=k��~����}#�L{�V��j�(ҥ*S��&%d�K$�Bj�f"��=��1��L�4)� ���/��t��<ީb�	�����T(���M<�n�U*�N�9\[��g:����t-Qv%t���S���:��>�aa4 ����5l��	]2��Ҿ�E/����=aW��5q:���ts��ƴ�����ـ����T;)�&_1c�Z���>5�vmԻ$V��O���&.�2ne]��!��4����=�M9v'�������.X������)]�ǡ����������\�u7\TA��� �і����g�5�ds��qb�t���R��VGˑvb>q�"ԃ�ʏ��b9���VWU�����"�}��R�B��=��@y1�iB�P�);� G��Vvk�jx��[-r0_rMԇ��R�x�5~iK�?֜�
�\�
�����ۜ����hMF��MQ,��Z��	©��)%|C�+vkUu�4o�����t��v��5��3�C۠�~P��oB��9�6�����hڠ+O��M�� 6����O,�.)<��G��g(%{ `Z��V���l4ib��S���>D�PE$]]E��(P�4ΦPYP�74`D��V�v�(�ibbzT���Q��#����� Ȍ�k����nZ�{��O��W�H��jNu���Q������^(��dr�����(ɑ�*+�%��)�0�lo��%���5+XB�}�)L�_�)�$T��}�"�cly����a eV���7J���4��h�S}w���AQ�r&?+)%��:Q����(�w��^�gڄ��mP��k4��e�`�c�nu��y�D\>��,w�!J� �]=-��鸺`���JM���ѷF���`«:�Vգ���Y���S%i	��ӭ�a��j��0��t��cS�Ȣ��OA�Ǻx#Mی\�G/���0d��.��<�\y��U�C��˳)ɺf�U3kD@�n�ѹ�����);�6#-�Ƹg��
�� ����͢b*4c�����1nw�gbF�/�1�����Q�T]^�A���"5M�@�` 
N�w���� �̔R(��΁j�Q���FSQ��x2��똫�cB���{�;A6�ea��6��h ���	R�Q����A�Aq�D�	��8�ι�J�K��1��z�f�@��[B��☰��ny�70��Gz�s�"�
O��ĵ���q�;|��Lye��#�m2?`�i�c��[�>��\#���&О�:�P�{����`"���Of�
ZL��G�������W�\OA�?����K�fa��(塬���L�,�O]��b͢��*DIcR5�d&~��S0�l71�d�UJw��h�� C��J.
{��suQI�=s?�������@������k�qJ�^��k��'�������%ۭw��<C���~O�sN?~RR�0���J�I�g�������G�q'3XCӯ�5.��m!���ۛd��T�¦*�am�"�.\q��!L��R��GV�Y(�C܈.�.t�P/`98f�)����:d�vwB9�����=��!�NZ���?�0�(�����\*��q�pv�G�4 �<#����<�F��� 1��K\	��
9�P�v���;V���G^� �H�o���_��1��,-B�Z����F@�=���cMWvA#�����
�!c��ǘ�z���?��Bt�4�E0����$�+.�q_F���y@���
��R�<��Q���w��:#&Ã�|L�J��x��C!����>��a������L�׏��!y�1_R
�hzGM�k�߈����_�$W�)Y���i%z=��_ҿ�#M���Cv��� Ӳ�M/� Kk$�`7��2ڣSq���*�zJ�y!0��Ƌ�皘�W$r�,��b0(���s]���_ӧ�z
��{����O�(K^h�$˓xj�	�G�+�l���6Y�a2#��в9X��I`�ؖ��fT�}k�ܗZ�	�����nv�h��u~0��!h��M�����~���$����"���z҆-�=e����W}vh�ה�	eWn�����������_����,du�����&��4-g�'���%LA߱�"T���w�"�6E�l1Aq���Rc���L��������=�ǿ����CA�#ݧʘ\ŭ��L���j��V[ ���[
��?�cMD����xH\�o?����%�1>�:�&��s��X�nA�H����]R��ߌD8q���b�b\!ަ�E�^���f
�i(��B��s/��=�J��i�����~�����}�9^���߫��3}��Oc��R��ñ��*N�}DV]�C`���T�c����4��M�����߳�t��XAz���9�v�*��(H����%��Z�1��u��t���U�Tu�P��\������w�	\#�+dK�h��e!N��%�oI��������ӯ���uo@
�M�k`t�R��ě#�m֔�1ӿ�J����d��B�6�,�0+B�������]��&%<-t�ђ�nV�h�Ɛ�k�������w����T.v�[�
Hؘ�\�ob�n�o�@��$/-Z~�����=��)Hˢ�ǯ�P��&�hّ�]cMX ��B��q'N6V��@�[GA���Ҟ�����*��Xۯ���!��_�*�ڶ���#7���g~(��JQ�"cƝ�Ch��hu{0��_$��L����Ep"��E�\�˘�����<I�(�tAK�k�2uMz���s<�#��\��j�Yg�_\�*S,B�_~%��!��|В�����R����u��+��S���Ĩ�M���^�t.�Q���\�ʚ+\hɷX�<����� ,�n��-r ���}Fh$uMum̎��Ż�<ڠ�1 ')3���C�r�Q7�X梨�*o+�=��L���tO?��1~����[�D�a=Ck�^4������n�J3��}���h���A:��چQ <A�ݣ����2�h�_�x�����B��if�L����Ί�w��q�k��9���e���(g`ǝ�k��s�nE&-<�ZR��_D/��\�.v�k1 ������2v��L;؝�H�N���@�a�V���:��N��9;h.d!Ӑ�*��-���c��g��Q}�]_����{���MtF�����A���
��*�A�&:�))�\��|P����W�# s�-��|a�	S�Q��){�|
�� -D�Ǐ�8Ayq���%A��@r��R�4t��}�t��t1��<e_i�R����2׿�V��݇k,~G'�u�%���Kr�	����H��-2���l�\�t�D�H�t7B�Қ5{2�j�φW�
F�k^�H�X�dq9+�If.k��_Qm3_Z��@ї��š���{\�S?E����=���z�m�Fk*c43�+�Ҝ)+�˹,��X��y��G���7�M�-z0#fWDܭa�̍)c{���nq�[�;`Q�ss&Z.% ��w4�oVt��2od�ם�>���^Ǆ�r�P`�\�v�� �����C2��I�;V�7���@�Թ�d��` HcD�����
"��SZ]\M]���Qp�]�RIK�3����!�/��m.�E٫Zm5��"��$\�^ebұNc8���b���3���@S��l��"���$̫*B\,�Z��x-�go,�(�)�NT���J�,�dǠ�'�˓��k7&|��h��,����7Ӹgű�e6��H�<eR�1;~���^G�fA+[f�U�zc�S�!�����R�<z�&5\��2QY���Z��;ؐ_��ȁ�Mp=)b<W}�	�$_��R%�@ؐ�Lj���u�� _o�q+SVԡ�2��JAuM�K��+]����I�=(7�6�,�H�o��-��c���L耄l���f;ƶ��zi�D���1ʠ��\��`Q��SJd`"�@����@w�����A�l*+ #��Ʋ�@�\��ߵ�04�fc��V�";LQvaDp+��$.��r���[Y��Mi�q��ꎂc!��h�B4�1�$�Ն�D��s@�(�FaU��1�qp���n�ǟ�|�+[él��niVi}+�9�t��Ѱ���6����)�����q�Ќ��"Y�a�߁�گ���̹v/�vg,kp�����1Ns]S�E6���EQ���jp42�Y�R��>7YD��>_k���5�U�\�-_%�N5��r���{��a�,�hԜ�E��>o�׹ø&Gwt.�4��|�� hƂ~���b]=��TJ5���r�Ӝ~-׷[vS�1�.0�3�ͦ�7I&��$�!8�Oט��=*�\��c��� r(�c�'��,�^�����^��'�^��Q�+M�z��8.�v�P~�B���\2_%��E�cW֔؝�$��$�%�2$s%�B��3���<IՃ*�[i��(;47�B��T�oӗw�6�&,P�1v�bC���HD�=�Ft3$�L��e�����Y��$��=i۝��C����nBԖ��f*빪�:���]��%""�QH�A�������Z@Oc����bTG�=SD�B�7�E^�oФZ[0��E2��#e"�Ф��
@�=��p�pǼhl��[�J[��D�U1,�y�NМd�a5��i�%v�k�Ȯ�~7���Ԍ�:�ܦ$C�+�"�c0&����N$�/���򓲾H�G2Fi�$�A���a?�P: Q��F�PL̥
�Of:K�i� 2��M�5� Ub��@�wk7�������W�*��f��j�r	�G<׼i]����������h@G��^��k=��Ѳg9�k��Ǹ��u#}�]��$�q	Q�N�4C>('�zV�*�A�D�RK7��i�Z��O/�Fp|CZ:�^�K��@r��WT�-r	=��b�;1��{(ㄪ��3�J'|�\RA����r��i^Et��z%�k���4��%�ʐF�^�-�rZ�X�}P�Sa�=Q}ٲ��|�xT^~U�9W.��B�K�,N����d��J���P�7	��#b��\|�K�'0�O�@yPT��z�����e�:O�v�D6#��}Z��E ��Bu���+��8b�)�h
�g������Z��~<�����OWY��$��,�	�4�s\9\5	W`w	���j�첡\a؊<jS��$�X�g����m�7M�9�Yx��2���,��
XX�i��Bꮜ%wJ����@��+-��w��5c�5�j�n�JS�\(�R�Ր��%d��������}���Y�rb�	� ��ҫ$H���HC<C�r#D����������&�~�dw7(F�9�@�/VԪ�*�E��@+D���6����_���Β�%�tNM�E/���o>�FsD��:���sⳜZ&�e�/���h�<�u�����Ѣ����F���,�ˋ=�&<��?K\������9�$�e�&h_Ʈ4���G7�B���Ԥ��^��g�ޥ~��o9U��5�(�B�_ǋ��:C����
�YW�d���m~�!ˑ��%�<%�l�φ`г�h�*���0���/.5	�a�Ze�����σMAF�30���#7;��L������u�B���V��FLT;�2�z�H�J�<��uk������Z���5���Q�-�� �~��t�P��5�D-�#��b�=�X���z��̬�����
nQ�ړ��S�%�+��Z�v�E�\�VH.��@�ړ5M^/�>MU�KTv�Asz��BN�BcYO튂&t$g�~B�����a�gpJ�*��m؝I����%

��<5Rm[�Kur�Z梏�`���l��`�Y����wl�����,H�e,�c����~�1c����gz=5��Xp����%ڍ1GO��A��l��@?�U���
y�ߛ��М�R�&�{mA�iO��rX�����/�ޞ�&�.���G$S�%�aT���`�(�]B�)��]/:Z���)Ҙ����h��?��̫Ԑ.� ��o�=Cd�yAe`��݌�w�Z�s�ua .n��3T��J��� >Ҝ鱇J�C���*��7�ͼ~]�x�Y�I@_�;$����(3�����X�HM�p�Q�P�k$$Ǡ�����8&b�}�� em֌��^��	������E��`4�N�̖�K���?MD�3�A1�}[> ��)N�T�JVS���@�W}9#�হ���ucx��k_>H5)V�\��-��n��&.��8��alG�X�v��qB4f�KI�ث���ɺLN�Չ��2�>�s=����P��ʛR��1n�&��eY��P������Zi�ҕ�e3}z2q/C
��/�s=\SAR[��
R��$O�P(V����w��0h&ϖ�2إ@ \;@/^B�M�ͧi�6�a���@�\��`r.P��X�%b�W�<g��E	���ϛ�����j�sn/��,1�^��MV��|i�28��Dr}�ݷ�*HQSL�	�ɖ�3�#��bԍ^�L��0�Г�O��ϏG*h͂�X��ٛ�mѮ�;��(]�:�9�Gs�.�zE���(�mE.�v� ʗ۠ܗ����۶q�נ �0�^#Gu��O����s;;�#�=R�:X�`k%�~���D}%AW�+�`�ʹʡ0��x����긟�o����j�NC��J]��W�5G�8^�Z?�!��)v=A ?�t�#����7�YI���)H��*��CM^����+�+\�/U��(��y�N�N��Tq���Y��()��h��B��!eDf{m���L/�:��]�g���M�C���?T�`��_�N���>K���q�L��*��J�>��h�N+�پ�L���}cS���= P"�������M����hXa5a[]/�9�r� �x��E�b�Ο�M�3	'�����k�U뷅-��.�Z�xU�H�H?��+��<O�B���V�C��ZCcp(��]����)r���!w��M�7*c{qj��ٖk�A�eTd�}���F~a���[��<q�v��۸�F�3_V1����zv=�tzS~�8j/5��JfLm�=��L���~�+�=gc����P6�|9�H$iaQ� IvO��|�����)��B3�Up���25bR_J:��'�C��������Ȋ�������F������Q��#,W�K�KI_ %^+��-��\�z���e60��q'k;)�j��]}�E��#52�^�������)�Q��i<iΰ�k>�SNR]���]��5��{ R���
)ER�^R8i��Ul����c��I�8a��
��Ɖß7u�"U����$����n�%�6��"B)��LLo�*����:!/��!l�Iڶ󴥁ʄ��V�B
T���H�c?g��oGU��Ou��g3�ֆG'��A1Hې/RPTyhߦ�����f\Q�ٵIj�p=��̟�e>���!Q�:��W��?/�Mд#��Ӽs0#���%H5x�=U����+j��*�г�l��ǐ[:���e��6#��>���� bb�tV��F��hߡ��.��&!͕�|
dQ��n�����ȷ)�ŇT�{��G[��_tO!˷���M�zc�Q�-0�]�(n�D�1}h�R��+�MOz0<�T�,̏�>��%�=��8b�x��rg��MöL�Z��E/�мg	F�Ӯ���Qc6xꀡ�-�����F�C,_��̪���d�_�
g��#Bl�ZT�Nfd��Lp�--��g��K#*5���6��^���]�()塰�v||��Ki!ig����s��ګT���F)�xTƎ��Ua�(�"X�ѫ"��m?RP9uN��?��2Ft!d*�CG჆Z�v�pm?�0l �r��	St�Gۜ1ɾ�k�&Fbl�8 MyO�nI�YV<��\k)�����%��
=S���2v��Aq�٧���e���,^!���[$�ڒ�7�N�Pe�0�Z��S����HXG�z
R/���k�P-"S�a��A\�S�Y�:H>�޵�~U���B����� �C�H��
6?Y������y�4Dt���� mũ�If��<S9򂈾���
2|�lI�V7QL��9�u=0~�İ�޻�����o��Yp���s�l�E~	��vuN>ˇlٽ\�%��u��e^I����ײ'Y������NWx9P�OD� u�\ڰS��w���V� �}��oɞ�!#�����j��~���Vb�>1���q�ֽ�}�"#�"ߊ���%��S�q�l&*����El*��гX�gK����$DP"���(
_�� s�}��4+�:9v ���j���iM�n�n�V���F���o�Zm;+�`�k��g��i]U���DBK������)<�}�ޠ�1��7�"�@��K:�Q������w(��N������<W��˯�T��Y��=ؐ��t#�X�=BO�ٺb�a/��l��or%
�SH�ZT_��=���]p*s��+���iڍ����6M�j�i��)��Sئ�kq[b��C��m�U`���׳bh��,j��R!Ry@�uE�o��I��և�Y��.����~xQ��5̗��5���Tݤmc�d������q��'������$yZ[
SUNL��m��J����~�
p<�Ӂp�sQe\Pj��
���h3`����Ds1�
|��Z�j �|N[`T~��J �����%;�L����;��Y��.s���q��7��-[�V��Ͻ!�6���16}�uxӹ��?$�*�Q��O^dMi���\�"��Z{�O�\w�j<��Cؾ�ig\�Uxd�W8�z_�W��4f)��.�-�2���`��{n�ޮ-�5�Z3�ޱ�7�EOݔ�#d�k�B����{�,�?�(����f%�ja8�fy�����$�����D^5Ç&L��pM����4��)��4$�a*��'^b�F4<��"���
}�)�[�r~͏�2Vb{	���G´��o��d�w��$��#�`L_>�m������MgD���A�����l�[B|�+�Aj�G�����ߚ���r�婝���/� w��LF�Ĩ�<���E�Y����|t�,�%�=�n����v7P�l?������n>�=�AN�������?��b�)A}1Կ�f±аE���bW�ǻ=]#���(�˟�[�SN�:�K,��p�������wvk��py�7�#�p6��d����{�rH��j>D�̕��Qw�ֱ'�s� ix[��ٽ|��Sˇ��<���Iu�5������Q�I�JUI�䌉����|RVE��t?h�餰��b��ոD�DE��l!gs;7#غ�����n�+�~�zk�ܻD�-��Z��y�9O���)H��<��,Κ���"b欅<����v
�h�	�G��>"}:7���@E4ru�J����I���v�B KF/����F�h)�B�'2X�$?��%�砖�ԤH�ڢ����-�s��(X����D�|���?ò]@A���w~,0�guT)�����r��|�QQ�'M����^��T#��WA4ͷ�NJ/D��ٍL�G��tX!y������u<�{譏��%Kծv4g����&m �k.&JU�-֟��Pg_�˴���
�\�T���{�,�g����)5�>{����LOQc�1��DK}�ʗ3�8F�(�r����#p=s�e�[�W���=M�υ�5�Mq*�&�XV)���n	iw�g$�R��&6z(�P�#�P�9�J��`�����sX�|eQ�u�܆�ڙ$$NR�|�Q�u8�N�/�\�{t)���H�t}=��V:唗�J�F�$%�K[����]y�֏�L�^�g��r
�wz�ˋ��i2�e���X��|�����듩O�E
Ym�~�$��sݴ����cwG ���uT-�;�q-נ׀��� }�hlŸ@��2��_�^�/�^�_�,a~����aآ3v_�.1�[o�A2c�UE�݃e=%��"����S���7�è	I���:��浹"8�++���2hh^�7P��z����y�mw��|8������ny'k�S)꺉��tNކ��y1h ���SNS��=�P�����o����8Ш�
�)���$�K�剟�O�e�fQ�ґ�'��M��h�k�|���4#��ndU4�Z�{�ma��� V�n~#�vZ�ӿޡHoC'|ö��w��S��ƺ�oY/{A|#�)[��@�,�������PU6?�`PS�AD�B��4PD�iHsbec�qg���-���WtZrMa��h�ϵ�' ��n<��u����eX�n�:�~�r9>#	z���+S�ۂk
f�,�N�ʘ�8�n���~�Qإ�F�8��>�{��i�xx ��x������}o�kZDD7��ґ~O�}ޥ���Y�՟��*H���\X� G��g?�ny�b7�Հvԅ�1I�m�+\��k�m,���O$r��-c8�ߚ�S����m(�+�������(J[�$/�iv?���>Xf�gWY+��vY3�rU��ٵϚuUdFsBk���L	kc��飴�(+:WO?`=�H]�'�`d�<�����5�`�LM��f�0?Ң#bP�MS�������Ź��~C�T�>�dc	M;�ѫ�R��`<�Xmi�(�(\ӃJΞy�����
�� %X:�Z=�q�Oz&Ҍʊ}���zGBq���u)Mި�kc�g^�*�×S�6�:D{_aF����ǈ	��K�o�.���|V9B�AYq�\o�05�G�����F�*\e����ﯷ��e6x#2J����QK[�
Z�n�X�G��D
�@y	�tۢ��rf��z­������"-6�xq����;�[���?����ե�t%�x%i+`s�v�����Jo�F&Y��c�m�#�qM[+��:KޤwC㪮/�k���F6��Q8�T�zd��Kc�x1� �3�g�7?�p��g-Ğ��v��52�j���0��0�a��4�mTŭ�L6ϢX��D��_+���ǽ�څ�%Nzx<��|Aẵ�.}ϱ���#��i��D}�i��u槦���[���h�5�D�Ej�~���$^�$�=%�����C;�$��8�ڰd"��V�K�ˀ�n"��O�����ϐծ��k���՛}Ä��W��)H��T�4����<�5gXz�ѭn�ZXݓקEy��5����J;	�>R����&��p*L�����0�o#�'>��;u����y?��bXw��~�[�'zu��4�ނ�[�V���aI[��ㅨ�����]��?��D�us>P_��� �i�T�
b3��*�Tt��ޭ��K�dAV���4c��	e}8rn�=�V�)��s
�/�Zѳ[�BI��~�r����D���ryH�3ZG���;�E�9
C�%u�Q�2鬆ʚ��*�&S�E��s��X�����8��fT�N�;��c-��f
����e���kT/[���}J; ʌM�̌Y�}���<:�A�%Q©Os��M�ɼ���hw�z7��-rb���q_IGkE��"��D��3M��d��$\NA�W�����{w����C	J#`�e�C����
��=c��v�6��j�4%�����]�9����� �24�:\�C�Τ2����/E���Rz�8z��S�0"�?{��k��ɳ(�Vf�wi輈�u��ʖZ�"�o}��^;�����~�XwT/$��lRck׊.�5�<8�|u�:m9����w��$ ��D6�m��@�:���^]*�h�nZih8]D�Z�F�;�!���;�Y8ֶ2��5�9SC�\OA���F�=�B�P�F�8k�]�n_k��s�u2,�E6���v�(��u�i�r=��Fg����>>QȦZ-��5 ,i[K��)-h����IE?\;m�bLG`�Թ���wD)��c��H�`~X�v�M����͠�{;�?9}�l�C�$uWw���׺2u��٘!b�fKC�G�������g�W�{�7�{��m8��.v������\�쮍��$*?}����ZKTt��H����v��-���O�
��b��u�y�q�" �h#�C�y�X�z���_�$(�s��s���~c.i��z��n0⢩˚`&�'
y��(	����#�ER���RlIߜ��������u�G)�[n$�����%3O�$Fy��~�ƅ����6����9���\6j�	�x�i�΂�ǹW�3w�ϳ�o	��O���³��i�ph�(�qB�uBz^#WDtk�"�~��^�ښ�o1���,�#�,/) 튜�ԴG��_NA�tם5��7��[`�SU��J?ڷhק�(Kc�L�}z�1? �Q���������(ȃqCH�6*C%2?�oT�H+I�ϰ֟
;�;�f P��;k<���T^c�ªtk+fI�:�4Vv��mou�����@�\G����<�{�z�~�<���2��t�P��%)�hgq\e�N�O��y�Ycf}15J�?;�_OA:�v�صHm�YZ�ʑŃ������'��Z�F��6�藳��"�j�������^��9�Wl$e�vk�v�:��c����L��ַO�9�~s;���\HTdL�r����/6��Ca���Õ��CmY��,��Y.B�poZ��1aZ�<ɀ�_XV�y�r�ݙ��������7J�`�����
8rIi	�:tO`\��=��\o��F��5��#�����Ʌ��"}[~��V��{M�C���ŭ}������h&;��<f�Z���w���Gd�q�ÜG2���w<^>s���]1A׼�3q��_�]I$�"O��	�Y�/��{\v��Li�6���d�{�n�u��.��B���U��L�_ѵ�d^��pO7��hvu�8[Dޖ|�]�HZ��xk�[z�N�0RVJa�/y5�V��}z%e�:,C� Y�\�r����Q����2 �}g��[=�'�T�qJGB�o�'�OrKi�s<�%�/�]a�,Qʆ����t��3qiV�a��]�WA������s/=Rl :�{�"����\��׌��w�����d�Iľ(a���Eƽ�u$r�W����kCt�{gT�hq���@e��@����}H.P��-�Qt@���o�M��8�@
��]-���ѫ�	��R}Wa4�ޒ�j*��č[a�C�*	�/��E�Й8֖��`���yl���F��9>vt�T�O��Y������_��z�ՠ�����*�F?Ӭp�5�Hu`FIQߚ�j?d2�-4sKP�Y�z��v�mq���{��w�Mq�|ֈq"�~F&�Z���
��S����8�>�/� �Hk�X��)c� Y�w���r���zD����:�:��?|ן��eu��/ȴD{I����\�ģ�c�ex&@G9�Cض�<Q����E�J]K+�Tc�
���(���l`g���9��J��`$��5q�V?y�`�ml�w�V������6�*)}�1�g,z�7FAa��Op��K>����2_=�G��gwu���N����G�K�Z��V۾�5�9ZzI	�b�䞵�rhg]r{��ó�#����z�Z���+.	��u"'~w��!�3���>�w~��٭?��W�3n9�����.���g�Cm��a�n7E��i�f����U?����R������BXsE���'��퇰��hT t�l�@.��}N=�ky�0r�|%<+n)S���m��B�?)\RA:�����m���u!�������V/�C��~vQW�i$�b�{]�+�	gǢ���ҙ�z��Ka#-������⟙�5�nu�|(�r��
 �s���eU2)I��z��Vܼw��wi����7VI�Tۡu͆hg������{����ْ0���0�s�������{����V��	�h!}.� �.��2�sI�H�-p�,Ԗm��Ei�����X_ɱ�9��s/�O%�ً	;�>yԑ��:u6:Lw2�w���*C��g
��Ç�����+�m���C��ƿ����s���T�=k�'���Ϗw�}��xޫ�����q���J3���h����~dw���Q؟�t���;�w\�kCO���)���d�c�v�m\�]���4�#g���?:fP;&D351��&H-={��2�y��Sn�K��5b�E74�_�A�B�2��)�o�`�PT�kQ1��O0W,�kD�]�dt@���X���\lR%,�3��H�n�:$�Hptel;H/�gPrs�1��e��=2r�*�v&S�o}�,����ZD���WHQ�A��,��:��s.�"����tƲ|ͻq�V��
16�0\���7���i.D�����E�E�}��>�)��Y���u�}�Q9z=��1�W����ѳZp���j�\ᅵ�Y�C~DT��yԽ�S@|�E��T<�i�u�p=i�*�xK�ʫ!�ӯ�����y���K��EY:D��^j�!ɓN��Y�R$��<�Ze�Usc\�l{`�ȗ��N䀬����.^��SWX#���x���@��J�/g3��Ɍ���V�'Iۄk��Rә=[\#�(ru���߶xz�sI`�>9�3l��x\Ͳ
u7��NZΏJ�����9��ԹUb�����Bb�淴��F㿯��>��Ҵ�ȸ�����7��Vw�(|��J��u<r�������4����W���g]�*��e��p"q5mU�hr������z7�^��N�:B|y����*�窩��"��SOY��G�`��Ƀс���=���c�\|�ee�kO��	C¤foCL~����@(�Ԣ����sE��i�	m.;��)�w�U����s��Sn�@���E���8_OA� �a�������@^��}r����g`qDY��%�W�K�W�>��<�����V?�����YA?�0����?o,���afG7��k�y@♮��kߩ�^��K*��'%��\F�Q�?��8\� |�pO|AQ�r
lH��k��(�'U���x>v�_�'��=��AzP���������ie�S��L�G���q��2�Ҡ��oR�&�I�� ^ �{"���o �C�~&��q��f��b$M�ڼr��f���3��^�;���_a.� -������U�>��gdȣ�$E~l� YSZp�18��?�L��2�݋���� ����1����F�$�ɳ���A�����a��)VI�.,�=��x)� �ص�4"�aK)��Ѩ�ѫ]��оM���X	yy#3�<�MM�4�G�pPN�ov"`�zH��ׂK*H��P}�~;	��iA���kD%CŠ��?�� �i�=.��Ht�&
���bDJ�;h��� l!#ᴉ�v`7��
�Z�/����v�J%����լ��4%B_3h��Չ>1�T�T���G ��g� �PY*��0=�X�̹Q0��Q�Y��/�K{!cU�"��ax�]�3�k��;�r!�9Y�G��"+�!S�uZ�Չd�3��>�Q&������E���8h���{ڋ�~B5t?!��9��E�
i�ME��G�G���-�"��.���5��	.� i+���� ���{�����%��Ʋծ��C�W�	�0D�Fy��5�"p��P�	�'�@2��X�M��4^�_W��
^9�,wO_���E+//)�'��xc�O߰��*��p�2�g��ލ>H����9�q��o������
Rb�O�٥#u}q�cKB'"E%Qi��o��;"�0x�dx1D>K/^������X��i쿷���4�v�fٓ[����Z�}���@�����E;L���9��H=�������^��x;@��3�yO3�������hG�d�\RA�rf���/��EH�]A���	N�]-����>�y��$E���}-|2�%ӧ#�)�G`3�s�Õ����/��-�w�C�u��~o��$��޲
����~k<W�-�vqx)�Dܽ�ui��A�=�8��\RA�e$�H���U�>ÏJ�*I�/)�'ږzy����\�Û��-�nL5�ߤKVFN�3���MGA<�|-����r���߃oCTܐrh3�3�kgKv�l77a���W�_X�.tav�'���m'�v
����h������K*Ht��L�a�k��7l�]�Q,�+����ld>`È(�)ƍ��F��0t���	V٣O~�z�H��T��r��w�MO�&y��;/��[�R�M���U�u�#5̉��,�a?\RAB&Ɛf�JP�f�H99�R� R��~#$����|��<�er&�42S��D���D9ʇ�ge�ZfP�9��H�fMlY�/ƐI��f��F;E�?P)��:��c�wG��C(A���D_N$2�;�|W+��U�z[C�B4?���9��5��-}������,�JU[7��X�`^AT�}��)2�oUY��tD��tT�٬#Lǂ�'�����"�j��>��	��|n�h��.vN�c����	�w���MTk("-EwUydLl�>xQJ�۽�$hι/I]O.����pI��:.��^}�D9z���N�f����6�h����=K�g���ݑ��Z�Z섺n��|��
b�c�vw 8��o��s(���r
	�Hs�Y"��xN�2��~���U%�e%E�ߒ��p��y������P�Qa~����>�A�ؓ2|�{��l`-�y�-�I˻�����S>]L6.���r=(;��{*6\z�-�_�.��7Tؽ����o%|;�#�7���ɫ����~� 	�<pB�����'n���]�Ow��λq�T�x��@q��ݏ&~p1~�� /`G��Sc��C��\���J�����è����%֧Ke՝��%��{� /�n�Nb�BƷ��> v�E�=iSXxj?��3�%���[ٶ�<)��>��;�*xm����;F��s�C+^���ݯ�7έ ���_3~�>��qI�`�U�{g���o�0���)����S5��қ���ih�Z��cJn|�A�x�,���蔣��t�Z���cԣM�9݂�+(�ǀU�U
��Ț���]I5=�1�T}�Ř��#�������_A����$HLǱÕ�"�ւ�o���?��:�D�x�a�~WCA����v�*�le�1����Qߑ�=�7������o��%1�2��`���w�\��n�oB�?	6�~I��o�����1&�~Ҿw����%������o��6�LN5iݙ�A�&g�ڊ��*.��V���@���o$�:	���5=# ��%���{=�da����K���c���\���ۜ�H#�nB@��hs�=h�������t�8��d�zO|���i�V�����@���Ɠ�uN�3���S�_���ހ6iШɂ%���z.^S��2�ys�3tw��h3�e�f�2d �3��=�c{�R\�Yf���c�z�ƞsTy]=���
i��Ȝ�lZ��N�3�Q�!�՘��#�S���n~g���J�M�C�"���\q@������-�˃�*,�9����=�0	=u�*��7znq�zc� ;�_Dy��lv�J�DZ�"ΟY)Ҡǅ\yP	q_b��]��h"?|���ۨ����v���
5]잁`>�����Ӗ���ДR��P�����VЯ�S��F�;��t�� Z�-�,H ��;���6]l���M���x��+G}���O38�1j��j����-;k	wg�k� ~D�����Џ̥U��^�~���Y4��.�F���m`0 ڧg�i��<m;���w���]�P��F���3b��A2��Lk���:p9)1�l)w;��#��o���!
@��(��V�Yx�\�4T�� -z��]�}��碉����-M<R�e`��RFz�{����~������>���"���r��Ƚ8�<{�|@��|�xP۠���Ʊo<�]�Y{���5x�%$�o��9�ׅv>�1����gHy�;�`|q��8xB�gYL��>�u�|�������V>�����m�r ��E�͂��\(T�O�/���<���>����`�$Z��-�U���1�o\����q�s%&�ŗ�)H,,����~S���h2�^�"b%0�ʾgq\N�8
�u������Г���06+8ݛ�&����o��@��/�<���o%�όɚ��5��-��������F�%k2@ǫlz\NA�{I")-1.�����Q�\�7|�L.Q��	��=���������g����~.f3�P9p��������\�Kr�L�h����u��o�)şz8el�t���HI�,�z�F�մ��w�<:4�t����a�\�֖�x,�}���u�<|}Q`\~ɴ��W�y->~���t��Ud�<N@������^��_��p�����}]�!����2���_���T�&�vp'Hf�������~&%���feg�8�D��ڝQ�p<�/	�,�o���q�/8�E|�ӻ���ۍ�S�i�Tv'@
G:�Y�w8b�и�D���o�"���\���#�Һ�VǕI?�o�@�.[�EyM��O���)H̼q$���ږ�)B�֧kA�}��{IQG�jʣ���a�m+?�������UMcĪRO(�Fk�<N,B�B���������C��_4��c�wm���Y�����Z��3�#U���q��Ќ���Ɫ1T��� �+����S����y:�s÷{��ߖ��œ��iZ,���&Zvv��;N�*ƹ�����M�n��ŧ�ú���r�%$�!�>�>�L�[9�"�458�#�Z=���$�����8ڲ�q���٩]!-`��J�r\^�SL>�`�댖F��fl��7��[�VДtgGtC�:Ϲ����/|x�=Β�E�g����р���g�>���gc;�m�?I�������5�<&�P��<����|�E! J���T��p��^
���^{[�d�:@ք���͎�D���� x#|N������)����p���h���mؐ}�v7>�\o�#r��;����vSW+�2J�y����ʘ�}j�ĄQ-?z�;��@���eL��U�D�-j���!���ox?�-I{��u�;�5��H��hV�l_��.��v{5~X�;������(�i����V������8	C�OD�A)E��r}�W��v��+�l�M0�5ͣ7_њt��$����,�cD��ǈ�� �怖�;9rl0t����gr���K����p9	��G9�Q��r���E��B��|+K�&�4G�P�6�!�(	!X��ۦ�q�����W��eK2�� Mw!�< -�]���D�kc�%�G럯F�n*�6�?;6�7^o�Զb,���6[��g�S�m�_waaD���(��`9t8��S��zRKe��?߅��h� �5��![���dW�2R��4 G��J��Y�䆇m�.�OyE{})]�|��Uܑ��sa��6W%r͏�M����w��9�[z��?Ss�P�h�/�����6�5�E��5�[>|#ĲW�j�>�S�2��uK��e�=G�;1�(�gl/�K�ߋ����D�BM81������x��1�S�j�=M��e1-1V��(��w�J�n�4�H.:6�
���}�l+�i��3X"��!�QV\�����Fן&2�@z��rs+�2��)���,n���q����n*�\������[�V�u��bFN3�Y�=Q4��2�� �P,Bͣ��8L��i�e���{�.FCG
(iB>��L謁��' �O�u�
��=!���� ��<�W(:'Y,�0�p~u��E�V�!t��d��mN8�|d� =DJL�ǟ��;E�*9�L��zeT,Q�l�SCS��������
4QS�Ɍ�Ac�L�Oc(wsţ��7(x1/q^�*���o��#b*4I+@�u�F]�Ep��gt1`�%	�Sp9iZ�²�i�2�o�<t#8-�;����U����������������"E�Ei�$a�ᾞ����l�Bb\}�ŗ��`[�)M�U���B�7���8�2�W�QG���`wҎ��W���tM���G2$�����H���
S�@ҽ蝡��g}8�B�j�R+���dr4vI�}��}Õ��
�F�V�D6���`��J��OC��ύūv�X!2���{-l���F��B��h#�{�2}�_)��n��No�5'���m�+h&�����W�lv;�;i�V����=t�9|�������VL�l�`�+ڐaÿ��rN^���΢�uTd�M���iCG�����w�����Ȉ�g3���ځ��ؼAJ��P�7\ ,Ri7�O��$��!R���E��C�0��c�FD�"��^�ʇ>1�"�	����k�y��Brmx�n�&��k���!�Z�-���H@���$�e��W�F|8d��(��`h,v�헦���u%t�E܌Rk���3��]���g��K���}2E��X*T:)=g�Av�U���Knl�r�u��a�1`=����_���"�Ww�>��Pl$�f�yBy1�ۖ��D��V���_�K	g ��O<c�t�XMA�&䯟q�ޟ\�Vi�$�v��c�gA�޸���j�z��T}H^�%��r��Z���iC�ԏtA���aW�1��e�n		����[�7
9�EZ!hOߚO�h�/5*�����2�Aܞf���d���>�����K���`���m�1��h`���`4 ��I���]�]k��$h"�8�P��>��C����6�ґ�ᬨ���9���.����_]��L��l�2x��
=.� ef��R}^A
��/������w,�v�R���U��úP�)�ڴi�H;#�@'�NI��cB���Q����m=*������tJ����(C�F@T��; )$�;Qg®��NA�"�����{7ĸ���=Q�=�䍛�-h�DY����%�g��.i{h��a�u����	�@nG5N�0��,�+`]Y�\R�+�r �S�=S	V�a� 
�<�rl�j���/�<��,\� �v���8m�� nH�3��"4���J	���W��v��dO/� e��]�#*�-�)C���RQ�N��|b/z�cFL��%����Y�ެMS��y�'���E�a�b����lR���D���'��yek):G��X}{���k�)�O~v����H&C)XH[�����kq�ೖQESu��͉&$��t+)K(���DZ���f�fU-����e�JgHg�a���	:�ە��S����?�uJg�`���
$8�� ������~�׮�\CFk�k,BF�["W��w�>�#p4l�Bιp%��4z��e��H�j���B�\��kᲣ[��}/r3�����^ă��-�Q�lZ[E��5�*:����53-���nJ��e8�VA3S�+n�*,{}	�a�"��x���ښR�46R�H-�)�"]w`�>��T�if9a�p�KI���<(A�:@�g��t�ԟ	!k�gR�J;H�|�hJ�ȼ h�o�;�o�k*HT	�M�0�M�5p�8�Q?;謀�g�|��CcA��F�}Q(�l��*aJ�`�la�U�KF��_�/�����҉���UN��{r��~���(qԈ��"�����^�_MT&i�NB-.Ț�|�&�k�I_+P�P��{# ����^�)==f^����o��P���>R�l���[G��x��w/A{48bG�V���&�|��?�98�TV��s�=�YSꞷ�RЖ����LT��!8jU�X�_E9����f���Ʒ.� U!G+��9�}���3�&�>�d��jԤd��]���<'��X�A��9�&8�i�#҈�R%(r��3J���̯ 1���Ͱ$�j�]/v�Hj�)wl*㑳騀��ى�[�ᨋ]��d<�1)����VՇ�WBe�O����1�T	B��XXp�h��bH��*��l�q�~A5l�߉������rd]�I��eT�"D��-_?!{qc�����׼����v6��!r��!��I�㡨FY�:5�'�>	q��X���7��~�������.L�*A�����>uX�S4;pku�L����g��Օ��)�;b���5�@U4����� z^��}���`�'�����Ӹm��Ǻ��A����w�:�mpA	��'�����y���s��Cf0"�%˼�6�J6�j�Kg�<�3D��x!g�y��vA�`j��*i��X�p�����ɯ=6=�{�C�4���J�y�%КsM�?�C��RU�����y~�`n��`C�cn�5��W|ϥ���3�q9�d�_�W�_ym����ݴ�$���p���Z�����Qā��CtV۫<���A�FPo�Rj�oz0�כq,�_�Y��{W���H�� E�G�B����*{�����L&(�TiUao��y��)�Fu�14 �?�9��C�n��CDg����`�6�5������km���{���"����g� Z���#������;W7i䶉,��c�CB��v&���שzt�(N�c.1./�A����������(���UΟ�� ���|LS��~���^���DT�|�y������sc? ON,�S͞�蔣�Y���$_�$+�����)�bS��b*����e#�X5�B+GD��0�
�ឞ��ۻ�8uّ��V+&�>�k"�Ujv$}�w�QO��,+��J�1����dS�d�!+���5V66Խ�N�j���
��o�i!E�W���8�����He��(�ϒδ;sn�gb�!��q@��R@�(a��ش�����Cp�ٸ��� BЎ
��p�Z���Ŀ�|�ٍ���W�`*��^���v�*���g���wҩen�a�TL�����f�"��Ix���b�/�Y�����S��
�[9d]���_���q��Q��{;���EnT5�����-��1í]�@�u]�~M^v���(�O1ݔR`��u�b�U#��X<c~���9G��
NP��r��RІ�.F��;aҹ� �[C:�n�!�eh�z����T\t����*$�b�$���5��Ǿw��]~��J}QR��J�C�u
u�f8z⊓|�{�ꖈ�Y�5ɵq��Rt��	]a�D0�U�xw �h�\�O�K�vT�v�Š�J�.���y�(���(5��	�r�:����l����ΰ��l���d~�
틈|��7��]��hq���	<ZJ�=yf�']�Yg"���V�K*HHV,.t���C_�Ͳ�'�y��ՀX�#��'�ϼ{�b'ݶC�[���1u���%,�v~�W�,x-���6�H�/sܸ�����1C����QE�J���-'S�������tC�D��Ӕ��9&®w��ҍ��]�ޛ��bt)����h�_�D�+4d��װ��RY��.(F�����$r���l�d�sχ��D�R)T!�7M��-#�H�)��sS�Y Y"�W�"��v3Kn���6�{��"J���P�jt�,0.Q$�j�3mK�\��,���eܖ��9hʃ�C]�P-���:�Id�5MȦ�2�gfT4�#�!D�<��:)����ݲ��l�fA��6g:v/Blv^��ƚwv!���j���-&3�SQ�<hw�m5� K]�:(��S4��4��,�M��Dڀ�j��p+��0׊^`\���zEH���\JQ#<ۉG�E鵢k��v��"�,����.�I���׽�ӼX��(��@=ĠYX�F8�ҡw�X��4��{g'�SϿ��C�m*��`]Ae����S�������T��/@�($��T�Cg٬�����⾾�?�!Ѫ^�D@̸9b��]����5%Ȫ�s���TЂ(>�X9�m����Z���#�������䙎?s-$h�'��lkI��}�2�2�?oX�xq��mFh9��:;�JX��
��.B��ڕ��n[@3��f�מ��Q>cX��,pI4�[*L�9�,[m}>�8u~�Z8rw���Ui|HL�yQ%��$6~zGSPxa-��w/.�=G�W�ի�2���r���?�-Zc�� �]��ܧzN������gWx<~�̣�D�&�4��e<�'��$-���?Ȼ3�sn�`�o�%��}U���k�Wl|,]
�)cCT��(
*Q��,����Nv¡
��~>��D��4c{��h����]��E7*��k�2Ï�Z��z�H��#��G62Եi�����>�;���N��WΡowEi��^A��p��U����H4�'f]����`9����#���a*��	�+q���M4)Wr���w�l�h)��\Y'5f|��/Ix�(���!$l�|�,���\�t*ȅܦ����G+��z����]�歨�N�����y!�E'J����O|$W�ć5��W��M�F���= �$ޡ��g��q��*�1n.�0�q���A�b�����r���d������rɘu�������}�=]�`���Cl��-�Q~-�ٯ)�;�NU-�2�\"�{^�(B��N�JQF����� i��Jc�P�Tط���d �`��{�z�my�V�Z-^���V�雧������¡S(�.�ǆ�_�QE��]r(��6��lQ���?&[��s�����ܫtO� �0z�lÂ����rQ��Q���R�
�Z�nӢ����X��k<�,	��%�ŕ���Fm�X�|���1N�Q�����V��ӏG����ꑒ0��p~�ʘ����D�P�I�N:�(ն��}�����A�!t=����'�"�� R�����h��%�*HĩR��ݲ���IO�x����@���ߎb�} 撊q`e򠲇L�#��\ު�X���j[d�K��(�Z��lQ\��8?��_N��KĝX%�V}bK�M[��m*��B������)#)�\J��m�ca�+|�-VҤV����q�d����q�:�]���"ӂDd�"�r+�y�Eцۭ0T@�<�Xk��DA"���GPu��%Т��<��-����m���H����p��@�w�;&�B0�n�� �d�`Y�7�~/�H�J�\����d�F:�����r7W<�e�*�˘-��	��G�"����?�У�Z�ۉ1$��%<����g*���q��i�\qt��_~�_�J�����:�u�n	/�حcPqw�60����cԬW0�^����TJ�ly���~�]�oȖÿ(=�28�t���6��PЖ�SA���c� W�����_�h�����SGB�t�2��8Җ�h�D��.��g��"�v&�y���J��D�y4'��NI���Α�-�N��+*H��`���H�����\ok�E̷�i"�i���� �
�\�X�Y� �����M��Bt��@��I��	w��y'�^f���D�{(?��T���e[�fUe�Q�>4�^9�F��g��9����4�������N�k�
�±*
su��v�a	g��c�}Ŕ�kl�ê��6`	3-�dA$[`���#�_���iZ|��-E۪���z��Rh}��tGV�@��!h�jڅ���uRX���畞>���c�Zo��K��d��[�D�%�ބ�lH6��"A�*a��8C�k�,㭳��.y��=�2�~�oE��tZ���S�=S��3Z�.7�ݣ�(M�?>��
Ru-.���&��W�X*�Rj����M��{�kž|�#)O�3@5�d�Y�
���x������n�kl��Xj��挲����r���OB�ڣ_�c⊞�ϵb�xR�R�Q+)���u��ų�ϊ�<�/�,�ݨ	tX�g䖖8A�_;��Qƕ��/ �|��i�=h�?�����g9s�c�]�7�FK_��/����#&o�����ܭ�7a ���_�[P���������[��C�d�.Ƃ��Sp=��-���2��Њj��H06�B8��<Orx�. R���N瓀5�y����ھu�(�zd�#�t0�:'��_,t<ƕ���-�k>��u+B�'���]�9%Ƀ��^�|$� ����a����ŕ ��6;�M�"jP��*�)�8%>h��9�E�Q%���ׂ�I�����5!�b��-�ZQ)�VA���(���;��l��2(��jJ݆դ���?�S~���>h���K��W�r��N�Sq9kD��%iUX�j�9�tE���p���1Ǖ�E�@fΤ�m��A�T�Y�{�\��Ӵ�0s�U=uxǁ��nOX��Ξ Z��2�5��T���/�En}(�����:���|N����(e<�ٕ������2
-�I�4�6�T���k��[i�'�o����3l� �:�
���,\YGEi\���1fK�-��ү�H���Vq��tѷjm���hk�_5���nx(H?���i�O�?�`���)6hi�h���e˼�Fi���ߩ#T���V�N��o��_��Gk �B�M���hjmY�S�H{�Vdo�؞M�G�\NAZܬ~��Je(�\�솕�`�~J����X�V=Qɑ��Uy9xG"�ӓ(�.x��|��w��� 듉�ȇ�fa
�>ݾ�F0�C���� B�쪮&�@T�C��1]p���%ܫRHK���~�E<�h?���V��Ͻ�����@
�ˠO���$�@N�1�3���%�x|ty��X#�e���d�)�ԱelE��V�_��9Ydd���VӣnT�����(g�
�5��PZFv�?�w��wH�����N5|�9ó�	�Hy5���I�[*�:�x�1��%����}�;����;�J��қs^P�o��y�k�k�ߛh'��Qjb莵��J�s���R��fZ"bN����:}�y|o[�5�������|C��;�X�_W܁h��E���(�"���ڃ�,Z`����\W��5�K-·~_,C���.vh�܋l6�(Aw� 3?~���U-�n"#�Ŵ������z ��&�h]S�L����5�E�����3}.� -����̵Hd2�Z ��B��	��K, ����`x����D�}|}!���<��!������΋a��y�@���yJ*��;
��I_x)v(	|Җ�3�����:��K��3�)��'�`<���Z���;)�F�9���XCX��U��TA��*��狿�E@�nGfie-��V ÿX�L��.�7�RG�Kh\Sۢ6���.ƫ�1 Qz�p�V\�(S9�͇̔y����E�XXu\��b5Q#�u�24�\]�h�#4W6��B(.R���9��_���2Ue�vjZ����,!zXH��(��oĽޢ�w���0dݑwP�����(G��J2��ֽXFsp�gp'C�
���ϣ%�n����a)2�Se�ciW�)� sѓ͊��B; �8oS�a��p9i���Ȃ�����?��I�7P���B�
�"��^��s ��0�k�P�ұ���\�R7p.�=l�˙�,�r$�.E�9�T�FgͰ�d�'ױ� y��g-º���g��ƫ�v��[�Em��J�"���(���=Uɢ� $l�5ޥ�@�m[6d]�����_]�1�4J<V�L�u�����g����]}����h[5>����&i�ʧ���^Aϵ�!�4ͤX��w~�G��+�����bJ�Qʴ�Qǯ�X/Z�c�~P��<g!fح�.���xͷG����bE�j��\(HIZv��Xҩ��Y��3���N#X���d�H4�;e'��2|(`�	����}�n:��oK�lF����m�Hp�|.� �Ն����P~�H��3�Yc�����Dyǁ"�r�3�݂T�"[�z5��IC��6��h�,>w^����'<cQ �w�ԃ�
#Em��ȳm���-�{0�0��&E�i}���J0̺8�u�[֣��FO��|X��vN�&��+6�Ƣ�Z���T���(��������wCn��&���9�)�zGH�n��LV�v����z�nȐkk���G�����yFr�����}%e�����	Q�H�b50�o�|�\EA/T��c����"b��F0��JE�W�*���]������4ߕGxj��OO?T<�lx�s@�L^�n�Wb��Nl�`��e�ʇ��,"O�]�f
�?��I��ع�� 3��(�W�.��}Ԋ��r�ڃ�e\�z{_���(�$FPpݛ��>*�V��ոD	�&�.�!gL��J�3X	4ʡ���$]HP��NWcwog�����߾xzL�;�|�8������74H��%@/�Jj��/.v��se^�,�Z9��1f��'���?PaS��%�SY�nih`�=��Z�N�/�Ok*���Ec��n������Y��C-��f�$$��o�H���4�-v��̲�L����h?j*����Sz-�"��*t���P:�8��Ӑ.� a�M�����x����0��'�J��� I����S����k�����hd���n6I�Fi� ��4�2�q7�i�ɱ�tbA�|>M7(�|xX[t�9�N��l�VgtYe�m�F�VR0�i&�Jp��B��r���(E����bm�t��4����t�?u��.�Zūԭ��$��䙚�T��m.OT�ƮcꖳZ&5e.���(GI�\���A����)(gs�@%�y �i��
yрR^�>��ag=��tƿ���VY/�1b��I�r �F8�y(��
NuSfb��)�fey��\RA����S�O��n�S'�~#��. >�RZ+�w�nM5�#��IH۝Ŋ�5�ֲ���@�Z�0�~5�Z�y�����3�7��{-T��Zbޭ�&��,�O��s���P;����d�L�[��/0q���?�����>-�)Z�,%V��>����ޥH+�(���*�x\C�H�t?�v��ȯi��B�5���^Z'�A f�՜�5F$;�3�tP���F�`-��R�mm��K�����hJ�����U �a��!N�\�6v:�����޻hK���b�s���g�Hz$���IN��{��JHB\|�*�����e�;BH�Qr/����B"�(�#�z�YV�j��hi����U�l�3�Fe�
 ����r_{����igA8�4�9C��x�h�\7�ԡ_�j���B��Γ�:2��tb=��qJ�{����O�Ѯ�Z���䂭l�������&�|yfz��j��P�� �\�얥����SzXL���m�2���U�M�Q�R�ۏyCTv�i(ՔW���z��<Hz�o��C�nև�#���j���Q�Oj���d��??K�h:�0?�Dو>ܑЩ�
7�Jg3|�%n��u��ߏ&���ll	LF��N����Ƣ1���y@:��Ĩv�,��ҾhБE4y��2�Y��fĤO֌���n ��gۜ��%y0��)��U��I�-J��N@�ztr�U�l��*��ˏ�o�+`��7�^�� �o�KFDotn�e���e��:_��˝[p�ϕƢ�-��k����[E��+ԅ���I�N�I�7���֧�~	���Y	��6r�Oe����{:ȅ$Vf��*��ƴ���1[-��ᆼ4��j9�H���z��1Vƺ�(/��)���g��joݫIi��05M���a>�I�+�hǧ|�X8�{a��x~CʷJd�̾x5����,[��uଵ��n�j��o�@��<K��H|�I���,Y���3qR)2T�޷Aף�3bQٮ��&.4�z��#���ه.{���g���t�B��x�:��`��T�c���.�(��,Sr-W�ڙ�zͦ��tn魹���Z�ҷi*3�1��d2l�Ju�h�?��\�����(l����Y
��YHnS lGӧ�F	f��Sk|��e�Z��|j���.��Wf9~�l��;��1&T���C��ρ{�ܡ|�1�|�\�:��͛҄{7�|Am]���{������f��;��NIB�o�f�<#*��{qJ�w�r@�ٰ+QEZ����&Z�{hEi�ݩck[��p[�8�Ð�+�##�X%)|�1W9�e�yo<�\�j9y-Ę&�įJf��Py�i>��ؓ�L���Y<S���֜���V���ֳVxjڕ�6��R��y��nEmK-%�>��dN��e6�:{�<	S*I�n$���mk�S�[�D��VQW�ܢ�"]>���4ƴ*M�� ���J�N��E������p� �'�fAX��/�tά�}�^�J&V�Ơ]5Zh	}U��⟨>�*g��B�5ain곳�t������s���K����e�!��D�L����Ȳ�W9�:ϫZ�D���vY&�����v�d�8�R��}�S�]4�E�l�{m���2�#�c�v�w�	Z/�G�8���H�S)��4�8�rL@�\�QM]����ֲs��&<X�V�{E�E P��rYJ�rr=rd��%%��)��壱���,�NT�z5.�� ��_�O�͈��GVB�ķ��r{���i�B��`�&b)�~Pʼ�"_���V0?�vΧ" T*[Ҍ���xdU�;����K��*
���3�-:j�CC�(2 5��`,����,��6�Q��|���±�R!+�:R�7f�]%�f/�^M3~����m'�$�mNg��Zu�:u�� E(tr��;.�թT0Q�5�s���
�ѡK��J�|_A�hM�&R1~��|�t�c^���9��_���x��`��4��@IF�l�JM��q�I�{U��
�'�d���,��P����p�p�AH
Q��-�d�Pv#'4)����(dM�¬��#k�R�M�?*��Na�O��q�@͛���5��\ LJEx��h�[F	���K�kE�+e$�e�\�rw����*��E�r/��ј�Yw�VPGa�c{�D]&f�ø��b��3E�v�����aΟ���s��X�#��[b1'�ij�mm��*�IU�x�^I����z�ʂJ�=�+)�3���ļO�l V~չ'y����TR�Ebk��dNQ��u�5�c?T����"�X[Ξ�2���Q�wWG�k��*y��xP3�ܕ@�\��9!��d{h���5��r��rEo��o��������@e���8a Q2��_��ì�?~�"]4�\���#b��qѣt�j���ד2����ִY���6��5�)$-�3N���Ho�m��h��=n���߄z9�<��">�T:!E��A"&�3r��t� ҈"���N��/��������i��:�Wt�5!�W�r��/�da�f�$<0��hPy�)R���V��$[t����nneX���wd�d��}Hy�cR"��]9ޞq��Ls�P���w���Ć��sA�`�D�l(0�>\��;��0�{�ی��L�^���Ѵ���keޅS*HL��ЍH�Q-C0�lK�C�I�t�Šs��zO��:Ɔ��B#�(H�6�u�Ǒ�x��4�"��6z%�E^�{M֌U�]G�Kz}��9K[(sJ�Q�33=�([2�[ٖ�iqn54�ns�J��G���A-�&Lի-β��o�8�dW���P��x�v'�*�QH��iT���vju�%��&��[��|G�ᐅ���nF�M�����r�P	�o_��]I�]�c�w��x.?�3�5%XY��w��BY��y>vB᭄�F���Q���A��Ǔ|7MbŴ�T��r�dzOMs<Dd��Y��S*H^x�XQ-8��E�VZ:]I_8面\f����\�R\6L�L����;8HV}'��Y ��%�_���sm��"�M&b�g�Ε��:�F��V�N�|%�g)�|����8[�6���ߡ�^+�w��{.�g��4�\�F�u�UE$�n�	`�m-9�䵌��>����ȧ>���b��넷Bʛ�W�vs��'l�O�����CBj��;d�[2���_̃���~�*@YI��m^�`�[[�����*i�|�6V��UY{�z^��8V[���F��M�����!�}e��P�<��?��f�c���I�/��5�UPK�<��� 0�s
�d����R�*�o�	$L*HI$b�o>?QJ�5�?Q�bg��`mIo{7m�۬��w���⿩��l#�3�D�� 9��v~E)IP5),	k����|#uKYcMэ���˾ԯ|�����RT�.����&I�`v�vY��k����z[z�տ���,
Z�:�4���W�j��yX�96�2�
�Fk%VxaӅOs�L���Nj6	`��]��*��:�i��.��%䅧.y*��1x��ô����l�m\�����i�7?ia3��(�i�����4u��qθ��n�O� ��v��P}9F���u8�=�v�p酛��װ��m3�1pM�Zq'���3k�<�e$uL�da@���ʕ�{)�E/�o�"�ń��>�I	c�0���5���v��1�7���l �za_��ve}���]'c��W�Hɟ
NB��X�j��H3�\ځ(���d�xy���>Tز�cX���:�in����G�n�~�R�J KKjc3�`B$=�b�YT�Ltڍ�~����U�K���X��<��GB�!�{/:���K��s\z�]�o���i/��@zc�sk�kz�JSŹ@+�h�����ݟr���(/�|���7|�-�-��V���j�� �-�9��7�Ŵ�4OVD�['�<Z����� �Z)�U����{ ��硹���0MՔ�+@T�����iH'T���U�B<1��x�%=�)K���#˘�F��6��Ù�f���+��Ѱ��b����V��Fhj+�`q ����i��v:%{��7VaK�G�@Cb�pMEv�JVE;�qS:Qe2��{��_�S:f�{K"Gi����x���
R�c������bl�Ԑ��NAN�`���x;�l6gt��CE�J�ncF#�UHQ��F��I��	�y�n���Ak�s���oS:�E�4��cZ�N|�R�{h��Gk�e���h��>;����Vt��ck���<�yt߷�}=�]eNg!�%5{q��}�	G F��!�~w��=*��̺���̋b˼�|���#��rs�7�r[�KQS�E��ޏK(H�`����_9T=d=���hx+	%��.W��O:>�!6^����}H}7��ëi� ��)��~�ʜ�y��[�,���aΉ����g	f-z�L��������5�"H��^Ar���z�T�z��A������je_p�2��Ag	����5��b�Vۚe�S�Yg����Qe��9���DW�/V֧�Xc�$��gє�2g߲[ECX�f�{iʲ?]IRV�oտՇ�u��5'�������N4���N����f~����wG7����|�����^�PA
,G�p�K %�e�)ۚ�u)�`�5��Ve%0?��WoT0`�=s36�Ys`7,�~�H)Ӕ�w�H�Y?c,P������'�߻����E�,�o�n8#�W�Zqo��w�]���Z�y�2����~���AQ��.�wO� -�˺�A�CV���rD9�����?)
1Ce�����v!*��G.G,�y�3I�L�y��(R�X%LZ�A^g�ɕ�&hX�ԷV=m��̓,ψ��*��*Cou����T�I�3����P���5�9��>O}
�iS���Rʳ��H���y�,��F��PQΏ��S�]=~��k��+��y7P4��i{ήUO+��+���ŤǓ-�RA
m��/�u��5�	&�z�\4AHy� ��ݳ}�z�ZP�#R�4�	�$�������I<��OJN��ҙ�Ty���H��9*Px�{Cj�	��Ӷ�����x�n�YYfӪ��R��� x��6�!�񪹈�r�M�P��\i�I�<���T��
�@��Q�7�_��+燑~��wC��)��g����k��v_��o �Ɛ�}N�x,���=V���اT��b��vfB��p�##�u��0��W�?j\]e�xL�4nQ�_dg�)&X箭��}��B8��dVc3M� �&g��![ñ���_�|j-6��X)��w��S�5��C�;"xE��hy�^�9�"�Z���g��P��<�Ek���.(y�Pj��n����'V�,A`������VeU���d�A8G��q��E��M/^i�y�TvB�=���<Y���=���I��(��^��Z���5�~���wt֋��B�%h������8l�W}��ߧ�ZY�.�<����B['��E�S�T��؉�0�5���
D�L?�w,���X�'M4]�:ߓ�6�塼�r�&�!Kk-?ce��t
�.��[��F�p�*� elMo%���]�[��C	�û�!Zۓ8KW���n��{IZ��oP��\V��F�ͪ���䣭+K-���X{1Ϲ��y��OOm�/�Ưw��
��1�8mr�Z�d#�Q����/v������/P����CiD%Ʒa��ҙ��*<"X����gmO\LV���6����eK/��W��q�p?0�[s�4�M2��)�D�����K�1�jO�U��0��\����k5Efr!%�a�z�VW���1��8c�Pzb� �쒋\^nn��)v�s����»����>��tn��L�ߛ,ӱ��i6dv���W�1���&,�����>:���	���V!X�xow왧[���T�9
nS|��n�$7�s���'��UZt�)N+V�j@ՇͰn�������z�։�X�{�e?��d���*,�w���!���j()�ϟ�	�� Ki�����*��7B{}Z�g���{{[iɿa��l��x���|N�1��K�Okɹ>��#��]��6hW�OB)gf��~ް�ǘ�8��Z h�Ý
R��4��t#�$�oP�n|v�-G�i�s�������q�����m|���g���^�J˨Z*��e5ޮ<�ފq�F_�%Ⱥu5�A���ɯ�����K�7�B9����{b>Em�Cg}
�� ��%����}'!��V�߁3�B�ۘi�h^_�ƃ����c�|��d�� �U��M�_�j�ڌ�g�V��pڍ5]ȋ�H��Wn�L�~��֬u%�#/I���O��;o��(H��yP��;t����Hn�	{i��w����(i�<{��GWL}"��4^�4�1�v�H�Xy|"��bt+���0����7�6���y� Vc�|�A�C�FG���ŭ5W�t�5��·*Uath�<�:I�\TA��@����F*M�^qC'��������a�	{[��Mk�j+��`�'���HB�����W;oEFwoqz3j<؜Mtcv�����C#�<g-A6�9'AY|w��������U9?L��$�� �DN���[��$]=��3c�+�W�!py��%ӽ���d�W���r�]Ic�1����|�}Ÿ��t�9+a��\�n�_����j%y��p#bT�}V���$�V����2���@�;�A�oE�����撼ǐ�,Q������G#1:�ǅ?�7�L)Iv�<7 Nx�\�m���d�__j��J�`K��Oo�Å�
���v=u@����p�:z���A8��)�Eۣ��K
�ߊ/�S���C�vˍ9\�N>oƵ'�'ߎF������B
R���Ԥ��$�1�pKQO?��N-��p��ѥ����B0W6�sW����P�Z�-h�#m��!��b��z�UT���+IE87n���8�hIPc��f�M���876Ŋw�(OGK�o���ݥ�Z\HAZ0 :����T7Bګ����h��T� ��!�:�x;Qc���Ӎ�aՙ���%�'\�x�uH�y���F_
�n`0`M{~�s2�)IW��p1��ޞ]�,8������'��B�v��g���"ѻa܇�����WM+�%t6�'8vXsg��t�{�u�ﵭ��wbH_��%	{�E�ֽc�����6|�2��)e�'��l����{��Y�_����&�?i�8P�y�����|%�F��0.l�;��w�F�h� �m��L?C4�Kp�qKWڣ���� ��6�z
�b�����pވ������Om{!]N����c��	�s|,�r�yĮ6JS��y�LO[����s��V"씧V�j\Y�����)�G�U�!��Q�=�k�9Fi_GkԱu^Ol9�v���m��P&z4�FЮ���gƐf�&��Җ��.���$����E� FJ��o�}9���T�o�1�Aa���{�.��� yP����eX�����R�v� x7Ř�5�M2���!+E76㛚���7�����;%��=o���FB�Q�-���E$�����y���^d-��YO!����qO<�{���5>1�P�竛����]��?k��V.��O����v���Z��@���+�wӚc�#�m�aJ
z��8	�y�k�j�_+��h�>�|s�|��$j�� ��츐<͕4���3���]'�i����� �=Nv�޼�V�£]�Bř��*a�^v����gR�eKo�Ӻ�(��nV��3�Zz�Y_+���˟gaʛAғ[*�O�����P�k��F���FI�lu��Ҫ���1+�UPV��Bm�y�z=]��<�
o�Q7Ƨ±�P5߫����(w�#faX?�]�zi�x�zv�y/P��������F��P���������k�wk2l�gJK���x�3Y�P���k'�?�sT��`��%��R�zJp��pGk�XjT�,�����V5�w�鈗$����`��Іk�)4Zd�k���A�M1�g�L~!����&��-���<�-&�EϘ�/�S*H�q�$��Go��Q���"yRxF�:��oV��il?�	��-�J��I�pti�M�k菶���$���{譨P�˯n.�PbY;�+.G���S�+FYI�(�/��7:�7z�=�#ށs*H+�� Ɇ�{x�'�.0Z���x��͔�Z�b<l��[3��P��(m�jPlK�-+��1o$w_�A���a�-A���"����ÈD��F��ŢP�]�����lъI	�7Bk^�����Y-����)���-|�AA���ஃa#�|�vj�rd\T_�r3�Y ^;d��-Ͻ��O�m�\,\��/
�UUY����pBi�ݓ��*G1/������ �܉Ѥ+%��a�,�Hs#��!���8�Ϥ�ϩ)/4_#d���X��J�N:9�?��t�pzUh$�	�����CV�b��5��*�'(G��v
ԧTZ]����yxC^
MX��A�ӓ��S�7K̟��%;�v�PA� ���"�+�#P�7n��SGO���Y��^`n�'3W�+�~��m��l;h�nC��y>=b��Q�g<I�l��b���������P�fuZ~�ĕU!��1l��g,���uq�Uɴʁ�w�>v^���:rKH�A��_�mTU��ӝ��z.-�:��r�񸈂tBv������:�}Bx�����~�jp��Ԍ�Ɍ��F~o]b�~|y��lx�ᬬ�V�-Z����}�2�v���Lv�`3]�2;4UK�Eu�:��q?��DM�a�ݘ<~\��%�>D��=ϡZ%��(�W�����I�7���(H7n\�{�u���䊥ta-�[�����ʽ[Ż�}4�P��������ʳ4�4�c�������ǭU^W`7Ɇh�W��Gxje�H��3�>�W׭��(ڡ�8��:�*�uYV U:_U�7^�s*HZ�녽q�(,p��9۷�kE�G�Z���ߛo�y>��/�S,Z�R�"����E��U�(� M"��C�]{�tnE���|,�o���ݯT�x��9$?���
7�^5�ά0�7K�7�P[KG#@k���:/��g���"G빒�/�:��]n�I8������y�婶�F�!����r�&�g���/|zk&����W$�b!R7@���J���g�9s��H�Zc��`y�="�#9ðV���х��}�C�	�o.����:�X�V�=嬧yh��ִ{ߪ*L�j���Z����n(j��O�t����1������@}n�x=N� -�0X��u�b�Y�S}����H����9׀���tפ?��N��-E3|#���X�PzV7���rd���ۋR����y=�}�x��dǝ�|�=6_{��P���~�E�������&�A)�Ż��n�'V�V��3н9��A�(FZCw�T�
u���s-�[S'�gĭl���f{����`O?���*J]�V�6�ݼP��| ��(Y����آ>kޭ�����]Qê����B��p%����!�Y+GŞ�7N��P�nܸ:P	q�%	dR0���^J�zk�茼��oS�L�h+��F���m�1�ٯ�XqK\���Q���W`3ݍi?���:�?��� ���r�����CaN����N32����6���ʍ�»OC#>D�� �du�<Դu��,o�k�Z=�Pw�����N�p!i���ƍ��b�'�`VIGLl|Ԕ��ȤT+]!uK(�-���B�)H�U ?�ee��b�9�lW@�DS�e̷RK����?��k�շC��Z�?�(4�&����iM�VT����d -1b�!G�w�p�V��O�Nޖ���ԡc��z�V�z��*oց:���ƽ�g��
Z/�<�X��=����q$H6�B~8\��$�ŗ� �m�%�be�����rD�L#_=�.���&Z_)�0L�E�7%�K呵�*�pe:��+'1�����Mo�7_����*[�Z5m�mVɷp�>g�!<ϡ���y|'�9eu��~��K��0�Xȋ1�¥�Ƕ,]i�]�⃞fi$�w�>b���r%����w�^�qaGPU��0�+oN<�X��c�����--I��<� �5ȿY��h����RT��X�w��ʻ5��S+H�p�aYk۞S�{L�x1 �M�'Fe�g~��#Q$)�Wrx�-#n��"�� Y6\p��i.�sO�����t�6+��-�z��tF�� ���M��r5����R��q1�Ad��ض*�g8�&�f���F�P�Hu*�A
k[r�A��j�0�.eh�!Z�4Z�n"��������դW©�`v.��},Ch��o�X��l�ڴ�@��	��=�$Q�%�N�db]��Y���H��O�ؕ���OH�l�fO����m��>���_G��3hr���ɛ@��҆>؁��[?컅�E�YP��.����w֤\���EI
���M�[����E�<OW%�y��<.C1�F�\Az=��Ŵq�	XKOZ譥��f\K��	h�1y>SP��kw.�<_c�κ����G;�ZbÅ��Eʗ��"H�Ў �b�b�Z����<Zw࿢/��0���H\�
5�瘱_��|��3`Ȑ+$��ַ�����/q��Z9�m��7��dj���3�UNӅvJ���u��+��������V��(l�7n� ��o	I��"����
][�����L�|cB�
%��c�B%�R��v����ۑ���ΌvK*����bk~:/.L�\x��u�>,c� ��a��y �/���[�ӂ}�VGW5k�X�H�^�S��fj�
������3���{��
�a��ݸ�U����Z���VX�sT&zʥJ�k�d��S#9�(���%Tp!ʯ�[����G�PbX��`]�%�f�:�Eق�%��*�E�/���`
��D_�V4m��V�ƄK�<f�@)�N�ÌX�#�M��C�Av��ש����h�s$�_���R����h�VI�U�$�%�O΃")�W9R�`�d(����"�Zu�V@a��Vֿ���<���Y|�]P{M�����o�S+HP�7_����Yo�XK�Rʁ��ǁ���ڇ�3Uoe��^���H�k�e�����G�cR;����(�,�m.«��V`>��5$W���Y�w�h$�ʄ����BN��x���+Ŭ��R_^�`mg��dGۄ�e��B1'��*���Ǹ��K��f�{jϐ�_넜�J�	��Q�a�o�=�[����量�ѣy�	h�ڃx��8���z�+ڹƔQ�:N�� A1`d�\0��.������2H�p���zڜQ|n��{�bɞ���
AQ��Ip��m¿ǩ�V缧���~F���2����0L�Y��c��e�d�NM���A��<1�� ��"�I��*�C��ʪ�%xy�3�u�v7�#�%I�J�j�<�<���`+Q���1y�'��$!?N�Y���ܬo.���/�r��U��-d�ʞ���_���CQ+�z��`
�eĪ���Y.�G��UUm�o���1�E 3��F,�D������)��@����0�� ]t�#�)��FXɣ%͗Ϯ������;�Q��4���7J'�,�`o�z3W6d>D,�,,�8��T�����@Y_�����h{����I��c�IW�4����|wA>����Q���?A�ReV�Jrzr�w�^��o���H����V�[s�ڢ_z{�ޢV���ґs�u��� z��8�iH*��Q���x�X0{H�H�¹���-gF�#s�-�]D�
��+�ǶR���ɧ�ʍ�A,#풤G'e=����K�V����֌��ʗ�U�oS)�t���Tt #B��qɓ�dn�a+�Ci��+hr���EW/gV ��].�6T~�%dg����V2w�fA��+Kz�@�����)�Z7��T%zE�ȨF���!�@o��B������R1���j�[��r,����ܒ�W<����Ȑ����y�Ċ5<���B
R��Zg��7����qc=<ml��N���[���O��� ������,�1p`�n���cuH҅+߹ָ1��26��9�a�ҭ�O��p���N��h�N�5�#H�r����J��t3]л�ݎ�V�e�.��9�$���1Xq����؊e����b���_�<��&��t�p�ۼ�?�6
9��M�\yU�}hC��+�������ފoں�XPiC�2<�e#��<&yW��֒ 0�c*/���8��㝌����{�fH���<�.����xԛe�+HQHۼ�f$���O�w7Ns)����w.h��!�U�c�-Д��|���y����qZ���G�F��ϕ�A�ޅԒkaz��C�Ө`��5�Pj/.-�Lg��J�}ɒa�������N�D����(}#,9a����J�hk-��I9b�]q�-I���v
�e�B�k�L��ߵ��4��N<K�g{��U�)�#�C�T2=��mkfב-�.̊���LJ�\^R*��Oi�;9�Z-�gn�ѝ3J�LUvx�(�[�k�l<����V�>G�Ȋ޿o&�*H����1����封�hrZ����x��O�?���͉>������!�d6&��0� Z%�j�dJzI�g�{)ˌet�� �{{Y*���0����U���U;4'��Q���I�bM�
SN�>��C�����<{�'%oA�޷JUfB��\��U�ԥ�FZL�� �g� ���>�^ϨKoA��(�S�b_�n!���B���g�!P&���?N���nVg��c�(�kR���`y!�#P����k�Ii�T�yl!ȒP$1��#�S>ir�Loa b�&�_�����:JY����g���~UبN�~�J� �dT�w��q=IX@鏴��K�2Yq!/2/�
�����/%��D���VT���x����� 	�^��� ^#��3��cK������[��YB.�O�4n�G�I���0JB~ڑ�N1�9Ņ"�,��:>v��r)����j̳�ݍ���̷�������n#�m��'�?�Y��>��]���EL�=��M�V��D��RB-˔�����x _OLIr�R�|'��4�ɼt�VqY�������]�֨���dE2�׷ �rI���8}�a�x��Q�'~�(5o��*մLO��J~'�1��G������4�"�8�D㉌b�����Ϗ�Ӳ*��S\����^���U;6�X�[YG�
��
� �d9R�5<-vyho!B��+p�y���q�1�N�K������vs
�X�)L���_�d�P����-�|�\&����H�s��]��gq.ǀ�׾­|�yJ�M{�ؑ���Ng����� )�୪$`O�� `��qQ_r��.����BZ���Bj��J'$A��)A�I-{T�]V�\�����=�[t���L�RT20l5���M1l2`��F?A�s�a�Z��"���Q�:61O�{�:�:��<��X����|p�����w�Bj��O����stnh�r�.�J������]���i� ɲ�T�Y�?{����g�ЮA�{���w�����onv�J�%�.�b	��{�O��($�3�Xz�[���}t�P*_?��+9	��]O$��鲠ZZ�~z�e&���Y\�3�O|�7�{�Gh�</+n�H*TġZ�{6�H���[��D��Q*��4����N\OA�s+��4�q��g�7� �[�i����f/���~��ě�g�w�9{Ac��M"��")&1>	ʉ��.�kꗢ�0��JB�����S ;�8y�g]ī?n�5��:%+d�Q�Y�Y۪�ҭ��J���J%I�������=��-:��~|��w_&G�eOK�֤⛔���9f��5�ۅ���/�՛����8��,�K�=FE�H�H�Lg[�����I�$mzQ�~�EQ�p��}ƶ�E�!��bm��t_����sq)p$�kE.1\��hZ{��<���2�����zp������[fs?[� �]`[y��{`q3��h'9^v�!�GE_��'v9��J��m�!E�F���������������7ަ]
��	��Q_��$ܒFed��3'����4�k��~@�9>�s�+p-�h���X��(�LF�y.�|�S�'��3�Q�A�X؆N�)�������?��a'j�����f�(|f+0�?Y�8%����D�	�aE��u�����ݸs'�S�VS��~�X@�Q>�����JQ�cu~B+L���Cxu���s�򷃿�r�����+J��|�&b�,j�;��$�,���ϣ��l�svӼ��?��ά�����\��y�</]�GJr�0�0N�?KhVh����g�6WF�^E��e%~�b�T�_�r?��?���~�)������0>旎�3���`�]:��(֜VN��I�?�8�ǯ�߸q�g�H1�i-49���v�LǍ9��]b�(N�F�#�K��<�P#���ۂ�[��:��B����ˊ��������/�/��q3�3_�)�B�E�H:�]��	2]��S]��嫽]~֍�"fM�A'y�,��ɔ��R�x����gSd���[�`��hh���=]�y(
������r�F r�Œ7yƔ��wedɌ��0�u���<��n��*�����:D���y	K�H[��1�	�E��'���<R�y<���t?�����{V�@��К����:?�抬��'Q���pzH���_7�?������p���\\A
�g�x��x��ODhҹ&9k�����р��œ�
�O���q�u?�sT���6�������{��E�R��s\5��0z�G����/�N};�?���������ߎ�5~���f%4�?v���z�0c�bb��$���0�3��s���&2,�v�w�E�(nU�gN!�F����T-�`����m���O7-����Z�|���!�h�<d�$@;��	�ԩ��-VE5P�㽗��\��$=7ʆ6�w��
��y�;;�u�#�NL ����d�u4
��uhK�e� �����q����b��=�"�����N[���Z��+619#NUJە@�qy�&A�L'�*SOJa�
O'��NP���P.o�Z$�Gi��߼��=�����mt!��!Y�$F�F 9fz4������ ��>�A���g5�4�BV����!+iY���G����8��-^�^�}X5��K:7�4�_�kD�ɲ���ǯ����o�}�r��.��k� �ԙ����!���*�`�q��+n��w�����?���ү*�|���H��w�m8�+E� 	ZԕNƥF�3�₿U6_o��`�m��gؖ�G{��|���x�j���v~& eBXv�,��.*�k��`"i��̦�N�uh�c�}{Uf��g�<�箱�D� "�p�F�Sf2<��Մҡ�����E�),�?Zb�;qK9�8�<� &�5����&�d�S�{�U5oΘR ?��aK���SͿA�]��LD3��0)%�e���:я���
l��!��QN'6YS�Oj�>]ۚE�	��
A5�8�{�}&I��3\��<�š�3�63�5Zj�N��(I�p���R�[o���u�	�0u��CJ׽�!��"e�w�%�(�L�� ��y�J�sV~���}`�JV���<�����!�1��>��2��807�$��~�29�GƋ�  �6K�i���9��"���(�il,�����\T�sQTբ+��$-�a5��TCwLN�щwpb�?��ܜ_��	���?��?����=.�9�_�����j$���+�0�h�h�kq������3�i9i�+E~�0�T��x.+��/[����?����~�?ހ��]l@�����ho옉�Fg/�/��|�!r:�"2���͑N�at�71_<��aH��.��\6����Eo�{�(���>7��6~��4��6�?��?O�o�%$	��Suέ�bW3��%.�ѣ���hh��:��Ń�X�nN�[���$[Y���&�%D�D*����x�i������B�\��}3�f[1�3�_ �����j�|�+��\���(�M�6�ؗ�&��TDH��ٖ^�А��]��/~�8��9{pC򽉶���Å,����~>�̕�hj=0�K���Ŕ�.}�W}6�R�g��l��:�8	V� @�a�TJ�Q�"���1k�U;"}&����w$�@w��R�y�f���Z�|�.�I	�m���R���ijI��͈�@���V�?$e)��:��˒�v��,V<
�s�b�
]^���n6�Q�qS�́���dB�PxX��ͱ��v&Ld��Ù<P�mI�u'/��znu���N�+���q�iC�B� %�A�kY�ڌ��\9�*.�F�Nawۏ*Hu�n�^��qD6��G�A�P��Y��W�u�y8��O+�!���Ο�ɑV���!V�D5��#%Ge�b~"n�b��� ƦT����`|yo��JPP�0�s�H�/�%%���K�}���k'|�v7�6����u��S�q^��F|v΋�4[���Z�=��#ч�3W��/��S:�		5�Vy]8p<��9"V���G�@��!bl*���%5:�^yP�Ȍ�gƍŞ��,��v���s��������&'"/T�tQ�LWq��2''ڌ^���C�?���d_�r�����+l�w�ٔ� d(��ˤ�F+�Ѱue������P���w������veĺ��f�ʤp���'�=��M0�>@��r`e:l��}���Z��@����t���`C�i�J��t���٦C���߱���ʚ;��x���ɻ�8�"�m�`��W�$ʾ���T-�ȅj>&*�8mBS��"���#��b+��3�!��Ĵ����@�D
�J�k�F��^>��E9R�	zF������,*�\�$�EzF�l:g�eM�nc�0ok�Q�#���E"�\8U	}�'=sT2.�e�l2�� (��~�U$�խZY��zY�TD9^�j6t��Xߙ4�u����6niP�M(�߫�(�d�&S�:L�����>��Ga�� ��(�Δ9ξ|N�]-RJ%�X.��T��,�+�+�Mz]9���Ԭ5H�����R&Ĳi<�u7���̀ݩ�����P%I	�ݰ+2�G"�3Et�i:7��{JA�8Ut�o�U,$��z�� ��6M� �c�!��HJ
_���Шt�t̂\�K}�>�7I���IY��-2�ƕ���ڜU�O�ʷ�w%!�Ŷ����,�hb��v���1ѹ�8��S�aX�ފ��_�Gւ2�ɐ\_cR���)\�h��[����^�Rc_���@浱��8��Ԑ�4�� 2�`f��4}��6�SA��C�������ڧ��畐��z��BH��.�,n�q�CoE+4Yߖ�K��mFJH�>P�J�\�:fZ�Syb�ǁ�	Iܴ#k!L��W�]=���|��
�JJ��9��;¿���l@*�4aI���`���$Wz�Q��\O�\c�mb>̜+��ߨ�V�δ.��\I�T�)ӭ!���hN�I9��å�P���&x�C��1�QX���K۬b}A��C`��X�]�ӛSxc8F�v�|k;��	s�*������s��p����XX��8qĲU�j����9�� ^?�����Ў>e~6�|�w�'���x�W�%A0�J����rL�q�`E�S�
*����4���5fv��S��b.�4��J�L
<������ϩ �?�na�t�pׇE�ݚ���&��!��.mGb����1��$l�q�W �\��-?��3�,[�%?[?�N,R�h,�ɉ��N�!:c��1�e�?/�&]�-�U��`T�hѫ��# �x��B�BQ�w��on������=ի�w��d���� �t����E۞��9֑��K-)�x���S�<��h��K;�Sp:�~�v�^�\R0���ч�ٺpR
E�1q��\!J�5�#��]��FJ� �W�H�ʆ��.��w%?�gG��$�f��L8�όC�i�)�lW���4�vC��o�d��rg�b�����|/<8���JN��"��s�uC����@}��&��^S\A�h���
MK���
"=1*�yQL%K(َ|j�+s�H��bI�z3�KU18��T�d�6���?�4��0!+���x?�A>�4�ͮ8V��F��DP/h�����`�@v��F����^�E�FJ.R��R��۔\%�ud0�zTm41hi7�K�%��䏦�Z���/����pҠKV+_�\·�<y���ºJ���L������]/,�n�)�]������ �?�E�a��׬��o�4��$���z�+mC�R�V�F�G���8�V0��d�ͱ��8�Gr�б6�3��.�t�n��$.�
-Y$"V���.nW����{�fd�n���S�`ShY��J.��y���9�gq�Z�+�r]Z�ɰ!��ƷM�qE+CtGO���m�,� ��Oך��3��:�@�Z�7�G��X���vV9�� �/���b�+=��ׇ�!E�e�l������x�[�Sȅ�S*H���@��?����vc=�-s�B�Y�}<R1jtn��_�����?U�I�n��M���	[�@1xI���4���]�2xP�e3ĕ=:CS���<Y+zo��DTF+?R ��*O��I�#)uP+�ç�����KEs�|�@a���9�c�?���ʷ��a�y�"Y/��d@�2F#��}���߭Q0(�8.�$�a��*�R���!�LJ��������%�|~L��wJ1rz7n��
�fl���4��������ݫ�E��5�Fk5W��\.��g)��-g+��5�Ry�	
������ ��#�mKn��ϔH��"�Y�����s��R�إ���VY�Ӂ�"��T;舯M͚jL�|��%{�J[�+��9�V�_��F-���nd��6���>��Dm�������*Fp&�ݤ$��{4��΢y#�m�y�6N��,Ad��X�p|��ͷ$O�_��Ha��}�o���]�f�ٛ)�33���H�������C�z��D������I���ȹ���p�(�SAٻaq�#������!�͍�ᙗ�	�%p+��;&M"���I)�I�bQ�,b�P�I�eq �˙�H�{_�B9�ɴE�RH7ӧ�#�DM*9L�q�b�/�%�,+WÎ�����=�Z"�W�l� &�t_��nԎڼ���i���g-}�w3}$��m9���P@�̨�� yCE�K�\L欀��n��g6����ݬ[�OR���'�z#EP��0g�qDn��5j
��ǎ�*-0�U�=F����\.�{��餠�R���i�o4�Q4�dg4�����ib���^_)�Nm�n+��ޘ�!y<T�d�H���8CU������pBi[�����Q�\��d5��$Mu%�2ה�Fd��^F.�g�H�B�,�9���E@[,��ǝ5,��ջf���1V�E�e�U�M��)
By%-m�L�󥞑�h5-�$FB�W��ۥF��z�~G�R}tN�Gc��k��Գ�L���+��^��j���0��B�Vc�){���>z�I�\����q#,�0GN��ډO��o�uǤ��P`*�C���b��|%ƍ�pB�|���A����ʞ�i�8�]/������0EX�<N���5ߌ��H
F�}���(g�͹V���m�y)pdOv�?SY���ӒoYw)�-vnL>!+���P��U�mg��^~&�۟�e镡O��k����hZ��z�6W�lIs[��v��3�ց5�-q�����h�F�/F�=�ؠ�9�E� �Q�*J����%�9��+Vl�_�[A* �+1qܸ,z������,�%:a\��a�b�g�5��l�"k��m�,�
0��/���p�"(�lV����v�[�kY5��V�u��թ��{�>�n)_a�h9���&��Z���c�������0;�z�,NH��=��blB.��&,C��af�iҙR�B}Fs:v���]���d�����֊q�1:v儊�Y�(�x�V}�d5VY����
���d+L-�jh	c#��{���݆;$NEA�-M�V����l�њÏą���e�1:�ߍV�4	$�� ������9��|le���b���e����ϻ�f~�p>7�iie��7���&�O{uE��D���c�`�:�x�ϲ���;�т��wK�=����K>�E/� -X���u�W�R��+Wy�*Wʻ�����F�m���J��ت�����zҙ�Z�g�cD�b�[��[�����4�v�ʒE!���kf���x�+k����l���mH��Pw����V�ԍY_]�Ϸ�4��V�r�XA�>ݻ�=��l��Mn| 
k?8��.B��=��Hb$d���du,�a�$�=k�-�d_9�N��@�2���;O��/�3���-a:�I�>���[�
+t�NbAR=��'�7��כ����9F{�n�J��R�9�к��I@C���|�y���Gô�d�Dg�,��%��>AX��ۨp�t��5��QY���6�U�[.�GH�-h��b{�r�q�%�	r:�K�JDfQrZy�'�es�4ɋ��5��ґ�|H��8�HC���R{ �v|>u*0���(}S���t�PAb�bk�1�h|x�d��wby�T�o���6�U������&�A��&Lkk�єh����#kh	&t/�w4��-�k��_��Ap�앥솙O�6�X�z�{�q��,�1��ؔ��s��<����쎂>?������eWJCR�ׂw��S���P�����>"�(�GJr|��v�^����������	CGI���e�<d%&4�`��|8�U�̰�?���B��� �6�@R�e��4HE��L������CW��ӥ�*H�p��ς�0vrH���ޟ�m�ƥ�6�a�ǻ���պl�n�ZI�:�˧���m�+]�[c�;}{����M">��G�9�=:$�K��U����ĝ���Z��-	��x�6�V���8���_~i��Ḯ����
)�����Q`��fx=��j��&��-�#a�w�h��L�DwF-�JR�٢�Sg�ϟr�֒��$�hL�%x�w��B�}na+�OO�Zs��+�zm�b�s���vlK3nt����[r$A����ڶe���m��=x1�SNg[
��'���빸����/G�!��`�-A�m����e�yl�[}jđ��^�NF���*J����]�E9�4����t�&�Wu�8~��$ w]<Iq���.�n?�%�b�?`<�ĞO0q�Y�Ù�iO�y�>>�O���j��c3epO�+�Z��<Ҩ�4^�rkߍ�DC.����{>BA�B"��������/���GM.��i��^��RĿ��~Oq��d�d�����R��bg��9%���h����	�#+��D"�#�������r4�V'�>!�����o���P"�^ڤ;w���y3쳷���z�8·���N%��g���%�+���zj��0�k����s��\PA���c�|�X��7��w�`"���  
՟�?��~���,�[޿�e�h�Ԃ	�@�(?Xy��V�:�*i��W0{@��(6�q�K8|�8�!*��'B����@dPٱ�JV5�����ߥ��pI��U�.#V�v�2�;��8a��J@+kY(����+b�(4,���K-�T�Dc�6��3VV�V��ޝ7^p_繎�
�d���8%�CV���;洔���O�O��-G$~��v1&Q�Z�`��(��l�ީ��w���mM��l��Q#����������z�%����^3���a�'���\N@�'R\@"F̮�)�/k*��[}W�=�^����C ����Ë�8�x�!�
�s�;���@%j���W��4��?0�#���	������h��N�,�wI>��x�Vb��A�����dop����p�5)2R�pNӠ�`[b�"�yA3�VA�A	��Ք�"����_���2-�2X���/��(}��k�@p=QNU1���*��΋pA���&�=^�OG-�F�7,��*���ëy�v^���ZI������%�􎬫�¾~䊱��+Jb)��.1�^���mg)*����C�k����Pf�p��+��;$�sk0��k6���Y�%-���Q���,��𛞳���jzcJ:W���R`��xIV���0�x9��$����f0�o�
#�}�u�;fm>���]6N�ZI��n��u�'0�7v��dv^��,�W3ƼR ,��bOa}��w4�R�^7����J��=��F�t��|��gc�J.1~��3��^iA��x�w9��]K ���̋o�]	�S�o2ec|��|~K�{e��_���ݸ1�*HzIu����p��Q+��Ls��p��/��Hnf/G%���G;F=?Y8Zذ���1q\��M���)$_c�����r��9Ц4_yp{s>��)#�l\���ڒ3v=�^f���|�T���Z��*qǸp����u)��ܓ�neTG��~�����؏���2��I�~Ox7�~�y����L���{m>� ?/6�y,W�X��'s�#
�>kzk�	��Ǘ���B�E:7T���or{J:�s��]ԥ��W��Æ:nT���%�v��ߍ#�	�"0fW�@�1�4��<�����2����1t���	ƈD�1����T�#��m[����fw�@�����
�������cxa�|I��[�6��p�z#�J����%,H�;�kd�/�+��}9����ڤ]�>�L�,��H�L�e^��%.*2�^��gF?�����F�h�����Wd|9Ϙ��SP�hX�l*rUU�%aX;�<[B�J%X��̕�M��t�������w�Gm$���B�te{����;��˩������¶8��e���ĕ���$Y�uXW��}���M��삇否�����#���j˙;���'�sx��q=�E_�l�����Y(�x�PA���W~NNwvB3	۬\ZX�rĭ�J��bm�{a��FS�V�J���"��.����V��C������ˍ��>,0ϑ$A�忕�� ^�g�� q� ��]���::sSP�lzI_Y�L�>OK���b��,�~���Z�����~\�̍1Z�<�l;s�Z��3����$i����� I/4n��.���H_���`l=�Mo��UJVk��8e?�%�HH�$�vK���w�]I-WAiJ��ԇ���vn�	�1�7t�	�����t���F�H�E+i��)��s��������t!�3T����-B=�d�La�ʣ��eD�R�`����&�:|E:��} ����(���vM�տ��ߪ��u��$$��=@�/��B���{��R-B����{JPo��ϱն��?W��#��J�4X�� ��'_m��e���˖�N� /Q����C�G�ǜ��:Z!�Y��Aнt�]#1��Y��O5�A�a��ۑ��G
<-�[[[S���1���z�g���[�����)�hcTȭ~�H5Z;�0ң�u�joN:M�96�ح��ޞ��J������^}B��U|sL{�����Yid�aZ�ەÍgᛶB�RA��$h���ߠ���O�6�la}S�F�:vg �
Kem�8����k����I>���zy"\�w�q�'B,UR�r���� ��գV�#�A���varIۄ>~V8��q7G������@���/ԑV�#�}�c�0�K�8��.��I��'|�!���|_5��Mug�V�hՁV�FYoR��!����f��[�Ӂ��X8[��=���k+�Q�C���So� ε��hH�on�/�pH&���bXCke�������r޽,y['�o,��xU�e	���]���v���$���x�b������+�~��_Lq�E�e�-]�Oܸ$nI�ې/������4�������P(1�
Yt��r=3%J��$��s��I������8�S��ژ�2�r��Zf����;e$�V�(�[+�ړg]`ȫ�4���BVp�2�u����2B�o*�)ɏ�9?�9=��n�2�W�i��ׯ�A��J[�'?2n,���ߤHV���hU�
�Y�kI�@F+���A�B6.��_�'(l^�ɩ e��slU"�D�~@PmbQ��b%8O�>(BV��F��i?��卌,���O�[AZ����EuvDέ�s �����B��Qk�Q�t�V�
OJ�	�:��i��W$��5k}p���L��S��.s��	5˽
�rdrg����/k�߽\g+>��S����h@r��ғ@� )(l6xߊ�JR�,^��G,f,w��LwV�*��%:��V��݊��H�7V��|�O��V$:�tn�[�;��b�I��V���;��'�[��	Eݼ����ʇ$���]F?]�c���@�����z�*�O��GE+�E~�9��wx�����V�?���E��0.����U4�|�Z�]���(�bd��[�]�娈1#���Ug�n�'⹊D��3�x�[�_�+�b4���z� b���a߄o��=&�qY����!��S��'��
R�e̖r�E�o#��`-�=�A��B�4�����~�,i�%�33`����pN`��������VF��o=����xXc"���R��Q"�L�Iy��)LgQx/�KL"��(x<Z�i{t�[A�q�����ނ�J�~$�o�$���`V�����-�4�xy����úv�M=g�Mq�cG+��s\5�%��V����H%mE�g��*��n<'T� ���Gv���Vy�d�y��Uz����2WHl�Ź��L�+T�1W�D����	)��,R��I�*��ap�oi5ˈJ��~�.���΃�+�Z&���=��.j@��A]J��� ��'��(�B�a �w�sPV�~�d�(j��A�A��B���xi`l7��JiE¢�=��n@q���F�\1{&L�\&�������Zy���:���dY(z��e����r8�_����3H_��'T��O��r�����\�;�x��0��:�[L
�������!���DZP܊X��P�P��/y��1�$��l�?U�R�&�L�(�W�8��p]�uQ���� �zQ���E���������h�6���|��~a��5+S��滍�c�L�[�-z)<��x�Td=��tE���Jې|w���w�1�^zP��2��|�o�n@�ϕUY�Tn�o�^7~�!f��_!L�K���V����5�6���M)�)��t�Wy�(����S^�&}Jә}�i�VO�����{�
�&��X�v-�q�7���+HA0�/]i�J� �<�8
��j\��ڻ(��5�𕃑���޼~�w�ߞP
gk �ݲ��Umhᚮ5��������u4[ :�j���2�/�5[��d�3�V`�?b�����N������Y�T#	*���Nl�K�d��]�<�5#&'�[�؎Cd�/���'�vM�O����1"�,`<{�[+�^����o��[��y���'��N��^B<���OI�9���,z�y%�~�籽��u�{�v�H^���%U>
�h��}��t��p}㥹�*u�[Iڃ�o��⚽}�7n\�0�����9�� �?ѩ��[7�Z{F�H:�������*ﾡ������?���e�b��ƍ�
R:���5@�R�~k��	ê脅�=�2<��k�8���aw�4��o�z�=q�<��~��XM��w����'�x7<�޻�Y��<%A�Y]�Y�Bw4����&K[�W�Rsڜ��g\����72�
����N"�`��h��Qh�1)Ga��؞9dn��sq)]~K|B3:�y_	vK�P�Ll��U��3��:��?�&�4����}������N����`(�������:�^J��{��a`M>3=�Sx�Q8����=4Ԝ���c�{1��	(�e�翹p@b�R ӓ��B�<�]ݙ��n����0nk�����W�x~e���ʢ򎶮�ն�$=-KE�{ )�|Ҥ�� �:Bs���,�Jτ���1����#�'���sa�;�4X���Q4���v٤��6B����|�Gt�I�s@��/���n|'�0�l-v���y�tлJf��U����h4V޽E�:��>筞�[�N��,�<�����WL�}(���3�T�����:�`��Ab�&7��n�|��*��.+��^=�Rǳ�e���F^C4�4���8�r��2橔U:��dD�uTG���b�8'�'g�O,W��ę��[A���F���G��-5��A��H��mV��A�h�;]N��>@���K���6R�����m�ɕ�B z[�X8�.]"^�lFkY�^'P�=ܓi �Su�����-1�
%�9}�4���6��7��Y7n<T����rږ�em{�7�SZJ��c���Qڅ���4����1����r�ga�x�F?B���/ވ������ؠ�3,C|�v�����R��(h���ls��C�E���i��a,7/"k��vI8��Cpk�ρҙ�/9�*H��&6Bf����iA�$(0�ĝy�]�=�%���x�1��z��~�粽.M��ֱ�t�M�vސ������ �)E}�d?��eh��r��@+k�wz��^m�:��GͬzN��j����h��n�Q�!�O�+���̔h��B��
^�h0�۽�<c�J[��>��o�
m�9��LO.��z�D+��)�#�+���O��{��\�j�}��^��F�Dt�㗼b���+E�!}�m���T�`�p-%=Oq ���M0�hL����7킒��Z�*Zdy���Q�r�m�S��Q,�aq�>R ̍�_�
�gc��={#8v:z�z��fi�44������k�X�V�ҪI�3�[�{��=ߍ�e�/�9�h~J��T�WI������k3�{п_�5��2و�+
?��eԸ2:T��N��km�)�2�nW*r[��$6�qC%���,=d�}�[���m���\})9W���)&��>�$y�����9���W���,���������CeR" o�ҵ<��.��9��'%@��� �]������(����jqbh��^��XL��{�8��F�ƿAj=���ܥ]�+���Goc��1��d�w჻��9���
��y��pri�W���-]#�Q�F��f�7T���E��S��.���2!H���-���7�����c(��',���x���P/w����V��:�7�(\�8� �(d>\Εtrwm�c"��7��}�VϖA�#��ι{�̐��[f��-*���n ֓^T.��o�-v.�w����1�غ�
��_0\O� YC��6}���W�4݃��Q��7tx��H,Zx϶�c�Iȑ�H/��d�u���i���: y/�h" �v㞨.~�V�e6Uj$0"�q�\�sfrن�2I7��|B�b����`.8��R}�q6�;�;�{A#އ�
����0�v��ُH�_Dm'�v�w4" \f0{���;o���r���"�jM�%LZ��Ѝ������Z#���Nb�:<Y:n��h�b���;Ff3��%��l�-VC�m��m�c�^��W���֡�pH��-mi?!��x[rNX[�Ҹ2o�TyN|�W�>��N� -�6�o���'Y*#A�����o�4��V"�L��u�Np	�"-�m��Y�W4�
?쎮V">F�މ�+X�U7�"|�͓-�>I�kn'��yaKbaD}w����-���ChMG遍/�����#4��$@�S�Q\
�d��;��)�(D>�K]ȧD�~���E�����t��p��J��"����6/=�Uڔ��VΦ���V�G]�?j2J���on	�c�s2��kM��]-_)H��t�a�憂T8o���0�|78�ѴC瑸����uN�����ڽ�3��� qA�����G���B��g��J���>p�ķvGf��2�9
�d���-i'aa6�i�-�}���)�.<׼����sa0��J-������i�9�����G2�Y.�&��9&����W�hP$b2�BS���ot���A�V��<��%}Պ�94P
����~Z[� 4��o�BĴҶ��E7�4G�g:���%�����E����.��[ȑ��B'�J���K:�4&&��,�Br�|�|���{��+����ļR��0-������y~yoyV�;�_��qL���'� �"�P�8�:[Hr���.^B�=�_�������e�L��WGs�f�wK�e��I.�ӷi����z7�n�$#$���>��Ω q|zܸa!�7�kn3@rg�s	�ɳ�2+�Yh�B���_���Jv[r�D���F�(��W�^�����*:�My�2�L�����Ch#�$�U�9}�Uz�k|�h �cb� Z.�g�R�p��G��EXA���?W�
�)���;��DX3������D�{�(4B>L��p��ք�N��[��*@��=(���FQ������)�o��<��ʆ�o�����ѹ�98 ˲�X��oLW���.@������ܥcXVD| �j;T(�0�,��S����ů��J�8��!��h.+�~�H�!>v��H8�!cHWY�7d߱�`*�JA�"ҍs�
R���*A� [���I��B��Oˈ�e�.	�Q�G�@
`�0��&�d´�#j`-���|r?�{�γ�@IT��K7�^���1��2���iiMjB�oy�^�R�Ū��xOi�cXZ^�0�ᎩO�3`L��-�ߐ��V����0��q�����@_�X����-ɕ)(�ǽ vvց���2P�Z�,2&���n��T������M��`1�C˄���/\�E�����$W���uC4��`K��}@L�C�)�Mw4��K$s9�W���-���A� ��I)��iU�]/>�sZ�����*�q�~�>�^�Ԥ}��sc��4o���
��F�����CE��[�Պ������z�-�"��$]hKE��
�F_���>F��gN䶛Qw���Z��.NR��&I�9g�2�<��+yrl�mIaB�����+�gR�byRI��}7n�� %󅶓B_ekĳ�{,���6�5%��I�Uګ��.�ª�':?��,B+��BC����@�I9�0Fu��P��CL��ñ��#MfRT�@��9y�G�z�P�,�!]%	�Tyrq9�mG�mP��\����tg�7X�y�虤^���Of��M���]j��D[[�ψV9'/�^9n�YP�e(1��b�?AQ��5o�V����+}x���e9n�"�.W�F,���7�'V���<9'3�c����q��5�V�>D�.,`J}���K�"5��!D�˘�
��q֙�R��$�\�����g�0I�<��BE{��r�ޣ]�Ɔ�9�.y��c�33wbN5�hL��Z��f���3p�uJ{G��c�d�uf�N�J[���~]A�a{���{<4(`��-�nq�>�)�9��=S�#o7BQ*S��o+�"Ѧz���,i ~T-R%�yFc��yp"��*�X�G�ۓ!c��{䋴dV$r�,U� �Lz���>O�y#�N��E���;\4 �O�J	����8v�Y�][�V����WK��so��7,�WArG�!������jtx�����k�èd�\�ʓ	�j�
6��0�VP�%\+�=���J^�Pt��V�K��S3pn`;�ȩ[���*��:WH[���� ��QxRJS;�����oOz��(�by���kZ"r�ʏ"�$���ʲ�l���Ӗ�HM���Ԯ�á�-b����'���>�W�qef0V�JzA
o�����.����b{�3G�xy[�:d%�ݸq	�XA��Gpk���IL�&ݸ�ո�ɚ	Zʾ�d��jE���ǠT�ه���3B�k76���_=fi���E޾�-͆Y����b�fEK�$!:�be����Z}��i�i)��>� ���9�Y������L-�\N�����޶��8��`ucB�n-��Uݟ�<08oX�5�u����ӵ�v}���&�zf����	H��+�u��+|^SP2��*}�hY��LE�
M�i�����H��|��o򱰒F�r�i'�_�ykN7΅+H��$&C5>�;��#y\ݖ�Hނ���Sn�D���d��l����]\X��[.�����( %�ar�M�͕��M�Bbc�>���X����E�N>�]��F�*$���DQ���z��d��v�BA.v~U1ی�M�$�'�,�&!k?���f�ȳ�7�F;�����uq�� �E�X5��Y?��t�5c��*n_hū|�4+I��1cQ�\� Τ	�k"�w1�̷lF�y)��b�v��h��$�
����E��4£�իX2��|hg^�F���9G ��L��k�n�x.� E�Kf��N�?�Iw�ֻC�K�q7N��.��kx
䳕V��6����f��z��&^���sOq0Swr8ĥ7&�[UN�w��2�p�2�!�� ha�.�\;Ԫ��8\k�	�}��0�O����e��o��P�]X8����D7�L����(�i��g�Rml�~)�� �@:�M�宑���)ޔR�}�Eݥ��Y�#C�%����Y�)�SLIr�tB�b�(�;��J"��J&�/ѹz�
�߱�#���|�:~�qM�q>*��iC���.��|��V���-ݸ�� J�����c��Z���P����'vda�X���{�r&m��&��)Z)5��I�]V����T�<�&u�����Z���ќgca0�I�$Eq�.cv��-עZ@n�>��km�kG�H�MT�g�D/��1�͓���>&�lWRZ���5K���E�9U8yN,�?>��6��?#"o�`��LCԊ�6�H3a��8���A�;&`ϳ*��|�k��8���q���
��%�R���h�;��^57ǥ]��d����V��n���ZAJ��Ƥ����Jh�Ra�ܓy��2�H�󭭝	b.�E�6��2\3�
Ȫ��!
|���f�h���3��p��Z[)��d�5Q�,%�$�0K,U�Б�{] C�ꂹZJ���(��Q5.��,xMx
�iQ����=5Ԧ�SSSDq���T��Ja����RC�2�	״U��������%�"`�I	��+m��䦔}�[���09�2�T$ږ3�+��J����S�u�$zCj�(�������������B��\I�o���Zf�"�l^^y�����5s�8�1�K�+Y�j�}�ȭ��C%?�)�����"O������"�^*g��r���9YΘ�D��Z:�D�IYS8Gƪ\w`��x��k�p��9p^i��l��ƍ��V���kD1�/���.���C���(�5�ʄ)
I�(L�F1Y��a�i�ZWe��H��)��G-�\��M�3��x�'��o�Qx)��kt3씦���x~[�b��з���4�ZE&|)���W�Y�)Ui,~�U�n���^�?����7��CZ?p")��| S��g����쬶k'T�a�M�Xș̜9�\�HK�ax�o��Rn����f����Q;}�t��pW)�2��{Ƣh�fRBl�q����:�·������߷�s��8�����b��'�d�qi�H�X�T4�VM<yKDVq|:)])�͎��ǉiJ��e�]"@r�*�S�I��*���	�
\Me�#քG
��O~�pE��"��y���K�>�n���)�v�z��l�-���v�q�E*��v��a0$m��rL6͏�X\z/+s�;�6�45O~���J���9Pwn+�XX��xh������mNws��c���Iw�y�qN��Y4$�ǁК)��MAHl%��C�f���D_�ɹ|�n���w�ۂ��9����F���(������V9�2V^���"Xɿ�mQH|Ә�a��v�_� (�I�4���U�5�T����%ˋ	�
#�"�2Ӎ+�
R�ݧC��y��%+�����ٵ�&�*s	��׉�{�d���^��.��Q�5d��◬��=�F���g��K�����P �y+_�i
+o��J��/:٨�=(v���0���i�
��aE8��"���))��5M.�<��H��YC����VK�q`X�|�,*�}O��(6_wT ��}���\�͠��K!P̋���80L��)��2���
��U�sP�L���f�E��okc�RS��^��?Fڤ��i]��mw�A�'�AÀTja���z�n�Q��9/��ü�7n�83.� ��q�9��:p����'�B��k�����W������w�����q����.��a���01y��5��{�T3ݺ^~�*��8��C1�ƾD��VE�B[���q�X�[\E�n�9��T�(If���꓈�Ng�:>�yQ~~�M�C�pg���:�UZ� �m�97�*�%�sn��*6�=���.}��5qY�c��Ӆ�(������I�����٠���e=�Q;>~�HOs�L����rT%���w��n�4��p��|�C�@�d�
+m��k���s���V֟h:Eq�+^��c�h�ͦ�c�Ft��ƍw�B
҂� �g����wkK��o+8�_y�z��~� ����H�������??1Aݳ���W۰,�xGy�j�C�c�j^e��渝����$rȂ��3��,m�<��$=��w�q�`˶�vp8�b��F"N~K؏o��AG���G���_
��Q��g{Xv��1B1���ʗ����hA�_�����JI�i{�/���[.\x����k`=5a��IC	���~���\�W�'R,����7�7}D��N�B=�t����.ɷ�2�v���j�Viw�rf��A�^�� �4���J-��L�am�&SK�[�}�W���&7�
�U���i��QUR�2���K9b�f�]���V��?��C��FZ�����96aD:��ւB��x�;����ܿ>��z|],���A��%F-*HT���>����-��[��Z�02k2�g���{e�qM����ꚪ�ݍ؈}����鮪����H� �dɒ}�e�ǶD�
�F�*t��g"?6<KQP��%h�]�Q�>������׿8x��lLSTn��\c��O�
{H�خ���2�`'ܯ2�O�~����"q���Iɜ����Ln�����~�yY����]Za����ˢ1Ĭ�h~;4���A{yһ�x��W��^�p�E��\4n���+ko��g*'|Nk�~��a���/fփnV-w��E^��Wp���%i�
E�P��B'�e������ǼZlǿ�����w���������_��:�N<<��˶Ay.��*퐩��}���
&���5���J_S
F:��l����m	+�û���<��G��/�{}vv������v���c��Y[���ۇ����E)�;%���o�8�5��ɾ�k�L��j�d*�IW��%W nh-���޴�)�J"%tv_�G��/���_���?����@�c|~����@��7��R3
�]j�L�MF�ե�v�1qM�k�&�*@I��QO�!?�6��-+G���J�w��3PS��B7B0P�]ͧІ�5H���+�����������o��0��\C:'5�0��[њ̴����
�����8�tOс0�W'�hw�zl�1��83� ��$����ڏˊ�w쏰¤iv'��v�����;3Fȑa ǀ�J�_��(�J��on�������~=4��ۑQ��/�y�Ȳ0���U3y�$_���,�</�8Fh>�*�uۚ#������(�ňZB������#,�ͼ:��%�=�٘�]��SVd����J��tc;٘Me��H�qI\�@����<�)��*��$��޳�
������>M,�T�p�b��7�ʽ��A~�Z�X�i���>N�Pc>�g�2V�i�&e�]Jٛ+HQ�PO<���M]O���2����3bH'0AW���jiU����*����"Ҡ����6{O��>`�۴������uE$[3��(����"�E������L�c+HC�V����\N�*�4�D���l�����p�T��_1~�b���:�i-ko�4i8�H������//��x�y���� x�H#��YC�H�A��f����~��]ߪ0�"����Q�d�d���`��� ���qe�^Q�f
��&�o���D�q�RBÈ�mb��76U	v�9��ʷ�
��t�x{��hI(+��+A�?���Xd�{	�ֽ4����)|�W�q�\�\���('�`����'�s��.{�ԇ���a����:�Y�Mk�z��*��c^#O����_i���� �+#{qp�`�XU2��a����m�/�/-IR��|֮�g��#��ⶲW��@�!����|ǀ���f�Fa{���I'/72�S[��2Ӳ�r�W���l��qn���2�yQ���x����W��O*׮�T {4o�A�?-׾����%�w��9��� ��%t��6������,�ǭ'ݸnI��y�_���슻�9x�hr��P�F��P�x�%{
  ��IDATzh�w3�+{��ʂ^����M�ޒ�T��]^v�в�8�:���U0�k�n5�IP����yD4�VvzR9F��5�m�k�R�\FG��H2�YU���葵�_q+18^�z[J��F[��>Q?^HT�V�)*�Q1+k���蠇�k��O�5�#m.�P�����󿌺�Kb������Fhy(]�����<�ֵ�\Ͼ�8�b+���;����l�}X��GVM�4���8!��*�B�0���8!��iq����7�m =��8�4��Ms�Ǩ2��-I���V���{�$,�������㵂c�%c*e�{��]� �R�[f��2�wnh u�|bXF��H,}��v�s�g+iM'�,�
�������H�a�Q��+*�KX"�;��2\}�<� T1\m���	�hMR@�a.� ��{r�en�Wa�B�Tjc;�Y��F�k%Ƣ��-z�hp�?[%��{b�{>�v��c��ؕ��Y�zd�b�#�9(�I���M@f�Z��V���������5)=�a>�L,��g���~@XU��g3R�?��~���e.�
�k�tA7�	�5�<T�߁�:��/����'�k]����d�B!x��(��/��KX
�C��zE'^�㿃a���� ��b~F}�ƨv����{�~~A��D����X<!8�-K��B}x6ym���\4E+<L�l�hg���6�D��>?�L�'�+����`����s���u�q95i�A_h����B�S=�
ߢA���,���qA���7��!�t�q')Z���z�������Ui�Z��DHlh�z�\�m(�bL���.ļ@�/4G�E;(�D��.�׈��d�VH��3�Bߦ>Ou8\(���V+#��u����I�U{ٺg����
��������Ƥ<
�~��ݸ�R\�@ډ[ݸq�}I�+�%���LA��Ջ��]���O�O�X�F��f!�F��9���O�){�g�&;�ވGx���4����� '����	~O ��o�ɑ��J��$hRX�B�1�v30��dō�F���؃��)��_�Ė�q|Dz���A<� �-�82t�ƣZ�2����an�d����'K{�>����\\�@�/�f���a!щe�Ha��չ��V��������'�e�d���/Ϫ���r��/`姍"�Mž9����E�i(��Ӧ�M���j���������g_�uz�-:A�ݴ@���½���әu��v�¡i��� -�hE&c`�Nz�t�����̀�&�t}I>�����o�+�
�ˍ��`h2nR�H@�e�U��<�#��n'ٰ�PM��=<	�vtZ �a���	�au7�5��o�����!|�iJ䍵�6�I�l�=6���.���V��@�eV�A�������\R��uE[/��P:�
	�)��~V]���S�����qc��� R\9�ɽ�,�Z�܎�AQ��:���Vc%�Y�M)�k�C	x�Y��q��(�(�Ehw��l5�A�Qe�8ڢ(E�J�b;E�,�.`�8K��}^l�Z��o=x��g�6����Sk[7#�	(�5N	���/	x�6ŧg���L��9
�RH��m�Yz�s
��y�A��Y�S;���<?z�����)W�z5����9�ET�P�M�Ѿ;*�[]�Wۮ�3"}�|=�4`�AL�V�ţx/QP�Q���W0N��l�H-����͈lé��.�
M�s8IH�~⍅���𭐯
'�Qd}R98_z�aع@�=5���
M��Vų�xx��e��A%�l/������k3�Y���[w��>x	귎�n��ӳ������W�I�e$>˕�g�ˊ����axg���LbV�%��{\`��DY:3�Dj��gB�*�*��e����иF5�B�2=�4Ñh��S^2^K���:x���Ҥ����=��>���^���i�a���'ŷb�P5vJ�ξ�������&E�+I�A��x����-_����'�c�I�&dV��qB�c��g}t\p��Ŕ��d�����=c��rM]����'���6��
?T��vta����/�����Z�Z����������1��i=��Ё��ȰI,��)�t��-G3���&U�f���	x,�����Q�2`�m��}��k9_!X�d�Py%�;zQ��/uFR�,e�z��u}���v�f��4��{����+��×�]�_IQ�u����MNX�W�S]� P����a�#��S<��T`f��y�WM]�槓9W����� l�����gR3E6付��Ώ���}�Jb^0�C���
��P/*�Y_������\
-��oX&��H��}Y~v_Ỻ&g׋�0'�gapY�Q�h���ӥ��	e�8��ٹ�3�P�8�`E��5�o�1�X�xr�)�Xx�/]��4�z��ܿq�=(֍���Tad�|�r��[��f�s+A(�����������tɧ[T����k"{9�Q�ھ���4*��$�!�+�Y����wp��3kxh,�ʎ�~��W��Bq�$#X�z:�M�\�c�}鲺�2}U���=����dD���\��8�:��)�ƍsp9Iz+N4OҞ�����Os�V�EA?���(�SoeK?�,�,A����ɻ��x�Ȇ]�볓��y�x�g{����_v3�ǂ1F�ZI�üe)O!?'���P3���"��)����J�5�H{��)�v�6�>?~\v�<�l���-���J��J���(���û���e��Tv得?�����.w��}L�M�C1M��;�s�S�o'��9O�6���_i�-�,�Z�MG|��ɾ�E�Ǿ��û��ˈ��kx?�3��0��Ű�PY�������Z�
��s����Y�q�&�P8M����ԻH;��.��0^�s�ڃ��\�b*6�S\k���[���I���SI� k����u����}�X�=���8�
���r��Oz�3��/�4�D��2m���՘�k�]s��*���^�Ǒ��R���k��1��������˄Կ@
sy�q����2�.�^p#d4��2o|�,�jE���&agvY���V��D}Z{k9�}�y�Ϻ���W���h�p�)��r�6��!6ΎA��X<^�	6*Fe����	yee��"_�v��������pM��L�r���$��f�?�K�j�R�TT!9M�
����9	�PW/��al�~��٢{L�FRMa�^����/+���9��ħ[}6Χ�	�B�c�P��y]C��G OA����"��yܩqP]GsdJ !Ӽb=��P��� ��`keiU��pO��x˂3Z�T��e:�b&H��r�(0��6b)m�ܫk�W�EW��6�%�-�9�!�>�F7�T?Yr��}��\�2�b�vω�s���,-�{��Zhk5�c�Hk3.�ɇGv�Q�w �3~��=�z	��R6�Y�����g=&˧���Z_ߺ�Ua��>\�4��ט�4>7.n$�W��
��D�_��]������%��am��Q/3=�$|���Of��������	G�V��%�Xʨ�ޗ
��@�٬����q?@�k:FC���9�|�TG�J����T�vv{�W��M��ʃ1O��A�/2�G !��g�TA}����i|�k����ѕ������-��}|�43�&0������(�ǅ$�ב-�Vʸ��F���Ђ�%�/K�t��ۅ����:� [��Y*Yu��_���ޗ)
e��^�P����X�n�o��K�b�OK�lU����c����s�WO糾�#�q�y����s��o�2�"E���-eM�2W���	g���_Q.��]1�Z�F�!�ɔ�)�H=
x�{����kP�4_���aC�F34�@'Ƕa����<,����r%�0c	ǸIln�Y��V�Z�:���Zq�h���G�ya�iJt�O�?�U
�)ww�z(�����Ҙ��ƍ��N�-�ѪLBqh���g�Ρ��J'���kI�c��?P.]���Օ��A�O�,��)�5��j��j�&\d�
��y��p��!������[۱[΄"��r)�ƍO�$�r�0U�nC�,�9��r�)��=^�d�G��ߥ�j��ۤ�޼�Z�K�C�i��}�2K������Ki�ګ���ڌ�U�����С���!{ܵz��mꚹg�C{Xb��SʰHk�׋޹�kX��<�c��Vǌ$�3�ڄ�
���/|�ĸQ���mh]��e���\�@"D!�����|ܸ�)��n�B���{�:���ӏ�o��	D�U�ɡ��*���[ǈ=����
���'�̞tғW�嵽鋯�{f< 2Z[CF�GL��#Ow��@�&҂�bT����H�����jRY�Yyv�&����wO���ۺ�g��ڥ�\@������(�����V��J����4K�d�[e��ګT���B�F��3���i�݀��F#׶��@�=T�*�U�F�8�O��[���	�<�H�c5��qm���2���v��5Q�� ~�|K���Z���q	Z�J=�P���70�VqVk^^��΄���E������p���H����eyG���<Of<��holG��l9S�XQ�3^���eyl��0�a/=����1���^|��ثu{�.П�^��J�H|zƢّ�[���p�|��[닽�ڳ���k�?�?>C���h�R�{�X���Pџ���ԚZ��sWF���n=��u��W��b'��\N���;�^(W9�e���B>|�o�K�B%�i�;���E�%�I�۩�fƳ����%;����P���b����ȩ��&q偺Y
�����Ьo�-q�%��&�U�K�E�7�<B��:Y��j�1cbn��ZnA�y#��3�T�֤y�_���{���8��k����^�7�5$�C�/|�qc Ch���|�s�cu���T�fC����,�V<T����v$�3b����}W�ṋ�V7����`�:�J.��o���#=����ws���:�T��ynEbĨ�Qt7DÔϏk�>L�4��7�n��A�m�����֛�[��C���( <O?5:D}����hZ��4^ï`����]㿣y��<�Y�Q��;�n$�o^�z\�@jP�M87>sϨzf��OE���Bz?��ؐ��?���"#�8���Z9��� ���]t*��j�5��
 �5Ɨ�i�ie�1^�ƍ�ϒ>�\��a�sv���:to+�u�_w��l��nh����K�����7~�&���?X��FͿj
�����Ϯ��������囖/���x�x��R%��^�9Tg����V y�SrW�=�4`K�������ո��nr�:��@ӌwn��Ƨ��hd�:W~�<���|�{s�i�� 1�6;X޽Oi�V���ӻ
S��=�1��O��K�=�����K������#��X��^���W�J/��_]7o��xU1��Fz�"������3�������U��1��iw{Y$��ȏ~G�-.~Z����~	G��(�*��ڍ��H��v�a ���$��@��h�X}�lݻ����O�?���A��`���=�p�k���s��G2<ɿ��H�jc�I�,��F�;�6�vb�_ǩr.YNs��:��#��wW�H7n�<��J��V����A��*`g/|o?w��F�Oƃ���.��a^e���K}:��P�KE��U7�A����{����;��<|��Tsd옿(��7�4.3�{��贶��P�JGO�'@���~���o��n��L�V >e5�Jh��ʤrU����ɺ�HH�v�>+#��I�J����WSJӑ����Ċ4;�"��0�I�{�����[�B:$n�~���Cf,G���L�_Y���[�;qų�[1}:���>��
�тN�Ox~C���OAO�~����KC�@~B�>~���y?��w��9�{{gxT?�&n� �nT����1��ǭ�У�~oT�s������t0���F���^�x9��U��NFd��l.�>!N{�a(�wV�'�{8fv}Bf���W�j�_f$�"�>ۗڻ��!x?I�ҍ7n��!�֞o����b�|�\-Y�̹qq.�~�`hύ�����qK���%àq�^~$F��WtZk����-�'�"z#��au/]=�����t�ƛ�+���(�7�@�f�Z����[+���e1��w1��4<J�{͕w��	��� n ic���>od A��Jrq��y��g��5��~�1<��G����=���VZ�\�1���α-mӨ�v������[��{�p��Ko�c�:���y}�U�?od �.Z��7n�0l9[�ƍO�=�7�/P=��ù3��$u�Ꞝ�LCO8x|�[}-��_������.`qs�)~�3�bҁ���<	j[úy`^W~z�Bu�����Q#(���*z���?ё����Iw�ڍ�(��o�d�
n���Mw� �8of �Q���27>���A�O�т��$?A��Q@ox��?��+�p�ƍ7�GH�ѐ>Ʋ�7z�*R�Qqot�q$�^�v�3^!���#��w��~���Z�E�����W�ϤU�SïX���%n���"q�
ݸ:��@,�2:^ӈe�q�(l�Ћ�E�_����
M��(��f\�~�𦙅�A�S▱�N-"o:h}��Ą2��8��qmb�qI�#�rA�}�@|�����W�Ɗ�2�@�&��ݸqqX(:�k �� ߳G�u*^I�ݯg�����	"���`�<��EQ��{��yx���C��i;�#�YKx�G7.��ᖵW5�0N�35[8ҡ7n\��Ҳ�~-�I,l�ΰ$��tzw���x�턿q��pI	�$ZL�Ms�T/�O�[��x[��jh����-h���>��{�j�r.����i���p��0*�9Q�q�Q��J>D���9P�;䔽/D!S�[*��4��
��<!,C��<鴝7߸q��@'�*�8�ߙ��0�H�ݛ������ݸ�s��h�c�P1�U�Z��)�Y�JJʇ3���R�sYX]�����T�u6��<Hr��%ъ�[p�i*�#1�r��!3�������|���b2CZ��7*��J����(�vڽ�&�pG�ƨAA��D�F��5o�,�,��I�ZQWM�v����3��ޮq�P��odx��8ѥ�I���y���n�_�(㈹rV�-
��>�k��4�#`�s���B�|B����Fh�C���|(M�Zr��t�]qj�*���%�?�>���Lַ����׻��-ÏԱF �G঩�1���}Vǀ�r�����=%�b�M?G�"7�J(pvop�ƍ���A0����N��7����=��ᨮ��ײ�F�=�O'�qe ��f"�^�&�|タi�������:����ٸ�����k�����ס䵽=�}�':���_�x��^�]�$ɣ���f����c0Jk֦�#V���׸��ն{�8�!��z_ܫd���{���!��!+A�m����U܋H�U�+H����B7���@������^M&]�7M�^Z{���1�0~���6ΠG�����ݸ���jw-\�@���i�{1n\;xzJ���!hJ���^	:=�~�6��n��x���Q�FԄ�^0�ȧ\�P�7.�'��.m A��ɧ��⭏��x��uB���^���A��7�R��:��Eƅ�g~a��[K��-d��K��z%t��x�%[�?ٙ�g�!�`��|�]I�D�g^F;����A�=&�k������c�^�ׯ5s/m ـ�{�?�O��uy�o�W�v����g*P���cUl�_�2|��d|/���M;��/-�Û)���^l�{�V6���&�1dO�.k^�5���j�z�ɹ���Ui����i�5
������m$���J_�.g -$2�2��a}��rI;ܚ�r�A��򅬟1-G�uC�ġ%��(�w�^�]Ưc��70j����۬��(p_�*�Iv��}PC��h
�
������r�[�R�2��1�N�D���q8nOѫ��ϋ���oNS����\�·��;M��������.W�၆�Sd6mT���β��[�^>�XAc�^Az�1�4�~3�:�f������	!$O'Hy�g^��UZ?d޾|cO�Í�p牪�p�#��Z}z�.A]�K-'6(�7k��h�6��ċ�3ԟ�
�~L�����^h�ݶ�k 
�-�Ag�.7�>V�gA�D(������jN��KR)[@�EX��:3�>G1�²�QY
���|utc6۞��Y��
��}�XMI�۲�r��@�,�|�]�so���BJ�	2m��	�/�}�λaa��Aߺb������qt��� \�⿠��<ы�#�(]y|,��gak���h|�00@��&�\��r�����Zy?/�c3@}~4+C|�-�W��h���u�YY�7�Q���25Z}\��'c��i]����I��#2�5��9W���(�ArAO�y�H�Hn[�5�>�(b�H�c���L1���p�_cpn��i��a�}!7v�V�þ�z`�5���Osa0]�KzI!�?	|� �D^�4�l?�QY柷��3���j��rRYv�-�:?��'��<˲l��v�S�@��ܳ��Vx�d���P��V�`����x��/taO�Z��{dt5P �+C�{c�����,S֥_L�,�����L��j!c��ӳՐ9�!u��ɽ��|�_����bpf�a��]�����gW��#��|F��� ���r]��w��~���)yH�U���Vz�{��X�<l���q>�4��g�.2�ۅe(�#l����;4�,cH�@�rꯣ�|�'�3�D�so����o=:D��������D��r���c�*jJ�y���4������Mɴ�m���d�s_uJ3�J��잵�u��~OZ�,`a�#��P؂�L��$�}�d�TƮ�4�޻�KW���qž���|�*.�t䘅\�&@#HC�p��ΓWJ��#"�tqI��;]�^�@���k����G<�L3���O'Y�+�~]��h-%Wt��s9��?��M��ǉ����p|�5�oJ�<e��D��w�y�͒�<2�a��09��_ ��B=�����v ���qW�6��Y�,<3״�w��Z�N�YYQ�|HC�]�_Y/A�+Y��2�f^�����p�3�Y�(9�U]X���YN#�b\���S-ٴc�,�WG�V��=ɕ�X@�0W��@�˕|����1b>8B>f�)�L�<_�SAN$j��k�Q������e|v����S˽�xd���̯7��\
c#���}K|y��Rgy��<O��P(�D�z9I��M����B��Q�.�E�<�ɲeD�a*���j�5�	̩�I�=}=��|�e����#���5<�Y�C�������H�)hs�2������ͤi#C�K�0��d�`�����H�=q�r�����?yt.n t��?���q9��a������Լ;�g���!�#�����0������5��骯=-k��H("�����֔�n�+i��O�c���!թ+4g�j��_�)��Z�=k��+����F/4T�=y�e�Vgo��7z��)s㽸� �,K��#�8��������s��}�<�	����9�o׵�5v
��t���CMF��x��ޗg^��h*�bF�r�3qۘ���&h�E�f�����]U���������o�7�Fg�嵤7%��䢽�DN{��x݅1��*�*�*ș�E rDE��;�)^&�s���UC�)_%�[r�F���� n��ǀ�_��C���sYE�fc_i�*���I���Ѵ7�r>���	4R��o�+��N$-�XB���ʛ�E�tp�p�����ֆ��IcE�7k�܃�������CW����8���>��7у��l��P�@����w^�K��ۺz�V���U�N9�Wd�yOe�4�2�c��-��aZc���ATQ"���ۀ<G~/}��/�KI�X��+3h��98[�^�@�zR#J,[(�JY��Ν*���N8%���F!���Q�a���'_O��A����������� 곖������[ُ�*u��4fh �j���8�NRHj��k��̭щ�-l�Y��k� 4,$ɣ���;W�E`S�gl==��9��(����*)w=6Z��X��@�r�.�;٘�&7AS��0l�t���=�,�U�|Eє��5P�m�N�{�Ko�8f}\�[m-�e�4���$�]�~m�`�GM��~v��7���	W��e��(��
��~�ز�4]��[@lҒ��?�2]Z�����ಊ��+M�ˣ��A�۟��Z��5��K~�7@�D��tl=��3"�Jdz��>w22�r�/{%Q��O*��LCi�O�R��U�G�l�Lbsɑt&.i i�n�-�1房��s��Q�GBz�9#d��w�Jސ��[�bJ*� |�	plBz��]��H��˅teov���f
/_�ѹ-��V�����Ԣ�B��ި�rw�ӣ��++S��9�f�7��Td���~ �LI+2�ν�����!9�-w�n4T/�!scW�)न&)7��g�JI�E��+E�������v6=�i��d�s�0�i<�,�åJ'�ѷ�l����:�t�d5�M���*L�ʰ垠����_���p��
�終��<G.�%�͟��=;�΁A�32U窔���ʃ}�Ɯ��`�=2�Q�
�(_UR�E��ŀ,������ɂWE��|?�4�p#s����k�O���Gܧu��g>�y����s��<`�9
5���Zg���=��������M� �׭+�E��k����k�LOi��d �:�)Z.1�$m<k�=�)Yn�)��"RZSI���|�N�V�}�w~`��ʣo� E��а��Ji3A��ָ"]C�D��C�m:�b��$?n\�&0vr�e��%��a)�$���<;�<R�+��Y�B�;�"�s���+I���-_��W���w���0�����\�+!3�&=m+�`11��#̣�;rK 5����g���I1��O)���H��P����Ώq>Y��ݥ��
Hm��h/�$Nf���Ӿ6nd�i3]�@�j ����qM@E10`j�Qѵś+�G��M��9�C�R�\�X�M���z���e�lcjG�N��+��ޥ&�t��<�ln�Z�Ԟm��B�B�)�M���R�h�gnЄAj¸`���S��=Te�M ��4�yZk��1�l���*Χ��I�u���Jwӡ����r;�'+�ymG@��v��2���!��HC��p{�w�F�:��8���'V��N�Z�dE�Tk��^V�*S�R����J��fG���L���*���2�i����\e��Q@)� ��d1�T��c9m�a>�����>u&~�A>:m�q���y�riX��R�R��NaY�;y:g��9Z���FJ��Qà�����B���[Ɇ���$qR�$-�T��imh=�������
�q�w��t���\|�ÕT�i�Ѳs�*@�-� �#�A�=���r�O�;4�f��ȣڃ�6��5�b��� �KGy7�/u���l�/'�Z�m)�� }��$=�����-)��&"�:ut~0g�j,<�� �jo����ɿJF�Cv0�&"����S.y���ɞ�c�2�c�zGz�̛�r���W��$��5�MC/�ٝf�;�3��)�e�ㇺ~!L�����dϕ�u��Vd��K��{�� @q����C��y��A����g�`�c�7\�d�{��V0��W�$�|����R`c������l1�M�۸���
~�����2�f�x���#imL�����G���6�=�j�Ȟ�!�2J"Ů�r�z'�6�B8ձ數�6�u�9����R�8vc���j��L'+HL@�$��� �Q꬛��z5��?=���J��F�8kz{}j�*�'To�\=O�^�@��$��*˛�'�(�o�
�V�������2�cUtk�RI9�����]�H�TcPX�F�m�̘{c�\E���PS�7װ2U<�*�^]½�d��w�gY�9���g̴��R�0�|�G*�E�?[sЮ����_�t�D���7�h��G�s�>��((���Ʊ�����Jf^W�B�J))��	��`�����hLp��֣o�|�y#���x����g #��/���9��g*{����22g��͋��^������~����c������t4Q�XM�I&��� �|o�D&��\A>i���z������n%��S�	�ᶟ%�£�'u�9�&�(�\$�0m���λ���
�~z#1>�?��7nx���>��O� ��V��>�B8ӦuY�� �N�J�f� �Hֺ��6l�� �+
aH)f߫@��9!#���e���)<HðΓ�)]���4U��5��3{a��HG����� 0��NQFښW�q:=,�^�K���(���{����1y��B����EV!�O�a��K�&���{��Z	��S}�o�S`���]�GG ��g|3Փ�i�c�W���:�7�d�ה���a�HH_3m!�&Oy��5Y�k~��/�^n�˩����ur�f�|V!�y�'�����y6,��gބi��ʛ=W���YBP�61YM՛�}=��p����������<m�%PSC=��'�BB<�m/��ů��D�4���I��ZҿS�=��r�$/$�������LN�,���$4ͺ��^�޲^X'E�����e�OǔS��qFR�Qx.��[&��W�������G�x=����j�@�D=�7 ��j��h魏�o�SG�m��_��$BvK��[e��x�P:�s�w$��QР�wA��I�]��)�:�� ����Fo�SZ���FB�oZU �pWzf�Z��k�Iz�s�͋{��+�����i�@Mu��;l�lm��QG�� Q��@!]=?�8	�u�T�hT����Ns�,t.��_i?�w�$:Z�&'�;�X^�9={�`�	JAV�c����<�����)�{�Z�q�g8�ю>-FK�P2<!�S��;Q�_Γd":�J9B�.W�o6�U�qMɹua��;�Sw��z�q��|�� 2b��Tʒ4�_���t�H��~����A��j��g8U���-ۥ���Fkj��P������{�w���js9�rE��l��M���X�����S�FM��P�����M��J�t4t�/^�
> �F�<f����c9��/�6�q�
��/ԅf�<�B:����ւ,X��1e��r�櫓t0rlb���W�R��:�0@����q�63dn&���Mt���Z:��$�*d�3��͠�x��N����Y,�:��7�nYb�y�H|�����|�k+t����y����	�9���M=q�%F��\�XU�rUͭ�,��ٔGT��R(��~J����٦S�?�����Ql�|��QϣY��cZ-�I�@"l�5ѻ�/"�_)������J!]��f������PY��0�Wz�AI_��M�)'��W$���yv���� 7J�B�bF��9|'�I次n���zh��=��mU�F����t{��Y�]�<��1�&��^��u==���A��UaA�ޫ5��)����lY����-���7�����H+�}>�6D�:�%�B���;)tj]��2��g�������kxBPX:N�J�	}S36I)	ŕ�~Z�v����c�p��ʍ$�Jn$e�5�<�y�4��gy%�@t����}oAkc)�
-��h�<%ANv��L��!-5B,�./�����x��HnU}`~-�zfLD2����#O�tl ��`��i��g�'Q��7�5������ˆ}韙�m&Z�Α�͊�H�U��@���Ov�k�E�������������\�TG�Л�@��;�|�3��B+�j�r�̪�خ�5�3V���_A�F'�l�Me_T��ɨ���1�>���^N��`�cdDz����[R�k܃��u��A��ȡ|���h��0Vj�pm� �Ģ����4���)���uTd��dr:_�5�d?�S=�=�օ�/j -��ۭ�S!m�w�Y� 1>>*�b$�b��	'w��J�sB�(Ns7������T�B�<4�7� ��z�åK'��S���^Z�gR<�%ƍ�^�@�B�ϵ�Ig�#�ݐb�SEi��@F��	�1ۿ�,E0�N����ی9�k��Svy�B=��Iȣ� 6uQ��P�o\a�&kW���g q��a��o0�����0!w�+�s��k�9x�)t�[^f�Ҋ����PȧȥĐc��:���e��>M�U-��̘��F����9�T4ρ9�X-ټf�D����`�c�(x�ot�:��ķ׎�*��m��<�"Fe��� yp�h��1��AAz7�w<9�$^�#m.M\V��$�)���Y�/'>��hd*NsxĶ*K<�"F#w�V���� �)􈨫͎����P��/��)�5�[͜����IB/����I���S���8��#?���*5��E���ww0kSL8��5z�4}������	%b��Ѳ'Cy��0��T�vſP��t
\&���;�M����U�S̥�rR
ۼ�d(�Te$�}ƪk�q��L�i�M�˵�;���z�P�.���~_l,9�.���q;�dx&�+��d�ؽZ�1��[���/�����V��VbZ7킟IأQ�~L�2�j��s�iG�6���2�a2P��a��T�� �v��Nߡ߿��N"IL�٪�a��
�dbr�Q�h�].*L��:�i-�S�cgM�K�?�I�sH^9���>;\S�<�+�c/4��	~�A!��{���N�3���"��/g�,��}{�R�`�<̓.Gʻ�4f��~�b��A��%?�.�D�킌��y����6R|$;6�;�P�+A�ҟf<(R��yPv�?|��^U��g�,[��-�ۨ��ƨDm%��CIǛ̫uj5�Sb��s����.9���vZ���'u���^s�q��r�z����q�t�����	N�(���Q���������%1'(Ģ+�ݨ�9���������Tb(�s���4i�����N�ʒ	�a������P��U�*���e@n�y[���'lj[����i�֕����_X�X@����N4N�a(i'�.!	(^W��b6�=������(I�R�����?�]W@KJVm �N��N�^�P��{u�0F�h��[���S���ј^YE:����Q�Nl�<ܫqUh�5��]u��jO.B�,����|,�6��ceC�J�\��4�<[Z��3�EN�Z���#���L��k��j2�~#)�)#B�W+��Y�R֜� �~��bU.��AP�1�����H�q��1�9W6=q�Y"�R��J遥��#��̛���B1tJQr����5䳆?�'&����inRąs� _V�4b��&>)�q��>S�;G�\�NM�2P׃Xϕ�|QP�҇��	>�V3���J�V�qk���
��n�ye����^a�
�����������'����Z�F��i9k��̙-:F#v���E���#�����ܜ\zO�c��y Y�ݣ���gh.5�Q$���j�̗�s��ѫ�q����a,iR8��9O��b��$˘#�[��L����7�M�o���&� �^��!+���D{UV�<�J?\ ӧ�"s^�G+G��w
+��S�%ˍ�5>��hj��jJy`x��=]\�g�zޭȅ���~�AC�^=t�;@���V�t�_X)�o�kzZ��;�
�|$�����ވȣ[�w=�&YV��*�^�6ߏ9�����`�c�Њ�,�r|��#�3��I�\��}�� �	l���h(򽮓��}�0�<j��q�����#G�j�h:����7T�2Z��:���GT o\��PK{%����Jc��e�r	���"NN��h$"/����*�+������E$�����J5W��e�K�}N��,���V��CK�<��,�l�0�%�Z:s��#�� ��uX{V�Z2����I]�	#L=���e���D�a��z?�*_��8��.	���BgL�I͹��=��W��x�za��*V�Z�*��)&�:����;��1tH��]���Ow�g -���G ?���0�!i��;;�~��.��b /��Y�l)��,��˯`�bf6�!�V_
��
\\y�YDᾒl��Ə�	&���Er�����c��|D����s��u��1��-O���:n��})�ӮҾ�� G��S��_��b��1�+A��1� >��/d/J��d���)��g
S��Ջ�J,�꫐Dc�������r�`BP���]�����}��/������.��z�c�I0��F�I�������_�~���t�Ac�P�)�0�r���D��� ^fT�p}��PWGs���A���nC�T���<�hLy�9�)�
���+�M��W�>8z2]�ь�>�2�W���JJ9�B���*���3z���O������_n�\��^�����aI'����2*�G�� i2Y}N��e���N���z�G�Q�����U�Y[���'y�@�7��Ͽ:�����m͓k��2��;}'�K�W���C���������_�r�P���^˝S��&5u��4MQ~��.�"k�4˕w�Β	3�������J�|� �p�bz��c��
�<R���j����Jׂ���{���Y����=���?��C�<�����cbq��ĝ�F~�����fGT�0�䍴	��I�U�%k��1�O�;L����;�LR����4�EeC�d������>�F,^��ܯ�1��cl����_��W6���r�N����������BbUج��b��C�嵏�-�G�~��O7���v���wP�"�X=�������<p���SZA�V��;�Y�F�Vz�o�9�%�J���u^�>/��^�j~��߿����_���nD
e^����!���������%O��֬E���v�(th�Ɗ-���G_���@z�[���)�B�`3*��B�Vn_g%&^�D[�$o|k���_�	{֒W9�{@?Y8=�~UP���YxكoM�RҗP�kr��E�)�K|B�y��6Ґ�ܴ1����,˹�`�/����v_��/����Y��}�r$a��W#`������6���>���u��,�Pv�L�����/~�7CtP�U�E����͋s���~{��o���q��Y��.�3E�M�YGb�X�g�q�3A����1EVDy�1���X;��!/>6�4/M�1��Ҡ���U�v�I`�u ��ܽ���<;�Ut9���)f�!#z�+�=���F�E��e>-2�۝��H���1��q�rnUz�ئ�6Z2u)�>�X 's)�|凴|�dٞ̽<�d��&������x�O�^$��$o� ��#KB��@���.�GzKA0�V�V0�Ǐ_���{��,
����=-a
�G��P[/zG�G��O���������J�C�֭�2��_n��o�cuZ�֜h'�ڡ_[�"�Jك�^�� G����,�虫�8X_H4.�RU��W��D
q)������2���|=f���pA�$����_2K�d�5M1=���S�Fk}E	��O�MJ=���m��/�t��TW�q�}�ûZ�̛��8�G�S8MOY�&����v��S�q�w�  Փ>!(�A�O+/[V5�����śk��O�O��E!����ke�L$]����K�37ot�?)��͝�oH)�b1*ʾ_V)��NO|0�0������$fH&;����Ru�^)�#�2 _���,���C-�*��.��43u�
��"#��C��b�-���]�+�d���Z���;IZ�N|�u��<�GZ������鈈:фH�ZơC���p�.���� ��&�	�m\����䊩��b��N�W�%�t�W��"�fA3~�	���FJeP�S��Զ����yW��T,�c���l�g�GW4�|���c+'�F�(�D�e�y:����8�yH1Q��|��L@)��T-�E#�	����K� z�ٲ��E9.!2��y��?ۺ�w�j�k��w�j�p��8Ǖw�ⱟ�˚����u}Ʊ^�~��W�M�k٘�By�Ea�.[�������in])��@	�F�vh5е\�FZ��Nd���Ô< ?����/��H�l��Z����n�/��k~�g�닾��Q���A]���ml(6K%ZJ� �{��1@i�y��j��G{�����SZU){��^g��Z�vo�k��iXF��Oti� �˺_r
�u��b�)�L^�
.{���G��~��K�<O��*iw�����(�ӳ!�^sV*L^�e�8+W�xr_�j���g~=ha]-Y�q��U:t�+��E�@�i�d�\�U�b�a�2�)U6�����b������+�i.�a�S��5����/�Q�\��ҹ����Z��q.���4�:9�X&�S�E�/��Q=y:��2������0�e?������*/�'�������R����Ǽ6�7���,�"m��@�X�&�^�r�S�k�u}?}z1~ēWzhșq=ɹV'�Ni*�ٿ#�خ <O.B�= {�q��k��S��>&�+��
L�P0�������^!��b�:5C}�`T@�>���XH �������,���*���<�G^�Cz2����ړ�>���T4V����Jn��T��U�/}�(�?�@��Ӟ,	�l"R��68��T%JH+��x�d�W_��>�$�\�ƍN��z���!F�Xi~0Ê	���y�*�S4x�y��$�l����2�����/&��[Ɍ�L�`K���'?���֟�~��"�軖5�C�M���J��9�q-�EVH�%��?�v֐�i����¢�T}R�0T[5��d�ύ�5c����b��?
��ZL^\�S'�o�e��5�eS����}��l�.J�	irD6R�z.h ��&�OroW�t�R�z���(I�(�2T�`�M�8�o.������q�Ǘ��R�+Xz���!���@��@ֈ�J�VƖ�$�xHd���:�]����9�B���"�pHt�ѵ�E���)UQ�	;f+A�wă
+U�>w0��� '��֥'qs7�&�R<��9ǂ�K�ə��UV�J��cb�-
h��Eۖ�H�p�sq����&M������/�S`WǸQI�e��=�p'O�\ç�A�/��(�bJ!������������(>DF6���!��+LU�ʦ.	�K��.�LL6H�v}�h�j=9`e�:f����C&|���O��G��\�GV�����{�4�\�3%�B����N��q�^����̾�d�ֆ���-<yK^�v='�%b0n3[e��j@�.1}������@QJ���d�r�8�^P{mX�&��˷g�GT�:Ivi�zR"1Fz�G�HP�GO*"����#�)́��:D�E��!�-��T�K|@��H�vx�d��O"3V�{0���"��MgBw/Y�uj	E��V~
��H���n`(�SH��l��Po�P�}j��� �}:�I��!wD��V:������_�0Scm<�xv���:���CKs!
��}5��L}C9@�.�KH�Xjʩ����%ﳩj�#��h d�&��5]i��±�S���~Ń;�(d����ϓ����AD�.�xzZ�e9l�u�|��7y���{_����.:x}�
���ZZ�*b�����9{v]���� �WG���hNx����8���Cݐ�=g*S4z���$H�S� *��
��I��r�P���!}D_�\�Y��8V#1�W8�>�R\�sf;I>prEE�
]���m\�j>��,ҕ�6BZI��І5>�sc�)���3'���$f�S���Ǯ�i�-'~L.�����8F�������]x������C��R@!K ���b�ʳ�����j?�`F��~�}��/%E㡖01�V.���`��!}|�L�^WX��aW��,5��-nP#+"�tP������Y�58Q��V��ƱN�s�����p���j>�'�F��;�e�(>6�G��X����[�t�^]��W�G����S->z�����L��6��t�'��H�0:cM�1<y
�yj��[y���iݾ�Qa��H3$	��
��5d Dۮf$q����U�OV�9��=^bu]��}�v0�Dt��v�B��\H[R3�?�T$%$���Nau�C���H��G�f��t\�J>�ϕ�k��; c"����'vP��Z�@~'��㊈!=)���Ç�_���^9Jt�_�Ly��P�'�d�)�%�θ=&�П�{h�X'�{����+t Ox@��J@����u[�ؘ�2��U��1��Y���J�(4.�\�Q�ʨ'LNu��/�U�H���%����r���ҴO��Ϝ��4���"d�1��JL6i �(叝��&�p���<��En���Mz��)���t����p��ǈb��Zv(��@�<	D�c�N�n^z���K�/��9���T[�y�� ���;"��ʞƜ�(����9�F"���@<��b�,Vj�3ՎAg�0
���,��8���ّ���6�d(k��[��O���T�oOBAg-W	x�5-�������P�xiN��4X�5~j{���S� �����Uf���ң�#�@>��>�_q�Dr�$"�/��:Q:�L=�H�_�N5�/^
�k����.'��';-����C�%pfZP$�e���#o�4R�U2��4��Qi�>ͷ�ʶn\N3��x���e?:�����ך�l[��b���JF��x��l\�@B�ww�Oqɤ#����7T_&c�]��f��d��ZD�q���4z)�t�=�3�!�}j��cD	�W�2(�bC�o�R:A;"��i���r��oQ�<�lԕ �,Y�z�u�	�:�g�dn%#��_�3��M�s�eS��i��˥zK/{4�2	(Y��K�ϓ�c��9=�`��K�|Ճ�zlA�i��js"�va����Aq�����x�ʷ��P����g�R���3�Rv�����PN҇�T�r,7(�y��v��'F������s��tI��Ͼ3����V=�t�#o�L�6�	�W�x(.d0NT@R?��{ҖK�����+��H�Y2�y+r�0^/Г|�T�o�V�트� H�
,�M���g+��y}2)U)o�YӸ*p��������P���F��W@u��;�!H��̜Ee�t_���rt�|'�XFP�>&T͛���n(���z�\)cn����AϿt�c,U�1p�"��[<�6�F)N��RK���s���S����Bj�����36��v��r&�y���no�.Wf�+��y����\k�?E���0�7���%$�_)��"W�T|�����19p��6䡰L�tW��U��EVwf�i��"Y���%��^.j{)���jISi�Bk�K�s��4��C��� ���G҉~�ƄJ�{��r?��N�hO�]rB��Ž�;�g�	4�&���mfɋ���C���]T�}%�O���R_�;�j��t]���N��|�p�4J���ʻ����u���b���~��}�n���S߲�����yg9�[��^T��u��,��gI����g�4�t,��hX���ʐʅ�;�yv�����s�z��i ����?	Q�I�]��J���8����yn
�}�Ʒʒ:ޗ�^���#)�
��7{��1X��@E@*�i����O>�T�8Љ�,���������<��������A�6�yՋ�����V#Y���Kv޺�Od����J��"����P^L��!�eL�X�Τ�sƹ�+�Cj g�� o��(;mC�1�?4���s�?{�C(|w���J 8�ձFt�/��n*�m�"o�Mx{�+�U�׋p=�d}���H��"!�z����jp�j���P8�b`}Q �Wz�w�EX�����:���͹��~��+��@���G��ˮ�6�O�u����>ݔPT��&A��x�z�t�`�=O�Pӱ�VA����
 �n�����g�މ0혲��4�A=Γ�eDH�SWCY>�6��Sz�w�n2Y̗�8L�b���'��VHKJ�䑺�,����'�br���rj��{\��	�t��u�s�Е�P���SF���S�,/f(O��i#ǔ9�M�!{W��bk�bx��չ�s9i�)�o��N�,�O%���W�J��}��G
ŤX���/�X3]^�$��i����w9���)kуm�d~��9y�AR]
;/�{�h�ԚU"YnFY����S��w�*T�Ӟ��������Q��Z��O�>FST��O���r�����ط�c��G?�B݆��p�7���4�|��,��g����tb�i%
t(����3n&V$~\������!�������4T��^0����p�G}�&i�Ľb�1J��th��([c�#��Y؁�R9�C��M.�d�}3k�̴6�sob��ֆ���SiQ��0�����yf�J�i�7��]kZy�*��A�b�<1�M�/�ks� ��)�&�r���R��Ð��GiJ�2v[d"�/�cE��O�=������=��ǵ	قd?��&�N@�(��ŲX��;�/�q������G8n@��(�=���x>�.Z�$��Zihr��r҂�JdC+�Ս~/�{7X���W��D0�h ���z��"$��*�x���˹_(�����=z��!�W�j4��'�:o*�c��Fa�
g`��?Ԗw2��2[��!�R���gJ�*��/W���4��%=�G�4)�v�q�̥��5��/�c�@��ԗ�"g���V��wdz��u�^_w�S�3��~���k�]5����0�*?���t�9�>%C,��E{�{��2��$�&A�z�����zuٮ�cl�Ϻ#�2��+A��w8 o���M��/M�p9I��N�_ٸ�,t?KF��{)��q�㍾����R�����fxF�Rw�����EbӞ�[����԰�anSl
-�U�N��V�.��pb�����n�y�>�-g�1�����H1�q�ː�"���j�=��ƌ,ԅ�M��8���GT���t�۹�(���RM�K���4ԒC����V�HJp5�n����0VX)���tF��Z���(>և�H+ 8�F����窖��g�*�o�U?k9>Ȯ��2���M^d��Lȉ���rV�Чɋ��^��%O�+V�i�(W��jҳuĐ�ґ���@��Q@���Vs)�Lw�kM'&n�m�>�;�zh�ot&A�ۓ�@��pXxR^1���6�I��G6XdM4��Oi��!�"��|��_M��2���ff��J���udBin�9�����<Y]�@��n�S'�d�c�Cn̼�^�����V��3��\�k}8�T�>���
�|��0�E �^�,@JD���F��g`�]�z��iQ�,�a����k�0'~��<�����e��ϧQ�赴���$�ɻ���O	T���B~�>^z\�������C����謔�5:�>���d��O�4�!�k��\��)��:?��:ړg�:Vr���$A{������o63=ù|��P%ZN�#0"+MW�|-|=ps��l\�@�1�Y��3��,+	`G�#y8�_��;lDwgK(��ֳ4���a1����;ZLZ�LƄb�w_1�\`�v�V�d$�h^)5ܯʹ1�A�ޤ��`{l��@<d3)"LH``3S���'��`��$�^�w5��������%�.�4$:,����g�~�X��L2�Ž{�έ��AD�%�e MY�����̊k��']y�םk�,�U)��J��[��QTyX�t��)2X��S�9_�=NS`�-�^E�_��#���/^�k���$��Gj��>U���t��I�	y5��y��/�Y �zH�˿p���"95�U�/_�[��V����#.i -X��ķGOˁT����ğ�pj�:Q�۩'V�y`�s�o�A��:�_n9�i�8�0�+t^�3y�YLd:@�AQk����f;|���pBQ��ș}�����3LtTEE���pW� #��p�w�`^d���0�o|B��%60�t.X���ޡr>��Ҝ�K+�Ҧ�X2,��R8��*^wD_�P��̔y��,��v|6?�R�;���9��79px�X{�Z���$�(�F��G�*r��5��y��a�?�-h;�L`=��]+ϊ���9�j�f��鳟�"Þ:���\���m����S�y�hjp�������2ҧݕ\6��q�@�4�7��;C�G2�6���&���?��9�������s#����+;��l$�����5��ɖ�ǝ+�Ի�<����nC`r�{	����{��tx'��������Y�V-�t�E?��n��e����z�|�X
��W{6�Y` .���E�ʀ��dc�5�
ML$��EZ�0�z���Qɇ-�(̷����P��\��W��L�d�~�E+u��D
Jw�/�y��2��E�q9GV�R�#|M�Ц�m:L�(�;���>�<�+�B�3XG��h�r/,�}g�-�t*-�j2�v�b���픭�S�y1.k eh룍�-�G]!"���#��)b�ۖ�XN�-�0�M�do�0�aCxe�%`�l��<�ICҝ�Bn�(��8�	���^qi��y���Q��\��%*-/)]u��-��������E�>��ƺZ�P�]��ս>#��;+�q�F�hG�4��L�(�\��Qz֛WFJ�&6�ǲ��q,�=��;�z��4�8����7m�}��g����+OBm��Ű\����* O��S_^Vm|��s(pҫ�h�g�ͭڳ�C>F+��`��×��u��#^jQ���d��0��h��|����B�zl_��%��Ȩ�x'�w���Ψ�����O�[�ʕ�ˮrq�;_����-�f;���^��}-��(B����}M��i���}d�U�k�$ Fy�8���a�Q6���C�h^	b<^�@���1T�V��XM��(�#no�!7x�+N��z��0��]��j����[鮁��xIيF�{�r�N)��G�z��.7��7��H�+���⯁J��� ���Ĝ97z��
m1J�WD����V��j�aI�Ut:b����4���2#�.���>��6����h�#+k��[�fU�E�U�FM��u��#��Ɍp��zx�*���2����[Z���r�.������gPt 8�]�;mwi�҂p���d�lx�=@��+Gg�_�Կ����L�?�s<V(51�,|��K
r���EYK)֜>h�`A%i/�����Q�e+�\�Ah��2�m���SH�e���]�À�\�����L�(����K'��x�g�Rh�䭖#k�xo�Sn�g�*�<$XN����؃�7���e���M��,����e�sr���W^@Hm�C<R?�ϔV8 �a��[X]�jaŧ{���q�J�ǰ����L�d����'�+��m)�i��t����g��Q�J�4�<'�����8��̜�9���j����9��:Ǟ1� �����̽_(��D=έ��ũx���V�F'ሢ`��YE��j@����(H]��[Kh�L��7���¨U�[>��=>����gi�wv��z67[y��0�}l��2����*hcs0{ f�X֯�I[)�+����ʞ��B�m�Y���%v���p���^+K���\"�9v��o_1�唱x�$����.��ٔ՞�ι�>5vy��x<8n��ey�����Q��b�_�՚}�����^M��p���A�[t���|�ׁ'-�������v�8#�U��g���U+ ����Q�ǳf~�<\�@2�
p��g�w�պ���q���Q>�	�̰��]��G׊�A:��z��3�L��#��К$S�44Kj�.d��f��W���������-����J{��~~�.C:C�ȒԳ6�&v����a�F�sn����T�����ս�����@���ls��ڏxumW?u��`^i�ʁly�����q���X�ɯ7�����U�>҅�q�0�ݬ�,�7�>��8ɠ�}��)�=�Go䬕�ϑ�s3,�c˖>g�/ːz��1���5������YsZ��vz+�x��m�Ci�R�1�v��cq�+~+�)/'�;L�v�8d4ųq{�RU:>���8JZ��C����&U��@Z;�w���5�+;����4���{����q�Z(z�R�My��^�����;4��ӳ~�sb,|��c��Z��`G"/�pl9Z��㦐�d	C):گV���K{)J�m{�1����=��_t�^F�vRfi~C�>�d{���Q�x�X�m�U�Qޥ��v�RHwZ�wg��oa i���L<��-���n��8�ܟ��H�Ñ	�'�̫hN����Y�3頋�H��;�݃�Wh@�{�W�ud9㥙�b���j{	���Lq����$v��Lzt�-І�Q�d�q��r�\-,�r_�sC������@�dm��r+|����2~�#�	W��J�ª5.�� �)�
�wu�t�B��{:��Sb�|3���~�⁧[�?�!PxR�)���5/���ţ�ҁEz�K+m���({�H��<ܽ���m\t䠍wA���p(l+����Ġ�.o'���E�3�\���e��]�H�����K�����a��kW��1�QzK��\��.�9i�醧��N_�V�G�V2���6]D�ʓ,�5��� �����%ݱ�u���O�k`u&������goU�}�K���!��@�����A�XO�y%�噳n�@��q�Le �4`+���\\����}��E�I�{b�u
��D���?�J`���P�%�u6��X�yWcLhwW��A�ZH�=2�e���򹚳�LƩ�'�4�ˑ�D4�`�ޛbA���A����P����}�����R�}"O��ϓ�u���G����zR����1Fs�kY> �bX�:�<Ke����H�)밢#Q�rqT��m�� Q�B���@����`����>Ih�]�O��+�o�?`��Bo����y�;ןEg���άH��t{���֫����|(7c�5�=%�+5�f���}ytJ��'u�����/*��Ծ3���H�����!�2/e(��|N"�#�c��^xqX�`g:/y��Kqx-�5����Qʮ��-<���ފ!�n�k�P{����ˠ�#l���ƻ��^8۪���~�������@��}%�ge	 �<��"�7���a����aQ<;�����CUN�
�����O���j�k����^�~�Q��4���yTυPVJ���#ڱܒ�Tzf7��C�F�c�̗#�vS�}�M��v9�%/|�7/��#D�Z���2;���i-�Wj\�6�w|#�s0OS�TgM���Oȴ��`�t���oe q���q�����H>���������i���7��'9mDI!�8�[�s#�l��iê�O௞�D��,��nO94���������Z6��Bt�<[���Z�8D��k��C� �P��;�F�Q�b^ƹ�nw��Ґp����)�R;;�C��Ŀ#�k�u�@<��ra~\�*2v�*�Sβr-<>p<R�qkx���A�-ꁟ�4&#�G�6�von��r,�S��3͹/���?�>�ц���N���`��r�f4�+igJ��*G�+30z���W���Z#>����	�8}�5=CM\���sE�o�L��e ��Z�݃��_WD.��#�H\	䱑@�~Dp�q��[��I��O0'5=�a��5#����3�B�x�U�੝�w��K��MN?V.�ĆYgz�|jh�7k���C��2���;*9y�����{Vp��C�C:��Y8?�%�T-�%p���'э��+4�xqԵx.>m��u�[�nK�g�����R�'@�[�("S6�V��@��rГqP�h����	�o��c�*��q��1����A�t�~4��w~u���#_�Cm�;q�_�@j�&�����	�����R��p>n�/Pc���+ͬ� �բ���g�� =J{��IL������=W*{���+�ۗ��ݞ.,=k~k��m*��k�@F�"����o2�@��������X�4Ȝ��{�3~�l|7�;&oj �G��$x�)A�F�+E�Vu�p��j�œ��?^�|Fy
?Y���1��vso�i�z�[h��`+����c,)�G�
|�aE-��`��H^{�Y�~S��x����R��K���I������1~�T�ժ���`��کn�>G���������+8��m-�",wJ^�3��w߆@�%3d�.�*R�v��؊�1��������Q���D*>��96t��-תz�+6�6�8:���tm���D��tkA��~������X�Q���Y�b�����3��t�|n���aHI��Q;����ϛ�n�KH&���P�6[�|'��a�u'|��e�� n=s6=��C8`�ڶ+���/	�g{��`�B?���f:˳��)z�sc���N�ἏS��c� �ְ!>P��m����[�)����7
�8��$���s_s�΂�p��e,/k	7-}��^����2`��EpzWjo�����y-P@�8�; l�-cCB��[�;�l�>���.l�؈�2��&v����3�Y|-h�G��]@��҃tz]�0�{��@�9����O{�+`X�T�C��b-��G0Su��{�H��ƞ8�ia�=�R��YX�l� �Z1�}��̔�!{�'oz\U��e���<����}��ڍ������e8eN\I2���B9"7up���+�S:� ��u����)W]Ŧ�x3�� ;��"|��R��g�8۩�/i�V����������-z������5Johu������w0~_���8�*4���'���n�ǵ~R����.�����.Ԥ�9�@9%/����ƫ��ob ��gbo���s�IIg�[��.ͼi%��?E���G^�&������Ap��[�@�k���А��� �=ZJ�,�O�}Q^=»>�RΜ����+��\���{��5�w�宀�2�n��L���L�l��PW�_o�e4�i�}��[���#�{ ��֊K���Ûy��CB�J$��U�`g.`������°w���<����I��&E۵� �W���p�ܸ��� �M�+T_��0����k����a;�g��[AWg}u���_�m�w���>��[/%^��O(��q��5)}����8b��R���ӽ�֧����~7���I�82�o^ג�C�Jy�O�%�� g%y�r��/��IwO��}��*��I��;���#^l4V��p�
R���]!�I��d�|�6��(/��JO�KH���w�9_�Y�����LC�$]�t�K*>�H�j� ��<��q���
�>K�b�5	��n<Ң�����ħ ۸����l�G>��?��;.��X���"7�!0sC�JcL��|j^qV��;}DM��m��
W\9ӫm�-���$�>���W�@��Ԡh��e#��}���Y^�i�h�^Fg�X]X��b8��'o�ǣ���[Kj?��E��O�<�}g"S���<U�W�'>� y�
D�>+��n�9c"{<���BT_��~���b%��+��qg�v�pg��?��·t��$�gw.i �b|�=���_�UKLT|��/=ш�$��/N�㫳�z��:��~+�A�+KpO���F5I��+��Z��,���S��yd�V�C�@�PKs��lz\?�HB�q&E:}���c�R���EX� �����Zq:<��H�uP�En��΄�{+����O&?1�e��]//��Սף%Gb�{i�����;��Z��I��X�:�]V;��#�>J� Q��]������|��R{�eivv0�����s�trА]}z��į�ܽI�y���������C�Gzd�����ęΡ75��D�^N�'�u�[7���j�Ua
�R�Hw3���Wa��  gx�y��n��O�G/�H�q��CV��k����n�}�����]9_���� ; �(F�C�:��춾���/��w��-:���(�}�k�ŷ0��dK�V=
���}�g��q����'�]iO]/]g�x��s˗�_�Yw�B��":h�PX�����7eQb��?�}@z��-�#�)]g-ۚ��b���E���zo$M���QحiP���=
��0;+��X:_dcf�SƳK)�@�k��+��l��
�S*����'ZJ:��^�ҡ";��U���T�~�^��8�6���$��;����:TB-FVVdL�� �0��Iv�y ��f\4x���%!n��o�v���@CU0�)�-K�� ���
�gV�bá���_��5@%�pE�ɥ�k���C*W�Ϭ��ě�Dlr�W�1{����q:�\#�:+k0�*�s��L=�th�NSӳ�O<y5�R:��A�SZ��.�,�hwI��k�\�`�"��o�X�R��?��tԲ�l/��7H>����8��#H�V3j��7�k�1#�$X�_+3��?CY���L��ܹ�֫x-��)��?~��hlαm~m�z|/���)�{�0{�0�kpe9ׂ���s��KJ�X�s1ɧ�<�1���{����c�t���v�t��g�}~�Y���̺�u��ϸg�m��X�� ��@���;Ă�b��l�d`���X�B� �kcy[43̌ml�=�ޭ�VfFdDd䏪S�:���}頻�̬���������S��X��I���J�D|��+{3H���ok�%�~u�)$�l�4�i-�Cc��9!�_�yy�a��0����#YN��E+�j���1Q[,Ԁ�����,��ky�������ц�D��Rm�����87i�ؚc��L�st�p�R��꥿����%�:�##�����f���Ez H� ��X�~��f�5��@��M���(m�pE�g�B��FV/�p���+*���%)�Q!Y�[�{��=?�u�$D6�\�#nĄ8�S���j�M�6ۢ�Fw��G���9ܳ���e(��ZgB8v���Õ�3o��p��m{nO�(�69�9�C`���qg<�[�w&��<��.����לA�qt=?O�'ҥ��=�4�6�X�q/ST�`�8g�s �se��Q�5��đj�^�Y�ڵ�*]H'�^%��й���к�ui�20�[iv�g�ȸ��k��-�q`{�%W0^���t���y��k덕��䮱i8E@]�{�K�D�(d�����1�FX^��%�GӁ���0�Z8�zx�z�㮠��j�F���]/୽���� #�4tBW$�@�/f�&�ka��{����{��Q�z����8:Z��!����Nmޚױ�W|{V���V���j�޶���0w���T^4F�(K~>T=���5���2����樶2���˰�k���W��V�ca���q?K�Q�z����^�Z�/��f���.^��-2T��H���#��Yy/�T1�kd|:� ]vjD���z��w(4�I/B�Ӭ9P!�)��L��^;��݆]����������B/H����<g*�}���^H��b%f�>w��5Hq��vi����{���<0C��}�*����{�3�t�+I�g`7E~a2�1S���b�Oӽ��i�=��ȻJ��fU�j����ج�+C��!����F�1�
2g�p^��P��
E3e`v?I`յ��f�Pk=n�,#�|��i�k.g 	�R�ٴ4=��=��4��g'�O�=��
&$<wrV��q"'c��y�T��C�10���w%�1��p#�
a��2��E��cǋ���H����%{�'���cp� ����d�ܣs��Y4{�ω72r�-W�@댻��m�"Ֆ\��/g EO�Gc.�ñ�@N7���`y�_M\��I�~�Q;�������!�\4��$F!Ofw�����48\QG��3��c!h��988Ϳ,\[y��PzC��.nj���{�[�yl;\�;�N\iT ѭ��ЮZkڪ"x����SX��%m
s��dm��b�W�\a��o�ݦ�.�q3���귤�|��h���{j�.F�і��z�:ҳ�ʐzr��96C�Lj�9z^ @`�p#�K���h%���,�$�����=���\�Y���ص�9{���	6�FJ��F��T&9�B�D~,̂N_ |Ss@{gR^A��\du�D�p'�2���,��:{d�XF��=����%�����q�F��1���!�| �Q���Bhx��( ��5(���e��z�m{ץ2U~�ᰇaL����O���H3��P�F��EP׾������R���	R
*��t��5���JFsP�!ӈ�:�E�~#�NRR�QpJ�љr��-t�p�u<x4��>��n?ϫ�A�PB+ĈO�%���Z.c �v����(�`�1��H���f�P`��9-�\K^fI �b�<q��^�f�]�躤��୍��������&*��9�t	h�U��œ��+�zA��>)u�{�x��ӳ~s�\yt٭<X2��m��c�جSmg��0�`ȭ�|����₀�r �w�;Y�:�`���L��ƿ8�!ϲ�hhP�Y�1�$���f����%?K��\��F"�Q<��7Y_j��`~RSN�h�Q|��M��@��o,�r�/�x����e���H�G�V3��ᲈ����
�ܩj�$�s��Sτ��bt]R�Z���_@���&������V���O<	���u��ʟ��Uϫs��cK_�U�1à��6��3�$�nJ@T3|AP��Dv�EK�}��C,�nx� k|؉���<h	�6��*��o`P�Fl�j�&��p����*��6ڤB5P�'���H!�|��$9Q�W�?�m��y@AyٸL,i��h��w#��"�!WEky8.g y��(F���i$��^��[v$�Gn���L���1��>�i��`K�h"��&�4lc��1&����
!�Y��2��b�~C��.|<���2\̣�+s�;���-����|�F3m�������|}��I�eޟ=Rv��䬋�i�tI�`C�Y����>�C�OG�#�����m�,.���I�Q7��|�iFR����{� ��1}o��pYL!�����b��B0����(�f�=�}�����v��-����0�_L��p��� ��;	�-j%��ճL��eV�4Jf��ݟ���j��T����J���@E�ǌ�'r�!HT
��.ͩ��<^-��/.���h�Y뎀�6� &�ض��|&��4�p�߰�}q��EZM�C��Fk��ߵ4�J�-�!��/��E��M���tnx[Ͱ�~�깪Y��$d-GXJx�,z���{�唂��8����Sy��$��@0O˫�ͫ�e:V9�?E/�C���5�6XX�FZo)����}�/"�EV�>�����5�_�ɷ�>����n0V�JRG�^��ƪj]�g�|��I�B��)�#�v!ے��7���'�w��cu�Q������l��tg%M���;3��߫�2���F+-*J�@S>9a<������Îb[s��h��Z�+!y�s�7'!�u[3�����M�)q�ӂ���S��d��|S��@S��xI������B��M}.|�JW@��1dy7�|T�������Zc�r2숸�����Y��D�| 7�rtp��J�3h��O��H�HZ�uv�0q:T�;�}���A�e�e}	)�]Ԏj֬�ݫ�%�΄�f:'Dg�p��9�@��ƞ6��sSE�+Oa+�\l�_Ī<�I�?�<��QH|�	� ��:Ɍ�uJ;�i��bp� k[���:�Ӈ��ئ �]Wn;▸ۿq�#�Ix�w)7��m�<�is�+�5���b�L�������q
Yec�BQ��^\p?�m��h��f5
$}.n��5�'���X|�Çp��9��l�v�i{����hե]��#�0��i�m+z���	���z�82�>hP�	��9�5��$�maY*���8En���+�b��+c�W���!TI*s��z��A�`fu{$�ދ���;��B��{"�EfRYo�UqlW+�Khs��J?�q��H�Ϳ�¶a\�@�웍NC��h0�{���ۚ��^jvA'u�d��y�a;@L��a.N����b�4�=}2��e�FV��G�=���Wt�"�VUR0\^�?�&3e�+S��/�D�@�v�4H�-}�Q,^���p���0�:FΓ�k9�+�Ws~"�"�;�6E�f�o����r��_4e�VyY`��l��2y#�L�:5�A���.�携3�)�|*���m�,|k���Ѩ�F�W�׸�g'�T8 Ȉ���ɋ/�Ϝ��-D�P.��T�PT���0�}̂v�ӻ{.i �<�]R]Ni!;t�hƖ�p��U3"j5����%k��j��7�pE�oݦ̑g�f��/ܧ<�TP��#Wf����=.i�ܺ�N��(��|R���glw:�5||?9XY!tƻ�޳��YF����o����o��9���+�͕�Zgkk#��3UE~& S�U8%WT��S��+��1?֧���5��;u���v0�3�OkVn6 ������q�q
9tS��6���4ꄼq�gT�)�V�C��Ё�ܖ�}z��l��4%e"XI�x��j���~(!'�����$�2F���W5�i[��Lۉ��X�華W���$��q�0���A�U��>Ÿs�bo?���w`q�EO����Q`9N�e�0�x��,ܧ�/͋ε�n��լ�|(m2��w��)�T�P��m����TcX����v�����;��V>;@v5)HkI��W��Պ�N�6y�u[���PO�-c��;��{�p ����ĻFxKV�(<̍︵������ �=����U�am�z􂌙�<�=��������!�"5�<��7�ƙ�q9صO�ƹѱ�r1���t"6_�����?��Z݂hQ\2N���}<b]}�H���b33᐀t́�P,h�k؟�KH����(2�AɁgT�4����xv"
t�2:�O��߫17�y`��IϢ 1pij	4#��Ng*x���Y0�V�^xw	�7�X���{6�PL"�G%;)�>�ߑ-�i��;�aٺNJ�GmZ4�C��S$Q�7S�4#*�S�5lB>:�G(�۪��q-2��ۂε�E���u�e��/R�V�X�����9R��݊Ǟ1�J�F�����,/�lO�}C�W*��S����,�N�h�>������W+@�r�b"�q��`ż&&�V��V�r�b,�
P����g�x��E|n�,��L�v���0{DO%]�0`�ި�t?���s������N��e�2�Hy�,�!�{��sQ���'�[�ty}uM-���3�!]�@�4��|\{A�kj1$��H ��ם�⺄ƯL���gj�E^�ي0��<�Ӽo����c�ͽ�[`\>�r�.ox��[�t����P���>��U:��J��t�l��++��]^6�������S&�ϰ9Z�o&d��|��������63�ļ�o�s؊DV��u܄�&����t�ޖʹ��[vo����&[��aV$��������;
J�f%i��h`
E�A2�g��T%=fU��G ��g���T��^�_פ<�>�:b������vd�OK
�8p6=�<�:�:l`��ꓶ�k�_ޠͭ�ki [���/�h��+�٦��[n��b���xs>)�Ʉĝ(C"g��Ρ�t m5^Wɸ�*��O�m���:�c�D���<��6���9f(�TH�k��A	@彳�s,-��"�d��-S��E:��x�̀a�n�)�j����<�F��M�k�<�ĽРE��R/�$h����?3�cQ�!��3Hhؙ�D{A���C�!~�[�m|A���3����
aR��|j�Y�JI�[D���#)�$��w���(�L^�}ʚh#��лc�=A��b��"�#|�>�����pI�)���оl�L4�.l�;��r=��m�3�n2�� ��O�+t���8
h!*PX���1v�Pk�+T¨���}�dAڇ!�� �pO�����E�*��ľv�Z�B0TW���睞��<e�N�E��px���҄(1XH�aX�G�I+����V�.�"ˆ9���t�Yqg�ud��NP��6�n�}�y'Hl�M��iN7�SQl�s_P��4��xG�"��`'6;��Q�� �f��7�D�1�Ɔ��\7wO�M �9�~s��N�	��m��p����1�ˤ�=Ǫ�JlI�Z�ҰS�)�X�g�q�DCy�Fi9��6��+�q��c/����!��Z}�'�xΙ�n�����(�]�m+�]�=2���-�2&*�����]�@R@a��l'����V�8�QГ
�m]�;�= �Do�u�k��x�CW�{UJ%O'.�S�s �"�1���fI�ר�m��C �c"e������ҍ����.� H-��A,"SIm���6��y,����U�r/��/��:�-��>*\2m�����m�C�5x�x�VhST��7�sb�)72������W�|4�R���X�iMgh���I��}i���fH�F+�@wj�k��~c��*�$p2�d���36��qWCZ���a�i���i}�x�7�����-b��\�9��۬/)i���/��\�i���'�5�S:A�u�o��#���Y�a�k�J|D��d4�-B�.�sP.f���2�m�_NutrІ��O@��G=t�k�I'��;�o�$#�u�]�0���,>n��NZ���kjeM�f�nݾ�`�T���G���X���uSr@�ȇ'���7�a".�;r[�j�0ي���:�����`�ȃ+�Ҡ<���v���(ّ�j��77@�!�?I��J�Y.��G��|�m��
���C�X1��R4W×M���l������+��L	K�+�j���5�}lm�����l��.�c�j�@�G$	��Y����i&��������l���Ljj�{����n+	�WB2ė`(mҦ�-.� :��|S>�{N�o�2�g��QgT����l��O�5:]�=͌����$KvOEf�7o~!���qm��5�b�/�ã�Υ ��I�_��ӶW�!�یђ���7^}�Jlmv+�u9c�������c|*4e֊�a>�.�K�{�{�C��۩�I����J��3��S����pmY�����o�[(�d�x:�:�1��V�]�H\�̋�R�1��|Pt�C2Zc�g0�	ٝ����"��k�v8��	>�s�-A��g �,�5���2S���?RFa�bkAe�Z4o-"s����{�Y� ���ni�έv��e��)�م���Ҡ�( ����Zm&�6f��y݄d(\	t$����z�'㬄���t�a�Ѧ=[���8��=>]6��-���V0Lå��}��j���=wc@��ee�Y%��N�N�eE�o��׸���7�㼅5$��s��2�5xZisN8�Q����F[�&�Ц���:�&�y�� �T]H3)P6��l��~�&z�0���Ѱ�9��y�X�/��a��OPx�k��]ѮD�^0�uEE��X�7�=}�v̊3Gi�Ҷ0�-�*��)^�Q��o���{���9�9*K���Z;��h����l�G������_����5[Eb׽W���2�gg9O���;;�Y�z����
Tf��Y\��f��dG!d���pC#�; Y���&�\��W�����#r&ޘ~o�j���l��ry����Ӻܐ'��Q1g�c~ ��� �7���U��ϡ_�ͅU�k~��C�J�鸞��1�oc�|����k�^�p/^�Nax�̓%p}��+�I�g`�>��X���/=ߊT�gjW�p��8},��.��}��-����7�ͷ?�`voaBX���t?���ޏ	Tr�?X��V�ޥM����͇���o?H�s�\�!b;|�q�������v�E���_c|We�$�`���O���hG��Rߐn�
ɢ����}k2Xb��?8�-|��훰�*���ֈ���� ^�eҥa;Yi[��{y�l|;�iJV�Tʹ[@���~�3�1�����	��qN-l���M��*4���k4egT�իm��y�����&�&^��M��Q)I�?h~�����R��i�_��\Om�C�,��ș�X�n�$i�Tt��r�9!b����dh��ϖ�%��d��/��4��{�j꭛��  ��e�d��[.ė�?����E�fw�xS,á�A@~��6��N��x����|a4[�͝���J�Ş�?.��Kxߜ]�E�0E�����2gb��a��ϗ���w�&�;�����W��:�����}�ڞ����$H�!��3L������z�7������fAӦ��J7���>��Kx!%�!F�L_[�v�v&�Aj�SQ�t3u�)|��̟Z�;��^ 4k=eO��G�������C����wܦ��A�2�3αj�r/��(�*�'���{\�e`��'��}�'�䯹�(�ZS�B�����7C4����!�qIP
�F����o����G�׭<��_�Em�Ř� ��F�������~�=Q<sҰ��IaQ�f�4�U�>�A�.��=@%m{���Y� _KPҕ�#*a�s?����'���7q>�q�n�W,�)��\�X���M�0���'����l4o����_̩�=[�r_���
�������)L���}fn����UGf�-��σ�kM�4��y��ƹ��h[��� �S���_~�kmY��e����vV�w����K�!���flY#=�Q��-��Ŀq�ʀ�H7�h�������-�fs�}��f����H chu�8��c>�l�r}ޣ����v��ݒx��O_~�'�ۯ�ع��,n2��ݒې��_����w	)#���T��X2�_�<����(��������_D�/��@�΢,9����=�3��CQ���oݼ�K�\�R���
x4��J�}J�;�(M�pǚ^O�ȧ?�B��V�`Gz�4��mXaЀg��;ܹ�3�P��~�4�=*���ýy�`R��������GE��Uf���Ἴ�I�l?����[6!�wk܄�;$��mW����0X��s;G��Cj��(k�l�Қ|V�[�z2�q�Y�܁��w����)����[��ے�����	�7�����@[A�v��JLa<��a���������	��(�C��Ū��H�|�*3��J�����}�0`Z�^(��Dvw������� ���7�w%6�Ю���<�����`D�)�ɼ��mv�'�:��خ?�3e���Jqu��8�g�#���u�U�xO:�����6""Uo�lkp��L��n1�6����o�	�J��d3tEm>�+�u*�ы akxs�w~��s���6C;l~0Ю��>3��_�h��M�&Ib���-d@�YfEgϙ+o�K���$���Un(A�r��.EX]j�ͩB>���t����M���O�p�-<ƣ�\��F�ڊW�ާ{a�ds Y\&�A�1�M��굫��e�=�=m�7�������pPZw$�o,�����o�:��m�Kڌ ��>���>�Hb���6]����h��Hj��1�o�צ���f\��k!ީ<�+�2�v���kN�U�/3[�ɕcO�am��5��Mq^ ���$bVH�&Ic<�����[r{��^Rm}�7���j�F7�*�]��b2F�1��P|��5�~�O��d�Up<2dx�y�[�e��W�ei�����<����B���p�1��TL� ��9��Jh0e S"$�4�v�~c������4�3���aK�6�� ö��+�	���_����0�5�Ժ�[7�8��^�����8s�(s� ��4�\C	X\��e�K]+쪍����6�66�C2����$���#'
� Ƀ7Q.5��(��z`Y��k_�A�_/ׯv@�;pF�*�: ���
�1�d&T�N���8Ho#��oOۦ�z�۔ü. �xb8}���[���̟�YcRxzӻ1!K���l4�����Z�V���w���.W���<׬���-x��hܘ`Rd�%�6�����F_�Z�^�����X��s���ؾ�=�����C�Ŀ4[Ǐ�BV�������*8���ɨ_C�,�g�22�\��k߉���8h������=�:��B��B��.�9�������k'���(
i|dFȆ���A�iJ;��_F�����zO����c(Tҁ���h��j?�iŚ����|P���I���Ĉ�M��6�Bܧ�	�A�a�2t&��f�I����}N:���J#�`������F�Z|	�$�v���:�iu)��nѺBo>�n���s���=^��1��ñʞ'yZ-L0��52pF��	��z�wZ����o�3���н3Q����s����<���޾��6����3I��5� �T��|v�`Q%��IS���,�^G�:p��u�	����6�i>���KN�w�Z�x��t{tj9�ܗ&[���6�[c#a{5hf���Ĵޝ�B=V&xSZ̝�|��בY�:�"OD�2�J� VD���MpAe�r�wC\D��/w�vp��
rSķ��) yjy��P��X���&�g@^��$�!����f]9�� (w9$cI/�;���Π5Ft�es5c�H�a
l2��C���R�("���@�z�M��k�`�bP,h�oEI���4�ؽv�x��7+}��>ˤ(ˡ�>��wh2����i��jt����8-�pL�y(�a�R[#��0�$�x�	���87��&#�fK0u�J��YUf�֠wiſ8n��5�ux_�HS�}G_ҙ|ɡ󆡶�G��k\g��<X߱��9�b=���d1��%b�RZ�l�eSŞ2���/V���37�M��3ͧY��Wv�*D$���<%��ҩ�ͳ*G����5��6�F�i��w?%Irdn��sR�ل�I�W�D�&�iY�����3E�Ɉ���7��d�ѥ��n 
�~y�:���H[S�/Q���4�B]�'��x"ƚ�:pBʫ�y�v�A�S$�(N�[�*
��-�6���}��g���Ly�����f�Fڗ����.���	���-@�ΰ)�g�R�<F��ƾ�-D|
� :��iP���+O��;g�;��4$�wB-��9�@�'8���1���Q�!Y	%C�s����٤t��؞�i�p�Mnl���-*�f׷�/ME��;���F6x�n>Й��V�r�����K�4�	�l��5V�ݜ�rZ��������=���!�����:���Ί�A�$Y�&����_��q_���`{���MQe��G�5��`Qb�S�v-|�F�������e���u+����J/�G� s�v����|C+qV!&A�*�IrWcD��T*��e>� ��*�?ب��y�O����x4�YD��i-7�y�v���K/{� �����뀡�(�=<�P����ޟ�j���є�>6<_D��,)�dL�z�IU��AP�1b�;g_�~�+"����P�-�!�E��")�*������p�[�'e�O�#0����^7���H:�83���Jf�%{� 	
3���S�-�~ϴO�U����"^�#[�Y�v'�Ћ�Y��N�ۭg|F�M������܍���g���,A�*E�p�.�!ߵEw	���*i�hVT�n��`�l�Z0�Y\�E#A�{"�رv���W�>�3	^D4������'��h}T0��u���]��a���օfo�I�|���0E���|�x(������$r�:~�2H�4[��ٖ&���tw�� �~�L�(�=_�f����a��Do�����h�i��:�$��+6��9e��B���q@0��Ya'Y)��NK��F\��J_��Y���8�9&r�3�:>��gi���X���M�c\�瞆�H��!h~����"�h[u�������r�_��1ԣF�0������rA)f����}�.�T�Q�� J����}2|��Q
�v�Gu��
�c�ԿH�)�IG�� �T��
ꊏ��bLwF\�� �(SP�gD�Gւ;=z���o�^>)�-���cxv-4�x�0?��ޫ)r��P�h�`�H�S�o�r�Q�"[_虡m���]ۗ Ґ�3�!@㌜�~5E���r�k��	�g��f4�����3mg��� �ƫ
"��?�q�\yq])@�뢩V��[ �5rb4��%��V5�-Rc�	��u643���B���HE�TmKL"�x�?���3͊I��:4��	�W*u���a/������*/�	�i7�[&��.aB��yiohv�N��E;78{\B�	���Y�w���Lʨ��y����_���S�)�&d��C]\��6uӒ��Z�o�Ep�v���U}�M��
<K�^{���N����V��)�����~��ָ����;x�0�X(�.?>9JA�aش�{�����|��v�<qW��Q6M��^�`�
���*���ږ�\~���Q�!G�4�#�D������f�T�.m q~���0��
�U��Ȼ:�/�p"1��pahZ�=#����+�uR�*�v�՞��/L�Z��4��^��O�:���KdX��v˷\�_>�-�J�"��M��n�C�-�o ����,��1㟤�YJ�ksz�cH���ˬ��r�vp�2o�cS=/n��L�zF��xա�1-I�6�O���s�
GJT�/Y�f�r(=�m��r��oz:��{�|�IsEz�F��!�k8p�wU��d(��8m����6BVU�#g���޵ֶ��k㽣<����҆1�
�{��A���+��+���e/�?�{������_Hڌ�3&i�
Z��UP�mh�� \�-�����2K�7=����i����,L�@��BI��@�k��mhy��{]eL_C,#li���`�����&��yV�f����j7*�s��u!5��W(�١�Lw��p�T�X@�hmɷ/���hV���ߣ�ÝW��^>'Bo~�4�c$J4����n����P'Tٳ����v�����׏i}��{y��C!.ucr?�.����l��>�ې`���qD��[EĢ���1�h�_��д���Q�&��v�Վ�����N����зZg.]���3�-�r�m[�	7H#��00���]�=�x]�!.���E�>��<�p���%��Q��æK�&&�*h�m nߏ���-�L���H},w8�GQ������C���'��6�4-�va��%$��!���01'�q-]�qǻ"g�6t/g��=�Ŗe�J�����'��S������#�ғ�g�m�l�ْ����0õhyp��Ad�J=�/�� �7�҇�z�Q���wfN�pT�;��;��ۦ�kP(�\%In�Q�V`�:�!S	F���r��W� ac?�1�����¤~`_,�7���Il�cZk-�jT��t9{�W1@kG�߶�5��?���ԎԽ@�E���/�;ܨ �sצI5���^��/�m���z�t�qN碠����ta<��zC����m�_.�S�뚯a߻2�a�<�' �_b�����n�.x�����q>�u��V�C�5<��
X��Kb���%l�,v-�8ؖ��x�x`)�r��gq�o����ZU�Na[�K(��sU�~�����sj�>]s�Ef���ȄWg�j�z~3c�ă�^�%
��J����$|v4��5KΉ˫j��Y�E� v����^��A������+��:�ʻw�O�o����L[�r�]�9��-��l��u{&i�u'����` L�Pz�����w��@�p� ^y��]�6�rlS���:��J͟L�x�LA;]52�gUXu�����Nz��.�8�r��k�<t������sc_e;�(�j.꜑��|k,��EJ��a�}n����R�S<_JV:���u�@*���9ҁT/_<�G�;�'�ez��i=dڧbc��#־#do�"W}������d����8�(|��#�Q���*N\w���~>�	�/�4;����~r'T]��Իg�5�jxX^'�ee�o����)���"��[�\u-�e���=�a��:׫˟y-ό�Z+ ������^<���TW����_�;Q;R*k���z��P��!Θj� qG�����LŘ8h%x`�K�g�0��~���V=��qV㇒5�-�Z(Ş��p�����7;�O�A�s� ��}�!��'vQ7�o�<>���)��C�	�g�'W�e�eZ��yYFJW��x�ȳY����|��S�Ow�Ģ���%=>�]�E�C�k���p��|عp�(�w����u�/E#,u���Y�=z�^�xeN5Ӵe,��a��?/j m���`�ڙ#'t�IK�?��s��ء��,⮱��܁�;���ք�6󒡣�B��3�9k�}���ݯæ�K��v���U��CUMc�B��yV6���_G�Ta9'vi�\��0�|g���\�p�����K������R�˙��਽x=��)*�����Ō�Õ�~s%�9�yG���i��1��O�͙u]~���V����S��n��n�������g��N1��5z{}��"-��������"��G�����րBu"���ְ������4�)�{.^�@ڀJI����i�̾��8#%wW��q���{��۲�3�֨��Ze��p�p��l��˺�8���Tu(=2<���w�kyŪt\��@8\�F�+�k��=Ҧum�I`Ve0��� uQ��X��+�sT}����������B3w��!HF2�y {q�p^fl4�U�1���Wu�}*F�5)���gK�V��'���j��bX��/@�Ն��Rߨa��KaЖq���lVmm#�\7���a`EdKE��j9B�h���=���N�V��܂-��$�������(C�����F��-�S9�c6f��2�l5�3uJ��c��}0a%X��
ٗ~ͭd�Y�BUg�+�ɸ�w3�h\��xc@��`h����O��z��ȳc�Z0�7&q��y&`0^?Bvo{�gI�-�������p�p@c�%���"HO$��'�q�n�oF����ʥz�TZ}4�	�M*�U���u2��ZrÞ!�َg�׻�M5�ⷷ(>���U�IXc�cHѐ%'4p��C�������]���I��^����`�\Y�j�n�J�~��Η�e�Vs��X�Z=)�X]B6���<�ư8R�Pha|<�I@�����lC{j$��0�0TC6lCeh�:S�r�h�ݑ�s�.h(����閻*��_��2�M]�4�p���ƵD����Oy�dA��rEx��<d-�wBXI� �6}������_���C��ې���۽���/�N.���w�}NL!rYu��:n��"+<[�6�\�J��I����Bh���1]6	��.֓ys5�^�.V��������p�@����NkY��*�}䷖��;����!@Y��m����I�e������<����ٕ��c�ã7�XW\?��*�%��z�v��}0��v5�H¬�yQ>n<µT���ې�|Y�n�K��E����}���[��F�O0j���v�~��K?S��6@� �=��^�SMD�!�'�'�%�\�O�"e#vdd6x�0�xH8�Q�y�.�{H[�3C��
����)�V�e�rA���:_֝�]n|�����󞸤���&!���������ʺ�Ӡ�=��Ee��5q�q�F���l�	�tw2u��(^��u�A�7{����Y�&�q����^�'�3<�Y>�ψ�=b5��s��+5X~_�kZ;d����`������LYryzI�`�Y���u���������r� �_����)��:��w6��;c�<���s=�7�������n��A�K�;��	�+Z����4xX����k��&{�r~.�5�
��S~-��=c�6���ʉv��=����SukK���7�ր��&O�Tb�e���O�Lq�{Ѩ�����/��H��pp�ԎE+Ҳ�θ�ʛf��rH��h92�c�� p����6;~�[���@�m��f���3T�N�+n����/n���4�1��U�]k�����O_B�r�Ӭ�+�Aʷb���J��g���c!vm�5f� ���%$� �a\��K��R���PF��k��T��+鎗ѩ@|��Pjk��}�X%���yߨ�O�N�:V��"[�r+��s���FidT�v:��~�V#űr���_n��\#Ɋ�=��uU|��铯o�{��Q�3+%�`�ߍ�5?�E��wZ�G�%��Z����ܼ�p0z��p@�����]�<�>_E4���,Z�Xך��&������~��9��c��u��<���/pI�橪���*�T:����N����:��a	:᩼��,{=�|L�y���| y�4�4��R���R�V��5P��U��u��Q�%n^��y4���W��1�+_�)y�H�9�׎��록N���B�A���Y+m?OR���n�Q+�<s�{��Q^�Xi����hj߼?nk���=��g1���\�(6Z�3\cLT ����%����-���]�Xng�x�w���l� �!(�S�D���Tf$9w;;<ӗ}Zv��� C�Z�w�kxa���F�68Y1����!dx�*�)���0󼚂r0��[��ˮ���$0���cz�ix�U*oW�7I� �:[�j=pf~-���ї�8��z\� O������
]ޛ�G�]�蝯=y>�fU�o�S�H�<tTl̒���J\_A6v�g�=s�v�?`�?W��sםA�W�U2���=]�-
����* ûs�ّ#J�p��:Y�xwVJ�u���v���]pV�%1�qF�C���� ==��H#�l��<��+4�uհQ��z�����BO9*U�E�Kk�lU3h�R�������]|�I~���+XGǻ?#7��|��_ݣiS�"���������H����hy���J�G�t�����٘�5^�K?�[���dd$�y^�B�7/�E��rR�Owc�/�"�g5�iw��d�7�Tח�6:�)���q�����2;��7�:,t�~=[�n����6͜{�Z}<qf���Nm�\�-�&tf�'��H� ��)�qٍ3��[ޯyz��mTޜ� Р�-��p��Za�Ϟ��A�B_�e��b�t}jz8�N�N���y-k�B�A�O����H�蕬K}t-�Z�PH3��#�s*vs��u����1:8) �����.6}>���,��;Ϧ��*��޴\�{��޹Ƽ�m�Iu�g�K�z{�5�+5vcs:���������ĹS y`_�I/r�}��8��]屓9c�!<?�1<�s�5}��R��0� ?!�ă��/+a��u������́�#i[�J��R���'�};�uX��C]H�b��!��E;��('��g��
��ky�koS�I+<�-��cd���#��5�G��Հ>=X��Tު�a�uT�g4�=�C�ڧ������ �VM�23H���Y�hi���?���sz6��x�>�PCf���x���cE��~�;L�۷��lU���� O�����=���Vnܦ�����L_��@ϔ���M|%�r���h����0�
��l�/�~H���ܝn;���n�!tF��'��ٰ�5����w>~fpy�Q����pBO"��h�w��*ޑvb?.k eݱ�RӭH�F>ix�%����j��O��7���'��W�;����v�=Q�gY�e������|�%$�G;u����b��5r�%F�ҭ��0�Nͬt�ϰ:������a"�Cl{UD����1����6���?7���1h��74<q���g�V,�p�Y��M��������Ϝ������=H�ⷵt��[�4�s�>4�=^��������'���Z���|٪!�IE+��{u��|ԡ(����}/����{��(*	t}�ڲD�̦k�'L�4�����Ѷ����أۋV��L��<g����Ǚ��&hAfq��k�͕y��k���Ɠ��E1��?=��|V�b���Ń���C.��۩�O��e��EqM�m�Bν�38
?8��H��-`���m����=s'D}��hЇ���H��驶���S��jD�A�QZ@��)�/����� �p)�*�v��|v��������s0��:��*r-^�i0�ty�$��3�H�	d��̶�*�;�+|��늠�؛�m�,�׷���T���/��\�@�����. ��Ӗ0��_*Qܡ��0��[�,�zG9y��%GÄm��]�T>�%�!r{��=��R
����0����'`O\�9x�߾|>�܋a�OP`�I�5oWB�Nב,���G���F�;�]�To�E�fl��m����;�n��2<��]M��ƣ�)�ҡa��~�A�d��dLM�S�2�A){�s"iV��Ce��w�L�6,:�֗-VG�ο<FE�Qۄ�\�����dg"`MǺ~Z+��_�Pu�q\��db.i a0[8)X豗�'�w�2T�_*��H�<suⳂ�N=a�4i��(��9�AV^�)�_"�
�ܚ��\���oc&T��x}\�@r�qB1Wzzq�lA�+�.u|3��dą)��e��=F�B�����"N�v�!�֧��Yxԗ�/Ëf���MH!Ⱦ�4��s��4Fz����|�1`��k5�W�vK�ӧ<�>ȑ��{ϛ4��y��Ez����{iJ�Y��:y9^^6��Þ����,7����N��/�� �-����л�Z�f��1b���cT�6��x1(#��a�_|6�,�:zĀ����M�yаε8��A��o�qŜ<�8�������p"}j���k]����u���<\�@�]�ϋ��v��8�����Y J��>��w
���P�A	�x���7�a�*�zD'���k�������u�Ȱ���$�Q�j�y��|&1�L��T\�@
ч��o^܇+	�_It�P����ݝ:�?d����a�x)q�l0��1�����O�ٵׅև=�"֦���%v/d�Y����ai�1:���[X�����P&F�[�'�
�B��\)˳�[
����N<��7��/����e�g�M|fg��&^ Vlk�S�^�j��t9:su
��Ϟ`!]�>r�]����c�ڞ�H��z�6K�<�3��I�d�\����3�`bb��8*R��yB�kqv�_�'��Oz��*�)a�@��]='�_�4�6ɻ����{���@]�)�u݂�<	�U'�Q��T	ѧ=���y�c�n�\�q��G:�y����Q[H2C��<���2�&��:h\<����:w2x��b��r^�6E���#{zY��ϟ�)�z5V�<s'�kH���~ ���hΌ�4�<�V��88_e�MLLL�1=��c����;2��޴�J�y��yq\�@:<���aǣ��x�(���R<��4111q7XK�B�/�@
�[��$���H\�]f�R��&V���@cJ��%�T|r�_�@B����m�cr��6����MLLLLD��^QPO��~LRxM<c��%g�s���/���֕=
5��l��]��@y�� �`�g��3�t�OLLLLLLLL\�����Q���A2@�s�{��í��}2>����[��9F��ʪ�����޲����������cD：u����/i m��)��J�;̥���kn�l��=�qpꎌ#}.�5#�[�͸,j	/@m;=V�Қ�����Xx�}�&&&&&&&����[�{���4���;l���N�6c�@����4*�YJ�s���������χ�0��07nt�A�qW���6浶T<���b>��ܤ��O	�<g�&&&&&&&*H3EWӠ_�@������$��=y�P�=1U�Y{�0ڨS��J�{s<LLLLLLLؠ]�.f!����h���3|\'D֑��6+T@o�=�!�3�j�9L�jbbbbbbbbb�x))�"q�g�w��I����#:���yVi��E4Í&&&&&&&&&&��KH�C]>�H��ul���Ŏ`m�P�NB�)�Q���@�L��J)�Ŧ'&&&&&&&&�(�N�x��w�s�q�?WI���$�fqĄ��݃��{���sibbbbbbbb�	��g�1�޸��ٞ�4� :T�a���x����I�.�/w��V-���:�2����YJ���&&&&&&&&&.k}>?s�2�M�Փ/i m �`U�'�[5萶|Q����9yǄ��[xW�g��]��W�����ĵT�!����������/�[�s���K��z����/k m��$��e֎����0��7ȪL�hbbbbbbbb��h�9h<yw�]��kH;�چe:��v�i��Lb�H��OLLLLLLLLL<"����M��l���zX]�n�M�!۰<�Nw,�ڑ�z�G�׉$�L�"�_�D��k�%411111111�l�si�����M��x����/i !LÂ���
{��O�@��S�b�;�I''��J_qNrbbbbbbbb����q��{����R��ƾ���S]2nZ;�1�	4;6l���#��7111111111т���7������3���z�~yS�ř������ⶉ�_�o��|�K�&_}�}n>111111111�P\�@��iT�q�M!0�Dt�)���r��R3K��kH���{�����������d�i4MLLLL�j;��(����ϊKH >lv���߶���d���po��nM�b�"�<	���%f f�V�I�4����5L#���xw�ۇH�#k�&&&��Q����da�1�"
M
F�d?1���Cd!�������H��|�u2�N��iM��Pټ�=���� a�)܎
M�'z�nbb�ʘ3��l�*V����NAW�/<I�ث���/�	�3��c�J�Qk��i����ܘ��軭@�i,ML�jLc�߯��@�u�⹁�AgNLL�6������ع�4���jt�wx��� <4u����sO�'�3�mu�{&�_��m�D�M�	bsj�S��V�Ia�z_^���������Qu���ʭ���$���4;�x�aH�=�P2�I�7@�,���}PN�+���3Ad�Vw�s��E-i��a��>�2�g���7�O��>S�}m��~_]\gJ_��jvS�X��H�6��;�&��ow3+4Cܓ1���c�!Ȁ9c�˔'
`�<��=Oo����KVRV&6�� �&y��la��,��>�z�]^��z���I�y��r�LX��� ��p����k<�z���_8<���4���6���-��3с��O�[X�.Cq^�-�"Z#��t��w���I�<���=]��ML��᷒^�H���y�|d��A����|=��I�4��VZ��0hN1R�dI�`�|0xC���-|g9�\���E^���<ǧ;?iX���t/�O;'9�_j	樹'���C��9�(7�b<������W�[�t���N\��¯9I����=�wd:(�.~�&.Vƀ���\�@��GA� �5�����y��-mM����=p?Q�	טM|.�!v�T�bn '+]P��!�;K�k�*��_�O�d<$��є�=s��J�,��r��s+mR�Q���91�)Аuy@��3UH�g�%��� 6��^�'�a>\g���I��=/���Q��#	������#kh{�`�Ӄ��:(�^C�Q&xZ�	���x]�9� -Q! 9��~�~��$�����z�ɮ�L17q��\^�,I=�X$-�GD��a���+����G

�\VqI�׭>����R1�2�;t�^<8!Q��l�N|V��t=�ilu��Y�q��[�]=�P�*��~�Y�JS��ݖ#+�����9�EQ�W{���l� ���X�M6,~9�<|�{�(.g �I�4��J��iY�#�F�̮���N�p4T��KzM��a�]X��_RFk�W���ȍ�>:{�t��QΓ�l6F� WB�x�+�}Y�E$z�_W�Kyd����k�V�ɯ �Fw�k��{N��Q�f�4eT
O��]�z}�-�	>�U���^?e�T%��I^~C���f�z���87��v����⹕���d���F\�~ur*FnR�Xi��+�q��8���|�|�ͧ�r҆m��v�Y�H��y&����S]}U�b�<s��۫��Uu��'�K��B��-"-T?���\�;q	�@p;B6�	!�����*�=u��U�Z4�epc���̓Q��_CR�!J�ݳ(�^���i }��۶ÜO��w��%D!�~g���Lޙ�Jů�	k�^~��m��|���qB���j^�F�/[֪"�ʤ��>ϯ��

�>#��a�ܫNՖpWF�>��\x��6_,�����[퓴΍{�h�9��@'K����e��Ō�����l�KR5o���!��$ ^�j�y�kx�F�^��D`��Q��Sad��s�l�=���U}���s����N��qd�%�a���W$������� ��Q���O���q
��&H6�{h���$����tX����^��}A����{�L�t�b���Xvn�#�h:ST0��'OȺ:|���4��z���y�V���8	w�`1 }}=��\��]PQ�<ْC�|�~��Bf��tP�s/���-�3����j�Ԩ�Xj�.�kR�b��LD�J�a���XP�&�̯g ��Ĥ�0�h�@6!�ԯ�}y�J�?F�h�	u�x�ԁ��6����բ�7��gUl�gRjIBv����n�e��	���e��U_O�f������/��L��wu^��������Ҹ*��ϧ��KHڈ��J��H+���m��g�^�ȹ�&�)�J�ы{
V[<����������-q/��;1ȻԞ��qe|q�G�o׿���������R*���*����q��e~/�ԦO�g��!/�Ό5ڞ����Tޞ{�W��Q���� ��q����I%�X�VP�f3E�⓪�M��ؚ�ꎡv�u�wIC�R����T�F;�~�]x�v��d�J�e����N6V^�@��yށ�ɕpM�@��w~���*�F�Y��܈FB��N�{m�����t���@2TY�d�x���D=��p.��=�#[(��|&���;�(C;<��~6�fSxP�v��K���L	^$�Y)��#I���Q�C�P�+�=7ft-]��7��6�V>c=hFL���L�a���ق��3 �Y*}�
�
֟���-%�GGR��N��F�1�?���Jr�,�TwS.(u-�B����6��߼Up�V��u�c��j�~�[ו�ͿA$s����Y(�hޓ!|�-�����V2�eIk1�ڕ��e��?��Y����7����|�&���5���L�*R�V(e�.ΕmD��d�/����5��^�Dh���w�3#j^�/�n/F�#�.���Ӷ"6<]Lՠ_:w�}�,��/$�S>7
���bW�.%c��s)��ێ��e�k
(��F��,ǧP`�b�RGk�*:\��+d�%�4(�ޠ9sxL��b�K�udZ���\`�FI��������1��{P&jd�S�~�3GlƱPo����w�mH���d��i�+�J*��˶dł�ۋ�4�ת!gY����u<�>2�g sW�6�����v*0�H#+c���g8a�z����N�{���GG��x�лG���X����=�_��kH�ʹ;c�r�J��L�ں����E��F���L,1$]��wx��m{=���;rD��ƽ���b6A��G���鍷;�dȐ�d,��'�����>�P��έ��I���c'T�e�NoP���Df6K���S�Nkawۦ���?�d�]�,�xq��F����p� ���{��j�����D��]����g�����W��6/�ʵh�5��'Ք�.��^�[sV����H~��Ϥ�s�ei/X��<0�\mۆ�Zˮ^�A�q�H���$i>D�Btp0�Ն �/�)}M[s�s&�{[V�H���#�ڶ8w��'��E����ء�����O���v#�UEa��T~�E=G�[��=HR����a{KWk
O���X:��;��w��!�棭@�4���A�y�{{��NV���f���� �Mg�a~��\������Q�����6�X�nc.�x��3�a�8)eMf�U_9Q�$%��a�-�H�b�>*�i��!Н4RI'���4���56!z��D�)�����ʩ!��#an3���j�KS!y�;�QY�.��^S.�v�c�"��$�ǝf#���D-{s�Z�*>�!��9Z��0x��s=^WF���I֦z��-�׉o ��uj1;o�Uֳ=$�������.;}#͊��@�ls��V��
=u�1~W��\_'(r��A���H���~�,w��X9�B����Y_h�O��0s�+g��X����Wp{y��u9��B�Mc Zr�+{��j8���~��+�W4	����᫚��gM�C巕���9:q��.���1U�	�v?X7<W0���������X�������$8N|��M��^�d��`��Y�|��5D�ڤ�e��w�ܘ��'4��������{��*2*#�8Ӻ�z���4��y���D�w`'��.FZ�f�P���3���i�h6<k�aB"�ݩTG=P�V�7y�<,�U����{�:��<��O2h���R���-��<���G�-��qM�]>�)-m�Y��Fۖ@��F�%|�SB-��n������*S��^r��ԸX��e������s��c�]ь9s͖��NSy�Y�!�=0Fķ��E"�n�&R9�"V��M��-g�����o�Q[�/�����H�:�`� P�tX8�s�7!қC�u�z�M�cz݊�$|7� [I�C}l��Ϙ�@ϒb�XU�EF���3o���:f���Xߨ[�٩�	��V�1�彚Q�G0X��W3_�d�����bKѦ�fuv��u��9m6��\�e�9��χkH�$�oх�Z�#��Ǽ� Ex(Q�M�G!��Qh�
�x�����j!���#�ӳR)uD)HU�r����4򵍦�1�+�`�:`[�DR��TW�S�P��~X� |\���,����L���~�nb��
E��q�HG<;���ۨ3	0꼜��t0�I=��{���,�)��IJe�B� ��;��ō
���M��y7¤Ē�LƑW���q瓕���U~o�	
�T�h�x�W��)`��5�H�Q�t^�C�t񲡌�h��;>󌢷D3�6�t�(�U���K���Rn�b�7�@�}�z�3�ދ���9�Y�W���a�hjڬ&ݓ��b��q[�|(8��O��u�bQ}O�|<��\o���aq���t���kH\�{�� ?3QM��O�v��F��,a�bЫ����ƕ�>	VN�w֡����wUX��I�QV�& ]C>sr�2G���}C�R#o0�ɒsC��Z�[b«��:��2�g����da����@��Zq�|<�߼ݪx��tT��R�l�6Lw�������Z�{���&	���5QL�V0��q�Ir����k����+�#�C��aXu_�hۮ[#4RV��U�e`@��~�6�Z�|��v���q��C8��ؐ%���\��杳9�J�CZ3��1�gs��l��]w@�� l��x���'�6ƍ����#k��ud���tM)�{�@RL�݂b����ϋw{�(g@�h��0���ij-��4�x����<��yw}�����Zf�"��m�y�D�
E�7�<��>���=��V��*E�:P�y��VԘ�'Y��7���W6o��^�n�M�ot��𽥕F[���Rw0o���6�=&��c���hR������X�EKQ�z�d]"�B��@���GeL��{�;N9������H�tX��e+:��ca$������Q�3�\�@����?ͦ��F�\#�R2Ċ�1�\��S��a��y�9zh}J�ap�|𺶓櫁�CZ=���&�g�s֘'��b���f�@QF��ʪ$��[׽-ـ���8cjO�7��ugh��´ێk��Q�ߴp�?�KD��.��?7�/�0�E�d.�rվ�g:�m��hH��P�1^��S�6�Q������ԞԮ��,
�㧛�)Y������֘j�d���
��f0��`�<л���hS9w���M�0�=g\'Z����0�x^�+adڇ�	VXU\��C��_�A�6���C�K�af/\%^���_Qt�n�B\h,�ߙo�RD�h+?�����
�~�{L�����]�9�<�<��^B:�C�/�t�=>��e$�����ő����������>��2L�4s��S[��vg�.'�
�@�JG�G-e��!�_�iJ�f�y[��pwM��f�9/��݆�7��O���d�Q��Gb�s�1bU�Z�Xƺ�u����0k�N6�JwK���y\{�Y"\�@JDI��n��UҒ���u� $	���.���"e*W,mϻ��TXZ�~��e�}���Σ>��mxRY�bz}�;ё�ޢ#aDe�fRj�Q1L^XǢD��%}�\)�9��TR�YV|���3��إv�J"𣏕v�$a�YS����1�TU�;�9]�kvhZ�����l�`[{���rt]b��x��B�J�Z8%�t�
���b��Q<�g� d���g�D?+7c��Pj���[��B��:��5�d��:���Z^S��o�u"�ǁ�ezg~{ڱ�PL ʗ�t9������l�2wn�K>��Q�:P����
�+S��ۢ��͛���oYIh��DO�l��l�d����e�e7�J�ֶn�:�_�Y��{j��k׬���q���	�T¨Z����5��Uf��mV�-� 2(�>Z9����üZ���ܭ�P+���퉏%�T����Ґrm�P*v��1p�^�d`!�>l��s��E/WQ�AC��s��6�|}���Z^^��(�������ѯn��at\�8Z�Z�^�|KMGNG�x����h�w��c��>�*c��o�c��N�[r���/#N���u$���]���X&�	�Qa��r��l&�-��v�7�k�r�ϡ�[������ܤ��Jl�[C�n�@���e�:)���v۳.S�m�D0~=�E��$����kN�5'�~;��><Q橁wV���-�;2u�Q�g#D�Rb�+�꛼E�c�іҤ��]�H�3}�<]g��i��-��F��~��h���a��Xқ�IWK���2�Zct����0�9�%T���b�=��F�/��˨�	���T��-�60c9��m97ZN���V��<-��w�E�on��m�da��m���>(����Q37P?�uٕY����!��Fɲ�:�w�Q]mc����7��e�:����>�N�#!vT4��4 d�	��m����R²���ް#� ip|�빚�<2���ᖐ�AR�2�r�҈���||O�\<�}�>�=\���gڇ�F�v�7����.�,�L�&B��2}���Sr�g�Db��;�]|�����㾵�4
,�㳃��g`l��Y�����}Nis)��PɊ;�rR`�)������{b�_Z�.�GƒӠ��IRQj������������5f� ��#�x�d(b�r����CJխ�!S
KԩU�n��}�Tjgݦ,�U�������cL��ݹ���aq"���.i �4e=� ��/ɛ-B�6�/�X	qh��2�9��
e�y�s6O��t��U{�3� 3���8����ՖN�A��=]զ7�<�,����hY%�� ˦�y᷋�I�XALpb|5�������0��=!|φ���<ϫP�S7�.����y�.���u��k�����2o+:r-��'|�Ӗ�ddv��Z���Q%��2a,�ߨ��nm)�� �\��}�gȖb�I*	�(�TJtvB�`y�<�H��Ǭ���n�� �g�j���>Dz*��0p+"x*:S8�`�J7�Qo.7�,��������R�et��h}A�f~��7������p��<��è����a�4�����+<�gk�%�������K�dv��t���S�7��'�P*�=#c������,G(��b�b��7����H��^ Y�8(�g���FhGW���*$oa��L�3��b��^f��o�>,0�m��U��KΚA>�|�����hm�|��!S��n��T���a��C}��	O�J�	�	π�U*����(�FTx����^�^�حV������@Fmx^i�FXa���y�@�;�O�;�p)c�>]�_���QQ|d%��tP�ӘE�1zjҢw�P�,�b�;)CD#�[Z7�������]8�Jڗ�Ǒhs�;�n8��7X�"��,���k�՗4���`$ᄀfv��`83g�1��	�?�[�w+����wծ�]ׁr(	��UC�k�V���*��-T��U�Su�e�g~���~�d`$��G)�gϾ�G��j߰�R>w+�J���V����*O��K�b~�xP٦j�8b���w��Vy�g���G�Z�_�Nt�������uQ� K�}!gnRa�Қׄd�Zр�f�,�Y�&��nAoƼ>"*C��:y����i�1'y�m�� ���	�i~G�z��
?��������)B��)���س��P�$�ꂾU��,W1��	��o0���H�	���/:?���g
�l�����+<e�2���<T^L���o��.pzQ�����'�dP�)����Py6PN4�nT��ց؋��= ����rz�t��sB�h�f��u����՝�����먬��$̰e	��Y�.�b��w���&��[ee�쭲��[i�r����!Ȣ?��4�
cRsI����q6��H.H�/�h�4q�cO���{w$�j �,��^�;�y�d�wq���H-�M(G�_茗���(qC��%l�>X��΃b������(m�����B�����������w�
]P���$z�rWeF[��C���Wm���R�<>��Z��k��EY9	b/j���]��l�,��'17�s���E�m/O��מo�Ђ�ů���v(z�e���Ђd��e���-l��
��fF^aQ�(��U��fqi��ŕ�GC�c�(����%���>�:�ذB��<�����8~L�8>�o�C��4mEOR�[<k(D�����e����@��W�S��Dz-���l����:�>%���,ԗH���DdYYu�5���bM�H\�@��,�\���:(��v8К�����k\��R��W�t߷��.�w(��()�I�B�N[
�G��G��LՋ�)k�O�Zq����gd1��D�!`�M{A%h⥡�t��#�7j�_�{�W���@dIe��C�:_`�"{#Cx��~d���}�i %�#G�y�U�C���aL�T8e;�A�m�a���&r�E8������S�}���6p0_���%-Z`,h�yj�Kw�0�'A�jukܰ.��߼���y��mm�M��JF�1��A�-Y��P�e�[/�}f����r҇����/I(.�� ��tH�����]��><����B��"/I��؎�R^���Y25��#B��Q�����`$v���%pIi�nٵ��+������2X*g��!/LL��I�g�Hh�.N,���x�P�š�}e���؇#FR���9��D'=]#������X��z������V�����c����U��
`��PM'��U��ߑ�g�ى�<����a�k�}�KH{è�3��ռ�������qՖTN6=Lڜ'�����b���8ȭ�׿>�v^�z��f���#�a7��IS�Hn��� =c��ς��Z�����=�q'�4���Xf��'��БZ���t���5g�:���0�B��_�o�����~�����B-`:��O�KHP�U�yI��=yG;0��O��@^	�9w�-�L�(<�sTDK��w~� @�o�rW�5#Lb�&$Xd"f$�8aC):u�n���?�J�2#�h۽mԂ�>0>�؅z��|}jK6��X�Q����;*SwUjN������q��׃0��"�(�{���t�+|�#1ޤ��JE��@_9���>jLc9w+o0_����-e������Y���Z�z4����I��Ռ$A\H�f5�gU�T|%\�@j/�M�zލ����̨PكQ>ފ��Ť���U�۵˩)�`I�F<d!��\�=��2P��a��9�:7�1����<�J[u�����;���_A���Ե�CS���9�g���}��س����ſ����k�#�ﺃ�9�xG����b{�����.Ry�|��9:�D�P�O�%$D1��_��)$��t3n޽��h���a���3�fŵ��3��n۬<�ȶ��Mи�:��v���ο�1����ҵ�<+��THx-AS$!�����3h�Q�޺cw+ZǙ�"�������O�<�כ%��bx����^�6��y���O^�|�0�/�����?��m��W9�����[`2��~�O]�N��B���"���(m誁<
/�Yz�$V��W����YC���|���A��eO��}uFh;'@TśL[o�1��b�m���c�w^EzX�:F�;ۀB�/�coG޹�u:`�bw&x[I��%�]\,��?�2��������[�ts��C!v5liVv�M-�n7���G�d�"�Z��T�|`�����٤^^&/�J	�w�)���y��ݹ.�B�y����Y�����q^)<���5U1��R�܊[u���zӋH��O@V�Pq_CS↷ițS)���B�ὣ4#�LT����!f{�qzf#Eq+:�
�S�崂���Y���}-?���g�F����)����u�k�H�pJ@R��]]�qJ5޾��R��Y1�l˪�rF���P����3g�r5��dкG^��2�I��{�s��=Jw������:!����ԋ�!��ߜ<�E��8݉��k4�M����ϑl.t�J�G�I�]al���φ��L�oJ\t^1���3���32����O�$z�J��-�Q�F+/LFgLPB�.v�h�Y�YYJT��kT$^��yV9�s�i'h�����L+'|6�Jcw$^<
�ȇD�ڑur�k+�c d���ͬ��_���B���X�K���)P���s�.�-�v�����Ry����V�ɔ����Q�l��`��/��6C�5�J����#s2��0��En��<��C#M-_A'��urd ��
8k�-o���S��������Z���b0�VeO�������ӿ~.,���W������g8�_���{�������r��?�g�3�O����տ�+wU���;���k}$-h�?�=���S�Z��?�&�������i�{���_s/�_�����甬���o��}F���W�/��ݽ
����ι1�&��?�~�~�[�r���w�&]�����������N�����o��s��,�����O�k��?�܏����k�zҧ�3��C�|}bbbbbbb��`H�Զ_��&&&&&&&&�
���h��Az9��b311111111q���p�وW����s���ך��������8�@��0 �ꖿ��Ο� qbbbbbbbb�50�G������8z���u���������������4��i]����Ϲ�q41111111�1��	���8���j��OLLLLLLLLhL��SH����C�����!������������������~����O���������ĵ1��;�sHW¯�8n�}��6��'��&&&&&&&&&��i =s�2��_��~�!E���̹�7711111111qmL�р9t	��ᜣG ~�݇��nbbbbbbbb���ң1'���_�c���?|HQ�����?5�}bbbbbbb�E0�c�=���#���=��m�h���;�y41111111�*�ң1-����C���?xHQ�ݯ9�������������ċaH_۬�6{����S���︉����������4�&>=�?����=��u���7�MLLLLLLLL�&��4�����;��_<�������o��MLLLLLLLL�.���h���Q���/RֺF?�[yOLLLLLLL�:���h�\�o���3�����1���o9��?�&&&&&&&&&^�@z8��]�a����:���)~�w��nbbbbbbbb�s`H�����?��~xHy��~��w��&&&&&&&&&>��4�9��Çq�{ο?�8�� X���������NLLLLLL<�@z06��Av�����m&���O����׿�{�o���u��U��������~���G�o�i�~�c7q.�ҟ���7��?���_�������MLLLLLLL<�@�B����o��_��/�����o�/�����r�_���������o�����������Z1+��>��yX�^/�����0�����8�w~��{�/��/�Y���������*o�{�;!$!���Л(E�"��}����^VaW]׶�]A��{GZ���PCi$��~s&�	JI�{�����<��ܹ�7����?eee ""s��u�N��H�@Bd�� �A�V�տ�����х�����#�Ꮎ�0}��K=���F����Z�����UJ8�����Ѫ�?n��n�!p2輺;7��3.�.��4ֹec4�:��r�u �zsG��*�z�'��0 ٛ�~77'�����Q�lTM����D�M�~ݎ�'�pT��,�|�Vgu����_-���m��~]i���w�m��)�X���J@�!������ہ�<�l�NTWl�ٝ}z��6�_' 4�<%�#�ѽ=���=���e(�G�TBQU`,NΠ����#��y]�9�)�����>U�����tZ6�H���M���84�5OA�n�Cоy �X�3�B���I�OH�f������U���O��5*��i��Mv���v��^���
k#��=ʡ�.��k�e�*u�u٣�Ƈb��HM7�4V�4?�>:�{��f����0�gol����w"d\��<���D��h3�ps�����/1�~؊���^I��͆�(�E0�6$	�~��m���x�ɑ�~�|����j;����k@�d�ּ�������f'��[�w���1yAG��|0�)�n�ؼ!FrMB����|��]u �pa��h���� :;�.&�>��;�Y�SW�GE�����	�}��r���2��v��.��\��{�jr^����ϑ��pT�z]��fX�(tV�!G��A�����_�Ƣ�	�3�k���@�^��O�fP7 ��]�}��O+u�G�HO�N̑s\
Z6���j���?[��[��\VOX�Ѩ~�u���H�lG%F�&��	�}�+�N��I�b?68���LDe����56D]�:-�OMz㵱�G%~'��/~��3�5rK�Ād`�A�x���j�7G���&�߭��%��t�*O�s����߹:;�%%(N^�߭�_x'm9;Y�uc��n��٬B�=�꘎��C�h~K��؆����ql�3��m���O۱ ��db@2(����7������)ה�������G�W��󙫼|��;ڡ���N�./ �o�{]D�*�m(��<{��x�Q�j�sh�h$E�٩�YbY'�K�߆$�)TM|OOFX�>[�D�0 P�ІxqT{x���w)��&�����Z[�������kz�QJ xeLG�����3%��`�N�<"ĿpS{S�N�)�;�ѽ=1�T��k�
�tu�JXk�\�Y%�R��j�Ӆe��'�la�����NGW1f@{��۹����U�)���q�}kE\���wF/N��;7C����f�>���KœÒ�Q*~G_���^�_.�nCc���[:��������X�U�LD��V���*7�nMa#�����r�hݥ��Ĕ:1�����u���pw�X�V�g�Άv����'��)��}�ڻZ4��?flQ�Gm�I���x��Qh䉡IJH����,2B���P�pwuƛcS�𽖞���Δ`�Ό���� P	G�,��e݈���9Eذ?d{���t�.-�kY_��	�e,nk���q��1����vx�U؟Hꖬ  ��IDATY "{a@2 ы�̈d4�T��{%=O<���8z2O�������'��x]֍��~aT;<��>�mL#���:�VG4���C��ΤW�tBP>{jK|v���	&�D^Q)��� �R�=�4Ս��^{�<2ir]}��-��i��-y]փ��+�6&*�1]���ǐd[�3).�ŀ�*�����'�Z��r��'�c@ҹ��qs�P��5����_�X��*�Y�/����T?|��N��u*#�C��3I�xjx^��D�ƀ�c�2���Aڈ�Ĩn�YA��Dyd�wiC<��(ץ�(Fڈ�W��8�"C��������C*H��ᖞ���J�P��?�%;��Ȗ�tJ<؟��-<��#��m}Z`�ޓ8p��>�J���zr�����n�����H�~���q)ps��u�?9��9���0�~<\]��87���#7�ck�i�>S"[a�[��t�A�p�W֚�K�����J�Wr�]m��̓A�"O�H�_>\��rNo�+�����mY%����Gs�q������ZA"m��'�%ᩯ׃�V�tH�P�Hن��v{�V�xa���u9��m�x��w~���'�&�E���3^��M^�R�G�ё4�c�6:��v?m� �-0 ���-8$oc7v��̵�S��a5uS�f��ic�ۆ�k�x]֞�V�'���G���n��uG�vk����ze,pC�ckG��
�e���|�۞X�p�� �`�N�Չ�_bȶ�u)*^q�v"}qG_VUԚX��t�q���׆�[*9�ȶ|<0�K3^"�`@ҙ	�q
����֥�xn���T��N�f��G��y]����������A�l�Up�fM�{-���2�{s��!�%� ���$G��j�>Do���-8��*���-�	�>DC��kb��M�����o�ND������L��Puĝ����U��5Ť5$��KȾ�I�gK��T~1��F�D��G�D*SV�27'u��l��-0w�d�>yU7v���ޮo����cA��V+��5H�>�ڊ������a����t�~�jc��K\�#R���*Fvi��p�m� �Р8<��F��Y �ø=���y��b(+ڑ��$���s�Gv�7}���O�7\i���:�ߵIa�t�nsn���=���I�!�ي ������{4�1\iC��)C�&����{��p�u�� 9��ti⺼A	�$�(�~C�(Vh��:D����~D `@�41��h�#�$w���Li�I���|�>�M��P�G�?Àt��1A��$O��0�K��c�����D A�Hv!�b}�r�d��%i�I��G�����bC"��7��fi���$pM�l�1*��9��b�&1��G�  6@e��?�
�KT��rw��RN���c@������Ar��6M�[�x�tj�$�a�r҅n��CT��t�d���y1!~jg������skɎc �/$�z�6V~��^�)?�j=����RD�4����h�Ƅ4 �!�7�����	�և�G�!f>0 ��$���^p�����sz�^p����zA��w\S|8o'+���=�������H+HRT?U�,4�z!���G4r��$��V�� �hސI���ĵ: ���~vɅ���tU;�H�4��M�Ym��I�����%�I?��0�a82^����ZJ�`4�v��-6�I��H�T"�HR�HT_HRT� %�8��$E�g��Rx]VKV��bZ�����xM�O����6�~�d�V�6%G�ƪ7!��je���8��� ����R�y�]9,��Q��ڸj��&]\]��=�,vak�)�THX-Vu�]�&�ĤG�ʃߑRT��鑸_8r@��tE�Ƽg�I�A�D�?:��n���d���[���ř����$
��F�z����p����{����z.�З6�1�K��tv��E�����p,�o��D�À$���t�덕j.<�q7��rs�u�Sb��#��<�/1M�7z�G~^�-f����<	#qqq��;�qǾ_R�1 I n���W���t�-A�"7�-�1�Gb���J�sϙ �VT��2�(����	AHTOl�`Q��%6��<��ǃ��r�������^~�Z���۾��C�`��m0�� 9#�ܛ�ꋭ!���>5r�}V\]x]ꕗ��v�x�9+���?1��6 �9��w�����kVVV�(���$ow�/�~�$qseCT�\�!�l�u�W��y���zP�E;n�Kw7��/�Z���f8�����!M�JymwW�ҡ�a@��ՙQ�%B6��́G��<�����㎸;K�aFFE& ��GH)� �:����V���#7D���X�?r爻n�x:n3B�����? 7'zעU����;�/ǽ�I&�����D�2���������G����F�e��ym��δ�-�a�:�Yp�����WI�ۓ�[�^A��WVI{m'�ϣ�ptM���yN�����S��M֚Mggǝn[S���*��/C�#p��~�������&�]��CQ�c��'�0 IRYe���..������������u�����&)�xxx�(d�9�;M��O�:t��EPQ�� ���,m���J�AT�{g�I�FUVy��M������7�������D@�U�Ǚ3g�g���9�;KZp�i��9�4��\]��R�s����IHݼ	zШ��5��m��D����I��ry�7% �u/��T��Rǽ��ټ��\P�)�q�]_ϑ����Qe��Q�;����Em**��/E9~��NfBD��C��Ѓ�J��E�Ā$�Ŋ2�����^T��9}z#v�VR�7��J}��aa8t� �JLS����_�I�虯��z��Z��{q%��	H�<�YR.�Yѩs�X��R�����#}j�y��'m0 I`�ZpV�(EhX�.��M�.�Up��H'�gA��Ցβ2}�������/���ա$��#��I�qA�:�yd�@����]{�ĲE�PRR,�{�_ǔ.��rމ\�}��6�����X����H�ڱ]W����U�l�v8����T?�[�j��۷B�ZĶ��k�.���9�),"R��qH��ɩ���S�s
K���v� �_�����D5�.�{¿aC�ɩ|9a�̃I�S/�{8;ə[/����t�#wK	��Kq�t��B����M���7����QZ��F�yQ��0�$3�q�U�ƅ��c��m()��^L�V�^���q�����Sܺ�聭�7�mz���L��^^��Vw��9��'m0 I`Au(:����H�>Z�n���(����GM��BN:�м��"�"օ�:���ب�]]]���$嵏8�Rq��Q
�Yll�8�U;O��
������J*������,Hj�^����k���UĽ�y��j��^�
;z�q$)�{Cg�����x�X1�idKj�z!~.��ȩ"]$A���8t���1�)�m;ie�y���FxT31ھ_�B�?� !���� �H�:�2����~y�(r#�#�3�g�.j�La(�yZ�����7�..+G�}�< �a@�h��t�m"�{S3�=���\i�C�����,�1�e^�,���O��b�u蔂E��\�Hg��P�GDJym�f�d��l柕���u|���CO�����"�8��]8�Y���t��_�#��qu���'��X����������UzV��i�dHmMϑ�-��g:u銥��\BŰ��FHL��z����pt[��3p��@���z�2i�ƋM8e��5#V~ދ�$sͦ � ��6G22���r���ڟ��Q5�JU����ág�:�8������ܜ��Q��K�����NK���xF�y��R~ۗ��b@��\Cg�Q��TQ	7�sx�ˮ�{`�e��~U��N���u���� ��v���|���~z
E���d�ʋ���G�>R��󺔿fSHn���yҧک[���k�d�±��T��Z�d��kJ���G�a^[y�$0 I$�Ѯ#yH����߅DOQ��=�v�*TT�~*�ht���z�8��a�=���$�=z��*1�d��vb�H����}���d����0{�����QxF�Z��je�t1-9�L��OI��=��'�;��ш��we@��c@����\� �C@�w�~j�0[�Is��ڶS7����(3���	b�BoI��>�\���u/��L�]�Nҫ4�����z�&��^}�a���4%{A=�kw�^=��6UҌfk�i$��u$WID�ŀ$������;N�>����#_�V���Eڮ���ԋ9��m�#8$z�z�	P���O���q��15��u���s����������OJV�𺬦��q"�t��[	�춉��r]v��C�i��?�IX�v7vn�o��n�K�ŀ$��#H�gX,r�[���@�Xޱm�Z*�>Ğ	bϥ�b�g�U;�[����et�RZ�ū�Ɋ������~S}��"J9_T��:KwU���x�cm���nb��];�۴�Hhx����Ug���A�ET�
K�)㎦��
����t`~�Q��W@D����R�`s��1��<���5{ �ƃجNlb�-ww}?8DHeo���o=��$xxx�M|�z�k4#��2Oָ؈��CC�լ���HoĦ�iG����6n��<t�	���m
�""��s'د��T���$u��ޜ-�����ՓIT�\��G�$�m�I�9��8��,�~�\���N�#�p�ς���塰��������������F"B*]l�������^�$�0�C(..FQa!Ξ-B�z�Ea1����K�{z,H=����H�/�[@����u�1-Zb��4=r�^��z��6m�N&�Z�7K�jb�\��'1 ��u����sm΅���Յ��:��U+K�s��U`uZ&z��g�ؚ�����r��E~ܘ�[z��mh���v舄�8z8�'N�����1'F���ս�D�׻ջ���Bb��c��5׳�(����+"�0 ��̵���h~��������+�)�Ň��Y�Š߉Τ�CٺE��Xw)�m�C#��e��:���rX�U��
W7W�8�订�ՔWVb�>��0�kṛ�d�����Ā$��1���fjz���?��5fSQY�)���.m��<l<����وiu_-�uy)Kv�0��(F��=�� �Ub]lE�	�.D����Miy%f�g@"m1 I`�̚����UR���ܕ�c9E���v�0 �ך='��m�y2*�6��Am��f�Q3���k=.Et�M]u OK��/�2PXl����q0 �p��$F�DŪ�a���K?m��U�̈����ѣ+k��l�xY��)�K[��(�vo�Q$;�GӔPJ�5$).��㋥{1q|
����<�^��tI޻�;������uy߭>�����l�
�f2c�Au��.M|6_-ߋgol�����3\CL�c@��
u{7��R��O�NqY9>Z�T3;��q]�g�Еe��c�$�¢�e����ѕ-�v��E 9:d;���5���0 Iq�`�S�=Z7��;<��ْ��͕jN\�)-��[�{��x]��������h?�KW�4�ս��v||_/��p��VDg��rKdl�Kq������=x`@H{{��a6+�Ԛ�.��0��m�Hv!f��\���s,��(�l~ژ���<s�A��=�=��="[b@ҩ�k⚄��t���i*���ڛ��0$�!)������PV�����]��� 8;q��>_����ji�}��O�v�(��sv�Ȗ�d�����7c�=���r�Z�`�N.���W�߄/���RC_.݃��A��q��l����Q ��s,�n>��W�+�7�ݻ��������'9�l�I�^d�Ť��1@�'�����ONa)�K���B�z�|�^to��Ͳ����������u�[	����y��bAb&��1 IQ�ͪ��<f��Q?"lN���^���=S�WglA���Ϻ�+*ŗK����� ��=��@u':�"� Ou�~�@="�$)j7_���;۴!�"���^�����5���D8�-�����th�����2�`�ߤ��":��ޠ�[ ���f��j�	���-~�����_���ZK�g~���u$�=q]�}{WD7����� 5=�� �i� !�@�W^Y��flV�WR�����^�>�xq���(��T�5��5�D�$E�+.������G�wa!76�q]>9e>�K�y�j�E�y]jL4@_�~�kd��4�ر�"<3e=�u[�sXC�����7c��S �'��J`�uYq��k�52,�`{�J��޻�;����7+Y��� ^����F�5�����8�\����ՈN�ջ���[32�c=����ˣ��ǃe�/gֺC���C'Ϩ!鍱)�.�`��ü.mL4�ž3, R7���㭟��lG���<}^��#��>^�ƠN�0 IP�zU����1q\
�p��b`��ɛ�;�ץx�s�ܟ}�l�X�d{�ۅ�@t�	�\Na	^�����@�����5xeLGv*��()��O�0��I"$4��==�<����@^(��R�/�y$��.�d5��	�B�A|�� �-�2}3޹�bB������b��%�G������r�>c3����LHv*�X���0�:4w�R�@���6��K�K��k�܍m�-6�L\�����^���r<��z�s|g4�]�(���W�Y%L��/�j��a��e�h�<=u�:e�H6$4�R��<�4n����ig'��f{�i��Y�͕�AL�ya��Hi�{��uȪb{��)��F^����/��ͱ)h�؍��%����A�^I�l����R��V�eb��8S²�H& ��L]�;��๑��������z?>[�[��D�"~>�b��._��8��4����AEUH.1�������-ЮY�w"���F���������֌<68~�����x�/܍k�HO���Mc^L/��x��x�l�f�]P�I��a�N]�;Qy�^�|`@<�M����򝟷c�ޓ �()���S��7�C��&���}�A��$�khw��S��"9���Hv!�1s�p��t�I
�M��),�K�mRn��x��D���CIY�]u ��d�%)(.�?l���ø@��΋!3���+���)�3z�ۍխ�ү�CNG>o��\5������b��]����pm�����(�����uS**9�N�Ā$���Ѥ�?Z���0�WKx����]����]�|m2&q]N��J��;�ie�i$⺜�`7����o���� ������Ֆ�a��4uj�۲Ǳvon���to7c7�Du�9��Eij�������H�̈����G�MoL����񂒘F��=�7	��qC:�8�뒤�|0��o��0����ퟷs�#�S��U7�ӭ9n�	wWc���;O��{�iuDF��$���	�E�_*7&�`�HR��ޔ��� 5�����#qS������>��9d����v��#�'��68�������|0o'��>`��$�'-�vSW�g0"�a@r 6H�%��R��6�,(*�������c8p� d~��v�~��-�$���v��.�˰t�q��|���d~T�;1��oC 3��;m;2��AI�3����I����Z��,���zL�ŀ$����A:{�!��� �A�/!�~rʃ�WT`���X�~7~۞�R_����%��w�e�ec�z��R�k� "i�rye%�����mG���,��01�A��t���༣wK�/��X�����s�|D��oV�S�M�:q��������GPZ�+��喃��:"#c@rpG�1y�.|�0���H�j��сH�
��z�6joF��9��{�c���(��!�����始w�%�論�MV��D�h�m�����D>R�O����8��n�L�c���X�4�����-�u�Uiy��� �a��r��竇-lѤ�r�T�	���f���"���U�9��2����FdHX�V�e ��#���c��C꿉R�э}���x#��w�*�=��cY��Q��Hf���8���>�EtB��}q��P��.#�0�\�굩|�պ��9E8z��N�h�Y>U�=���H)�yC�*A�m8�o����yEe����Y�190��#��ǴU����G��kX��k��7kSO���{��8��;+�},���L�I
c쿱?3_=�H����g��	�.8�Ú{J�A�FeE**�v��#]Ε��sצӹ�Ս��_�uYũrtub4F�rqĄ�aP�H�K���~
܈��9�c�֣ ����\���d���qq�t�.�P�<��lbq��M�SD��I
c7�����h?̒8j�si쏇$9� >�I[�3�_��ù;ѶY z�A�V�����S��&��w����p���ET7����q��]�I+L�����Ƅ��U߰?K=����N-��&�-����]�G�(G���)��V�o��ȶ��0����Ƅ����s=�EZ�6@d�}=��|�T�^��MnQ)�J*PXR��J �wB���~�+��iD˄ĈDD�s8��z��1 �`������8Ŏ����$a@���@��g� IDDDD���D��'��}LHDDDD$�fl�k8*�}�����H$�!S�A$""""`@"�����$� G}�������H������L�IS!0�"""""GĀD��p�� �&m�>HDDDDdH2p������H��$�r��,V�!�HR�pIӷ�xDDDDDr0 �`�:�V�>""""r8H�-C����$�	��Śp�������I�	��S�L�������d0a>�4Ԙ��!""""C`@��Ȧ��֮e���Vo?���RYK��&��z� �� ")+����&�����ڜ���~��$R��M=������<��������a@"""""":��������$"""""�s��������a@"""""":��������$"""""�s��������a@"""""":����C�ǿ��\V
KAN�_���xx�T�*a����TVO����HY�r���TV7w�/ DD$����6��),.����5�-%Ű��=T�Ƅ�/L��NYG59����% ")9��S������ �Y0 Ia��X�<�	?""""2$���	]�j�i�����H$,&� ��|DDDD��HG�D~4a�$""""`@�@D	� -G�8EDDDD�0 �`�t�1~>DDDD$	�fL Z����!""""#`@��sȈ�����I
��p �����L�I
� Y9*FDDDD�ǀ$�ՄC$Z�#f-""""��I��#mY��H2�p��b�p�X3$���D��tDDDDD�0 �1!�H2��ODDDD�KH�C&\�EDDDD���$�\���$H20 \�����H$)���������da@��C$W">f$""""��I���� ]$���$�Y�F�������1 ��4J6`#""""I�d0�����#Hf������H��$0k�_�/���1 ��q������H$�:���F�bGDDDD�0 �v��╈�����I
�"""""=b@��b��3"q ������I�9S��ለ�������ŉ������H$L���>HDDDDdtHDDDDDD�0 ��&d#""""�c@����дyc�'�����da@���	@��e1m�$""""�c@�¤@��e����$�Y�I�9$	�Vs	s�+""""r$H2X�:��~>DDDD$iF��b������H$� 4�c'Nc֏������I� �B"""""cc@"�1gx$""""#`@��-W��DDDDDr0 �`���E��g�χ����t���c�*�p�������`@�C$�r�9?""""�?$Ҍ����1 Ձ���A�����Ȅ����$1	�!�6̻O�R�o��)$����U;�~@DDDTG�Q���� ٟ���(��\V��Jq��wEye�U�;�z��mX����<�7z'E���Z��r�_��c@"�� I��Z̷�Z� �������A���[�����z���_/�s���%�u��gK�Qt���Ҳ�����V����b���C�r���GQI���j�I+��jZ�sȮ��H�|�=���͚���(��7�y�aGK^��X��mv�Y�g*�)+���C�� u�T�����IC��t��c�"Z�kҏ��H<=�΅� 4Fs%�@�\�{@E���ѡe�?��J�+�#=�N"�`&R�gb��lTV�&DD����V��$��9��|WD�������+G���m�H����1ᮼ��-���yť�خ��LlQ��Jx��4C�1�O"�!��h
��]�A"���F~蒬�����������<�]ѩU�z�WRV�M�N`��,N=�-�O���̋�,WF2k���}�����ɂ�1MлM(�&F�}\4\��@W���nq���̘��/*��m�X���o<���"�y0 �J�v�5(�r�#}hD�մ�/��o���#>��-����g8�K+��gcI�!,ߞ�U;��k���ȸ�lH��tU;���h�kL��ى(�=�k,Ftk�N�����ZG��C:��h��#J`JWC�(�@DD�dC��ҡ�j�֊Y���5���P%W��q�pb*�B~��9g:c��]�f�v���-]�}�"D�����έ0�[+u�������A��cۡ�����J`�-,��'s7#�L1��,Ņ@e�&�zz��D�.���#!Zc@"�8ڒ+"Y���k�0�o"�y��/1�1�j�Wo냹��ai��t�'����ل�'rA��t:(+��\U�n���]����#8���v��׀1�㺶��-�����3�v�U�9g0m�|�p+��* ��M]�c�2�&}[D2�"1R$F����G� _��s��������M8���n""��l��zx٥M��� ?<0�#�^�/wW�y��i��w�o������f��H�r��u0op�Q���*KQ������v�Q�mO�Ai���(����MX�8�b�v��GTwb]�#J0���f���Gn�K�{�㹛��-8S��i""�2$�p�^_G}�Du���{���C:���QH�����~�_-܊�
mJ�ѥ1 i�z����b�&���|DTc)��xq\o��Y�.@��|�-UG?Μ-��Z\����׳��VX����K��}�|=����~鯗�7Q��eX#�M��&��O]���oWb�4TY9jODdH��f"�,5�F���G]v�ٹ�O�EȄ�7�+��VKv����<TBЁ�8����9r�D�ͮ����u��1,�͚4Ds�_�C��l���@�z������K�|[:�H[�Π�9��Ƞ��u��|k��VTJ[�T.���l���-�&m�3�]��*��ȮwM"\��`$Ǖt��)<���ףY�w:�*wO  z#F�ıb{Ɵ�"d���,D�'�P�S�^�BLɜ��(5 �2uRd���������$�+?�Ǝ�r��c@��s����9��e�K�lE"�%��	M���1n����X�[��W�u;�_X�Q�:���˶����'vd��>��H��_���^�QX�3V���߮T�Տ1���x����v�ū��Ah�/����k������T	Fi��Q�ܞ�/OY�����6Z�0�G	M��z5�G��~ހ�߭Bi99��V�6��|[�Gd`-B�{�C��p����L5-Q����ԐD�.8���w�� Jo���7)Z�?[1uS��ҹ��|5�Q�1 Ia�)vD����O�l��uFb���+v�����k�v������u��r��n��+^w��C�1���j���X���"Q�1 �`ڑ�����A�'�4�_�A���Qb��5{0]	Fkv��ǒ��_|3�~�p�z��aL�%,�Q���ō�[��v���7+���T�'"�!$���2m�#�������ҥ�d���԰�kv�l�ȩ�����ѡeS%(�ax��h��!�[SG�&�}-��MĄ���I�u""�c@�¤	I˷ee�"����=|�Z�[D���P$������o�������1�S�Q���)-e[���5��O����&]��l��L��F�+�H��]]��^��N��_��0u�v|�l���ǜ�������vm�ۮMBR���ӛw^�Acp�{sp"�������`��U�#"�jߢ)>|h��MEŴ��~\�O�m�[^Q���W��&KQ���3!�߹�O^�Y��@DDc@�c#Z�+�9?"28QB��q��~���ƿX�i�v��G�G��@<:"�z�I�>�ڹ��k�7S��B������1 I`�դ$�s~@dPb���������vH��^�ײ��b	���W�:u�	�I����ݿ�:��]o���3ADDH�%MG}��HĆ�>t=���������ά�X�� �|��>�g>[��߭ƽ׷���!��Ӯ߃�7i����>��7p "�ǀ$�i>f}_��4��Ft�ӣ�����s>�mM��J0Z�����:���W�S��θpGx�����섗o��I����_p��DD�����uCd2�ԉJt����y�xΖ���oW���xvLw��'����')��_����y "rDH2�5HX���O,���썈n`��=S\�I���ß7�HL�{����߯�0��k�j�׎j쯆�[��֥��a@����M�.���C"]��O�:~^�v}��+v��/�";�,�.�==�����c����hn����<�Ë�����;VL$"ÀD�nI��2�@�����x���v]o��H6�p6�;�+��a�z�"O��f�Bn.����A�n�I�W���Q0 Ia��ە�#�Q�����]����E��Ǵ��d�fՆ�ff�܅7�ꇑ=���5E ��c����*�>���.��$�9��Ί�C�lO����2oHii�ל�d^�jrK@T����f�ٍw�� o���ؾ�h��y�g�-��1 Ia�ƿ9s�����>=�[����v�g���'iEL�[��޼�F����뉪�s_��^�^-"ADdVH�-s�I3$�C`/�za4�"���zb��D�� �5�{�W�\���h�Ѥ��@,xc���g��Ȍ�H;A"�h�kcѬIC��֩�"��֏,�L6�h�A�<�	�q�5�;ަ��$���:#_����O���l�HCZ&$!��������GK�R׉�.(�=�Ѥޟ����}<�l�Z�����cp�3�j75&"sa@���m+kϑ��P$I��ʔ�xw�z����=�z S��6��F�����	*�l��4��LDv%��5Gbz�-�>��~`!�.#+=��9޺�:�~]��^�ݵ�dC_|:o��̀I��D�;ҡ����T ?/w��΂M�)u,�Lz���6�(ޙ�_��/S^a�Z,�����d��tI�PcaB��k��^m�p��g�1y�&�ь���b
S���N؂�ł���e�(""#c@����G�X4~���Ȏ"�`���x��5g�S��GDzv�D.�<���f�[\�M^���	�?>�^��U;Y�����I�IG��BQ]5n�^�~��{�c���sJFIY����Z�	6ywWu�a/�-,NDŀ$���#W�)vTG"��#1�d+s7�ø�?�Ȉ�p.v��k�����Ey����1n&KDFĀD��t�՞�N'��YS�l�����}��%$���O�����%�zb�s�p��_!3�DDFD��F���)vT;n.���(���7��¿f��,ߖ�k��3�ߛ�@_��ࣆ���o "2
$"2��>|=��������߯�"3�w�4�>�%~zyZ�j~������p���L��W����HCZ�YYȎj�Q�0�s+��[4�n�4��iC���FE�3Q�R��vr���|�Pe�VU��J9�(��BIY9*�x���������j��-�j~�	����p�?g����H���jJ�'��d��%��t��Վؠ7*�Q��Ղ�W�V�MK��~2Yy�8����|�g�aW�)���j&��C_��o��=�@���SZ�q��ʔ� "�;$)���*.A���R������g�*\���6]����5k�ظ��T����C!1dA���ѱ՟G>����H6��R��V�,�f�4Q|���᳿��.�����a)�<�,�""=c@��j�ֿ��;1C�U4��ĴgG�ӵ�&Ѣ�(�t���0�Mi�>ʑ��\Iz�'q�qDD��^�zK��GPVQ	�ݝo����_��}5?����W;�mM�^���fb\_S�cGW��섯�������u�x��-r�� oOw���J(R�Ȧ�/�71�%��tT�0�H?��JPZ����#LPKً��k�I�w���u�LQD�iƪD?s���޼yW?tn��y�~-C^�������	ɭ#�@Իc,:�7S�)���
��,D=���g�p���x@e:[ZG��G����;�hz^?/wu�%�FIo��K0i� ���S���-��$����q��.��q�rhM,R��Q7���$���A�1�O[u��*���>	�!�X~�h�z�>G4n�,���-�wH�m��=rƾ9K�NH���
,X0$_��X��Ɂ��a��#�1�H{�~��W�������:G�[n��;��߉�K����Ft��M����T,�z��f ����{}�:-QK׵o����de;"�$Ҏ��'�L[���յ�6��5���e�	8
7W�	cuF�v-��#�<1o`��!�~:o�Y�Mut��e��wX��x��iznQ�n���H�^0 Ia�ƈ�o���h�޻�ڣ��{���:*�DC���qxpp��՞�������7w��+w��9����)���oj�K�0���jYu-�R����U#�H7�d0��ߗY?"��	7tP7����`�4�����Z��~�s�n �?���/I=�n؏|���AI����$1����M���F��=�#�.0 Ia�$���;��#�:��8����������T��(8pϠv�s@;4�� ن��&��5cRd¬�RbM�(ܠ�^�QxxX��{ID$����q�XҘ����C����yŨѫSW���,�ѿ-�ӝ�Ȏ��9���KS����Ǻ��ju�)O����O�;cӾ� "��I�6���ҲL�k��QG��$��uGf�-.����Gq��,�:�P+�}�0���Q�V21Z&�Iz����St�|��`t�3�����c@""]%���K����2s1~�l�Q�F�J0���[�����5�F���;?�Ç?m@YE%�d��m���_��윑���M]Y����b@�¬�#ڍ�3��S��=��?0P����ב(�]l��iwWg<44�OQ�$���b���7vo��>�k��IO��ۄ#A���t��ջ���I���$�I+��m��==�;�Cjz�'>^�=G�a&��C��Ѭ���i�MD�9�݄׿]i�)d�N�+ߺC��v�c�����3SL7�FD���$�Vs��hZ�۔�Հ�=�Z��f7�.���rwU0���N���0���|����;�4�o�������WO�윉э�؈Θ8}5���I
�6hXŎ�IL�{��A�N���`.̢K�0|������}���x{����5��2����{ղ�w\���9U�،���\9���8|���hѢ�Ν�	&��Ym��4j���9���Z���cԨQؾ};�iH˄d�IWt瀶��e̲����/��ۯM��Ot<qS7��=���c�g`t�|�൪<):L޺�:�;9�O>��;wV�<~�x=z�>��&�~���1x�`�ϱ���׿�������1 �`ҝµm���3��U؞�]�s>>y�)��I��D�> s�W�u��t1���	#�P�O�+�u�fCz&D��>	�v){���o����������ޯ_?";���L-0 �`��_���Wn�omys7�S����~��t���o�K���큏��[4��_/CIY�JL�{��y�~FZyy|o��n
��@�H\]/�hpww���{���5�\��wrrRCҴi�@HR�5FX��g��G6�=.û�jv>�h|�~���)Xo��_H���]��q�?gz�ͬ�i���}��v�y����~�D��U�V�����D`b@�ƀ$�Y��,�c�0�>>o�{����|�������:="A�E�_:�6u!#O+e���׬������iز����-Z��
��Z/QrtH�V��:xtxg�4��|�,���,U|T0�<5�U���O������B�1"��w��7�kr>1��ϻ����SLQ��H���,�j]b��#�����q�9� �$�'��s��p����/�d&xߔ��㳿��o͎���	��/y���`Db���y[p׀����mL�k��H�7.�( 	bIT�st|
�`1k�v��j֏�.�����ݢ�G>��ҥ>VĢaL$��//��A�^x�e0�׿]���Vjg���?���Q$rH�z�BE�vE\,��3���V����m�mD7��n*���=X��0��ሮ��!����'?Yh�Σ��R���2|�� M���7n�d�
�Du��lۊ�}��1 Ib�'\Mi��L���{al/��jse���t���j���m���ߟ���*�w�v�6%ԤĆjr��Fu��Ui(8[
"�Vpp0���c�82$Ҍ�#HTC�#5-��ƴU��+��0Qm�ԣ|<\q��?���F"���{�.M����n�d!"�ivHD�t$+Ӗ������k��C.bg8��ر�=;c�1�P!i߱�x������N����a)�b�V��-�����Gj�������1 �.Y,�ɬDk����C̅�0Q}�L��{wA��%��Q=۠qC�z�KTz|dX'nKE��޽{�l�I16b�GZmh�������q�4;״e;�۞c0��q����3Q��ؽ�����`ť�x�����񡚜�k�����8�DD�c@"�p]�}��59Waq^�j)�$6<S��Yq
rlw\����W�,�Q��nVl�PG�ꋣHDd+|J�`5����U<9��f�zYi�.(�QD5����G���DZydX�Z�俿l�Q<��<l��^M��Q$"�$)�$�~\�d>b��[\�&��u�>��F���/�R�i�����ȩ��~/� #+_]���&E""[`@��b�ƿYsiB�Ma��#Fb�H� ق�łɏ܀�/M�ƽ�a����^����>ר^�x����'��ıQ;g�ępv���ͳ�5a�6י3g�������Ɂc��j?��Z��sj>�^�k�ja@�¸��W�)vt1M0�sKMε��I�ܞ#k��yz����Ȗ�H�7O߈��N���\������6hR򿡏n�6�P��L�G6�1-)��k[�޸m�9s�`������y����Xp��_yE�z����gU>iG�{�YC���:jU�m��k`/��nq ��F~��������(���I��lR�Pi�.�����ͨ��mC�H���n�޽III�;w.&O��$�%Q����1��59�����a�@T��� ����xi|/CLC�(?����\�s5m�!�[a��4�Eaa!^z�%��1 �>Y�hb푘���I�W�����Gn �"��M;���ֻ�~ިI@&�О��4��D��;�1���m59������]�;�`^�#��d��}��~�Q���e�ŧ�6���}��-��C˦�)TAD�ŀD�ѲH7�5�^��h�-���:�7u�dL��S[�<5���*����O4	H��<�����������T3whT�[l���T�]��&x\	HDz FTD`��󩩇��1m�M�*��
O|��\)_"��a@"]b<2>QQ�_�暜K왢w����_��S��B�E[a�>}���=k�&���C���ۥ�ADTWH�!6�w7�������J1z�Ԩn�n "=������_"��zu�x~Y�7�������ŀDD���D��r܇.p�F����E%eг��Ƹ{`{�Q��_��/x��Y�4	H]ۄ��9#+Df�����d�i�M�6���,��`�Z����'N`Ϟ=HMMEU+_iF˙E+��YBT0�C��l��9;Y���ԯDz%��}2o��?�J=������+1�^��"�~'d[ ��pww�ȑ#1j�(���OE������˗c֬Y�1cΞ=�3$ҎU�D�usmF�~\�9g��gMQG����w�C�����MY���I٣&}���~�4\\\0a�����?��>�rk��^	!������7�ҫ��\E�X���˧(HW���{� �t�����y#"B���w�3���s7���y���~~f����C�ǌ3��Ga�����������Ab(�{;<���s-�~jV;�^
ƴ�e�@h��àVk6j��puVtzm�?����F�X�p!:v�(���+W�g�}��cǊ#<<�$�Nܭ�Y����O�&�4�a�u�YϞ�Ύ`L+>z���@N^�('/+���=�)>������5i�7nD``�Ş�M�6طo�C��q@bj�}�5�pQ"����f�z4��Ӓ��^�4�-f�x���;�H	H�B��_���Y���X�n]���ڵkزe�7���b}ѽT�X����С��郪U���j�[�fڶm��W���q@bq����X��B��k����h ��#�:0V^^��m9��Tu.��s��o�!�rE�����6;�i�fͺg�9s�X��bŊ2M�������A����C�fwވ�����_����q@b�H�GEE���k�R��h<X���nMP3��i���3�=�]�c�m?��F(�	�mvL�jժ�1c����s�aYY�0*((�ʕ+�~�z��\�Dmv�N�<	[��I#�����iҀ�r�Gs7��Zq���My���}��I���zJJ@�6;�UT����l}��͘8q���H���L�4	6l�]���Y}s���J�S�l};�o[Wʹ�x�W��8:�c�!����t%.G/ŠU]eӹ͎im �o~���p��s�; ����q@b��Il���m�H�Ҥ�?*y*>ϮSW��5����"�7'���z�u�J�բ$�9���w}����ҟ�^�"%�,�$&�̶8NG�ӫem)�Y�C���z��H/m�7�l����,>}�����jY�,�ƴ$//ﮏ���J�{����l$k��"('$��Ny{큲j��W��M���WTe)%#����µ�������j+ӌ�Kl�݃�hD��y�>OϞ=��X\\l$+���Hl=���)���.B�Z��"2s�FC:6���WgGUW���Ni@�#��Ŝ��ۓ���{���g���c4���EJLL��*Tk��m���r@�юƁ��À�u�D��ZM�����ý�c�ҽHNφ�l:!�<څp@b��a�ddd�����5k��;G�Qt�`��hܸ���:�0��q@�h��|�S�lV�zʫGd��+P��U}ѩQ50�Gn.Nӽ	�[}jCm��qlhce��u�����<�iDRR�������w|�nݺ"$-^�Xl�z���2m۲eK<�䓘0a���������{���HL�S�x$M	m\]�9N]���u.}r@+^2�t�������ê�/h��H�ɧ����3�iŻﾋnݺ�S�Nw|���	>��8RRRDH����͛7�yj�

B�6m�9�Ç�7� �dE�k�+�
�M��_������{����ޭ1�3���lQ[�]���:}��	U|��&�9 1M���ŠA��r�Jt��垏���F߾}?����1x�`dg����8 1U�!���AF���]b5kG�ӻ��Qe@�.J�ڹ8)�d�ܸ�*�+Mrr2z��-�)���K����z~�x��/�ī�����8 1i�츄d�:7��6g�Jg`��G�Z��t!J΄,�hU��hߠ*�Cb�D��)S���ӦM�E�uKk׮�;＃�G��݉���4��C�U9ޛ�O4���l��ک>>Y���Df���!1�;y�$����@����ѣ�w� �>?!!;v���m�D����������k��t�5���C�����\D���%�;74$�큲S�E����i]LL���{qZ�D�����nj��A�94�����p(�GMhZKNue�J��r@b6�n�B�+#������Xdd����Y�y�"��LH�R�	�T�#�	mB����	vt�H����10k���*R���nZ�ڳ�1�o������T
��h����]*���#f���60��P���"�F5��T�,�yd��$�J\@҆��U��^7�]]0f��M�mv2�*�;�p�b4c�$��*Q�3��р?á�4T�D��܊�l����E&"9=�<]��n�p@b������տ�R;�u4ڛF|�̀�ua�m�̆�Hm5��m?qE� *A�]s6cj7v�ػ>�n�:ܼy̲8 Y	_{1��\Y�9NF�A�x�7�um����9y�P���RH0_aڰp�»>�~�z4f��r���ի��z�k�.dee�ݍ��pB*O�S=�1�ۓ��(�6��l������������$+>G���;�YK�~�0}�t���Ke��5j���o,K�"͜9S�/''�6H֢�2I���t��)"F}�6�n�8d��э��h����E���O� cZ��/���������y�>�����Ʋ��>F������U��	��
`rɚ��c�TO�]Xw�emR�1
H�Z�5��(�<�"��iٷ�~�.`��_�NNN��xӦM�{�n�o����[l���@��N���+݅U*B�-v�6�eL�Ժ�ZB*��y):U��Vc�,����l�2�k�����?���'�bŊw�U�V����.]����IO8 1�(�q�ѿz�z��\M��Ș�ǘ�vRt���Ę����cժUEzz��ǟ={���Ø1c���5k���w���&M�W_}[�����!jq�M�d\\D�H��PeL�cz��J��vo^S�9��WczЬY31�nȐ!(,,4����x|���駟�x�b1��x�|��w��WW帼q@brIZ��K���_��*\��#��Ԥ�?�&"V�{G5?HL{���+�rӘ���C��&O�l�233E%��J4����@���7n�-�d-z E��؁�������շ��3��f�Mk�0 I���$�Eyyy9r�J6��������|���&��B����:$H���^�NH� Ū��Ԩ�c�54�&ho�B��e�\�!3j@��1��+U����?�;f͞=׮]�LE��[��6c�HL*;Yc����Ůf�J`�����:A>�~j!�#��"�o�1��J�СC�u�V��ܞ(����E���}���t�{M��T�r@��n�*�ӯ�N�hOQ�H�v�\��;Ѡ5$r96��Ш�W��,j�{衇Ġ;�����ܰz�j�&G닌����$+)*���2� ������b��.��}�DHb�݉����������9�4k�ҥ�̙3�����6oތ�]��ҥK���v��w},1QΆ�Z��j��"� )���ˣ�nNP*15jS��Z1vO��xCm⒍��bL��VaƬm֬Yb��O��it[�l���ȒG�<����Ry�;HVb�c�Jeg�� ����򷍌�<�M5�j��=�q$vzV��sxy(���{)7K-a�k�ѥi����9��R����ǔ)S�q������ի�uJݻwGTT�]�G�&�~�o�6m�Z��xnH;�::���5{�[$�gyR;H֣ŗ`9*� �V�b����٪����3P7Y*�s@������~���S�Ʋ�i�x�QTT��'�����=��ԩ�ݻw�JѩS������/�/_�*U�����/�	yja������L�v�|O�q�I'筅�z�:ɨ �/ �Wc�n�*lE�q����+Ӌ��\6۶mC�֭���h#�cǎ����>G��K��:u�\���Lҋ�_�����
M�b�ݍ��8:�#��j�.���-vLcjժddd���OKK�}��'4�h����F�S(��$4oɒ%`��G���\��=W'��PcI��*�����i��yݦg˨ q@b�Bk�F���s���7n�gϞ���?j��j��4iX1�"`R��	��k��#0V2GC@�z^��b�lTNN���$''�w�����/���}��裏";;�$�Rz-�i���M��8�΋/�+����QA�1p���D�V�Xa�c)�<��X�`^y��o�Ӛ%>{�llذ�N��`-v� 4\��A�7Z���+H.Z�+{�$m����g*wk�"�--�m������Ճ��'RRRfR5�Vq@���i�lt���)I�$�X�d��e�q�Ņ�2�[�z��seff����`��w��i�DR���N�Br�cc���^])�o�0�,���K?z'�N�ڦ���-c�R[���
�Ab�����*q�H����1V2�iHJ�R|^w�+	$�R��a�ns��2U�c�%$�JeϯƘ�d%T��Y?D���Z������c�1�V|�b%vz�� ���/<\��&4B�1V�B��F�]������1����pBb�/��T���1�((T�{�������|0�ؽp@bRف;��MF@�p�Ę��嫫�"�=$'�c��8 Y�Nc��}�x��j�H�*k�c��Nm-v2����b�+$k)���R�G��XA�#c�+TY���u��b�+	$��iI^	�阧
� тm���{+���ln�c����ը뇍��}��+���Ԍl�y{�1v�\=�A�
c����+$L�r%\T���t33�c%P[�ENI]��1����+$��q᪕����*�p3#���Ѻ�,�$����e�1}�d5� v�*c����Bzv��s���v=	�C���SrZ�F�{Hz���2Ƙ>q@�}����A�;}��*\����ťd@mdT��S��ؿ9�zb�m`��ު��j���d5\")�,�
����j� E&X�M�1������2n��k�1VHV��:�����Y�k��q��{�KV_I�f��*�{1�ԁ�K�"$�Y�E-vt�8���A�+�� -+j����{��������)�c���J�	@�@�_��ةM�J͠����>�U���X�ETB��j��c�t62j\Y�9�8 1�J��Z�z��S�l]X(�3($�GU���1�hR����N]���U���<��1VHV���L�hѶ� Q7�jC��9 1v[BJ��Zњ�P|�����PO�/cL]8 Y�^g4��|�#�CT�N_�ǰ�`�;uE}�#�>+��u��Rp@������I�d�ǭ�|�l��ā1v�R]	��=c������!s��r��k�\QQ���ߣ#��pv��l�����5��6�&��"��72c�i�?�1��O�d������+!իZ��Q+����foT�t��i"����T���Y��Ȧ#9yH��Alr:.�$�r�M\�5�����,t�ie��I֞A���*�٬�Fj�� �5czp�Z"�F��EZo�c%�d5e�C���&��Ѵ��XH���{jSr����nO7gq�jN4����8�:��g"v5�y�`�$k� �������_��Ę18wM}#��J�r��0�XI8 Y��RK�EZǆU���p���y�� �q5q``�1
GG�^��㗰�D8������\0}�'
��o��	�v�2�d��k۽	�u{�F��nm)U}����+H���p@R	Z�@U�":��3cM�N��м�8^D�梧.^+L����p$��!-�JK���#$��fϙH0Ɗo����G�!tx4$�X�8 Y	��uѩQU�QM#oW蕣�=Z6�!�g��C!Ά_ai�1�q<7x�>M��VJ�[�h �%��S]n�c6n�i��,������Y�X�8 �3OwW����wB��Ep�E4=�qݪ�x|dw�ݸ�����M�q��U�
Qv<ML�dL��q7������lZTb*N_U�;	Ugn�c����8;�o�&֧������)�rE<5��8�F'b�!(-8|M��c�$c������M�����ZOǘ-�}Z}�H˺����cFp@����n;�#&팺��LS#�/N�g,�ڃ����5S�ᗱgP��ձl�9�	}�������٢]*|ϥm+ZI	H\Ab�����hP��a����E]բ��|�g�!=;W�sD��\��Fz�Q�M�d2Y��1�cq��9O`��Sb��>
G2���D}��kP�Ɗ1-�+(���6]�2�qo'Ƙ�p@��a� ��`_���延�6����$��ld�ӳE�u�dd�|>7C��ɕSqp����U�Ѡ���(�j��U��#=���m�ժC�����DĬ���R��6�s�#۲=�9 1���h����6�%���,H�1�8 IоY��P_��d��S(�p]�K�Ɇ��^MDZ�ܪJ�!|Б��kC���{�k��J��TI���`Ch�R�׀�К
J/���ŏk�� Ȭ�pX4��6Pt�Z��5�C�s��x�/��͎ٖe��C�d��x�c�(H
�h�/M�O��c)1Ii�s�Z�a(jۻ��Utl>!��.%����X�Z� �U�E�>>����PL�F��oW�d�� �hQ������tZ��U$fK��~��p�ME4��|-��1`�1c8 ��_��xi��jTS���'��ȿC��X�Mq�CNnv� �[:��'���N-C�=���&��I�����D�]B
o@[^�\M@vn>\����ti\Mu�p��5��F���NNgmp�c�p@*�u����B��R�K�E�>�%;��dD4���f��^qws���-0�_;�h�P���t�g�o��}Z`���v�!q��,�ZU��� �p��ղ6Ԉ�옭Y��Ԩ���BC�q@b����	��W���bX����oiFv.��hۉ��j�6�%�������[�F�m�Q��C��� �0���w�c�Z����d��7�0���4 ���޸�5�;��v����__Ș�Q��CaP�.M�W�N_�!�1ƌ�T
�ئu.��o%����gE0Xu�:��5\�2���4|�x�8�T���0���UQ6-Ч�~v��*���V�8y�2hP�� [m�,�v��	s7�@~A!Ԇ��  ����1f*H%����<7 �C��+&!E�Ek �f��Xa%?@����[��x|��*q�:�F���n�.LV���7G��%{0{�~r5I���r6�5�߶���К@�ߨ��+*����(�H�:��g��1�L��_�oҠ��M��Iٗ�.�g�ۈ�k��V���	 {��a��,|�p7^���0�\���㺠O�ژ��UV)��Fϟ���&5���[Sˍ�W�.�o=�'�czE��4$H�:7��Wm���Q`��?T���/B��7�3��0s���R��8.d��Q�����F|�t/�����Ѯ~0v~>o��� /M�g��ˊ�C���%���'4a�-C�vs�a՗1����Zu����?J��	�JeGvi7����kS�<7P�:����˘��zlګ�q��F���KN�������mź0�]V�Θ��}��M���z��)�ڃaxah{���._�8 ����>㩁m���P�h�qu��-u���I%[��g�
G�1�s婥���`�`b<ܻ����q�<f����k��|a�]�~�pf.�)$�F��^�e>�=3�����SW��9����B�?���X���[��kG{0�'_�yH���=�H��8���V8*��:H����=��!��9�����Ǯ#��7�*d�J��M�g-ۏ��c;��Ae���[���������w��W��j˱��@�yhR�8������?�_T�wdLMnf���MǡV�z4U|�ys$�'ر��+f��ڴ�~��X�o������������v�ILH&|���h���m����Y퀲=�_C9:5���f���X�`.ja�Fum��~�5�u���|o��V�ڴn4�r�硛7E�����p�J`s���_���X�`��g����+p��y��Q>��L�t��3W��_�X��xk|�2�z5�];>���؄%;π��5%��~���H���Q��4��5���15�ꑚ�3���H�y����S	�(7� K�J���G�{���֫���=�M���#ط�w�h1�Թ۰d��eg)�x7ˣ0nEp5��j��؟=��Bζs@�ȱ�N?��_���ʽ��c�0<�a�>�֣}��@�hQ��v�ܕ�����x��>CW���Y���=�ۺ.���6�QHR����~/t�f�0v�R*G9���l�YiOUd�"�*��:��{���D\��:ܬE�n:!�h�ddC�Z�$�In
�䦢V~:��g�j^|����p��5Gw\s��UG�s��igo��<`9����L<1�O�wͬ�����W�>t������?].�(���9�8 ��]�6 Ѹ�;�`lw9����W�h�u|(u�R� ��V�mu��~��HC:6���}���4Z�B�Cҙy�!�4�IG��8�&�݄��6�.:���S�pʹ8,�r���|��Am��+����a��~₻,z����o�ƃ�,��e�j��⨴���/~�j5}�^�V��HL�hr���Ge}�.	Va�o���t�h��z�����<��
�$Y�$ZT��H������Q�SW�֫0��	�%א���W��s��d;3��$�!���f���S���DoCH6��BU�u>�Q,�c̸��dqǶuH���x�9c`�zXs@�7W�R�ժ�R�~b��ѾG_�T�8}B����U|j�[���̲�p8be������0���e��oW��ZVɉ͡����d^G�|mmf�lH6}S�1#/{���V�R����'���Pk�֓8f���65�+��y4v�BҰi���?3n��K�ݵ�j���~<г�Y�p1fM��ۮ������fVIh���x�wX0�p��H���E�>�]����u��b5������Q'C(����2��W��և����.����_�ev�2%����({#��$�8��������[��NV��º����iy�tk�a�]�gP�z��D�K5J���ǋv�'��1������95%��n������p8bf�]@�]�i�QY'����/+ǻM�$jQ�v����Z"k�3$׶�i�xװ���:V�!{��\��.�i]�S����4��hS�?���.��Y�®��dk�=��m>	����8������1-x��6C�轶{�ϓWP�돘!r8bf�U@�!s^��Z�)���PZoT�c��
3�̍�`F�E�mu�WblA�8�ڹc�c0V9V6|�|��x��W���Ja��.X��<`�t��L�4;����D^�yV�;��ݢ��5ե���l>.&�2�f��ሙE7���?ֻ�����0��M(/Ջ�19�:F�'�	��7iT�����J~�0�?}�GA��_#}��a�[�Lޭ���	�^����5M���m9���v������6��zU+�b�z/�v���<���YRZ��j鵵�=ܻ���,�v��Z�98�n��O�5��6/����F�W��$���Yx1�:F$�_B�R��/�.��H�~��!(Y��k����\Q�����Ӓ7Gb���系�H�wp��Q|��m�g�Z5{{�6�iU������=w�IjF�tCD�̜<l:�,����*s8�#]���V�p��竰r�yXZ�����AI�-SL\��O�.���X̮��y�F����|�S2D%���h��)h#�?��ƈ��pH*�����to����A���QQ |o���cjCm����ڽ2�����hoZ�Ę%Q8*���=�#=�|@�}�ʲ	m�I����ʒ<�
�R~�ʏc���̂��i�<q�"&���W�kZJB��g!~�|��X�U|<E{^�)��dv'��{-!�����y�k��6B�~�r}[��71���s_����h^�jH9�#��̡�D�nޟ�����f���ͥ�$����ah|~�ȋ����lm��*z+����w}Z����Ş�*�o�OƋ�;��xZ�4��:m�ؔ��Fwp��+�C�둾-���{��5{�uhZ+ �˰�c�DߓT%W��Ft�r����|cL	���5����C�pS�&��.���*E����^)`�ΈB��8����=kZ�y>X����1��>&=�m� |��@L�l%؝ҔQ���PA}fP[��G��n�c3Va�G���Ę����7[��]�`tjdZ{�1߭>��mc��4�h!��7F���L�x3S��d8����"T4�������\|�B{��]t�����ɭ���[���rr��X��o��cx�U�����YO�+z���]Lz������P|�d�m�b���e�lQK���3�؇��l���K1�d��>�3��Q�xKS���#�=�IJ���<��1�����;e��c���w�zb�E�<���Y�ḯ0VC!����(�����$�9(0e.L3!33�������zg�`o�Z����<�[�9f.ۇ@Åy+�O�d�1��}�Y�۾[sXJ@ruvĤ�m�Ѣ�P;jl��e�v�1r�D�pV��ۼi�Q�������;ƭΌ1)4�h�����X��ՒS��+H�����Lՠ
����y�WG�SRss+>��BSZ��#��6�jҏ�{�?3
/���M{�6|-�u�vv7upì��É�8�o�X���,���Q|�����+��j������у	V>����x��-���9y�i�=��`D-��1&��-Ԟh8L����-���CQ��]����Q(��[a��o��opu->����;���o&�}�e���G"4+t�aW��2*���7tiZ��c��F�C������DV\|��� ��O��=���e��_���?��
���MkfL)
	s4jV� ISi�f���2ƴC3�Y� |�Xo���?���|
r���_w�(y{ſ�i`�7U���J��%$ qq_�P��?����6�WA~[����a�����1T1���A�����ZXX�����>��Ɩ������G4�JC��g�\��^�,m��+���q��$c�%���oW��3��M$oW�2e�Xd�w�m���I�s4�M�o��P-��#S�"C��׷x��Vџ=8
n��つ$Xj��75+�Zg�A)�δ�S���#�[��=�ZU��>�֞��=����
����tU|._/w<Ի9~4�$-Xw�ޟ�S�ߝ���G'a�t�LҤ��Fui$�\t3Ԓ�w0��n�\��`�C�'������Pk�Q���u��ŭȂ�b4d��D��ڨ��V%��$��W�,�z�Pz����P$9�kmJJ���wa��������_��g"q�b4Xq��sCۉJM�I챤��H��r� oC�k�dK�������_�b��ݥ��oD� ���]b9-k`H�CbX�i�w����h/��|�'��\f�T	*���.��R�P�jqP����e�cK���0g/i�JL�v�!�gG�j��9�e�h}���N������F�O����Z1�Ǎ�W�2�7c��0�?^.*HZѵi�����5q0�+��h�{�HT5���i�u&�d����ء�&ƣi��r�>D4؀���e��Q5��G�w��OL����,�OQ� �7a\�n8(qx�sCm��>���c�j����Z`I����Vd-x�+��|g�&@�

�Ч˰j�84�&��M��X+*�Z2������S�{N�����?�C�",�TEv��>wO�Il�g�c�k�$څ���܎3��JǢB|�p �үB:��ԩc#c((���FE11R�(y����m�CjH�6N�ۧ�	��h���S�X��<lMv���e-Ξ=�z�6Zq#5Kl=����"<3�uLh�}����}�S�Hkᐕ�=*GK��_BA�P�;{0FT��to��!A&=v��=8p����v)*�Oq{�?S��
�ƈ*'�|��TQ��;��ED������I!��*]�ݭ���>>sv�x�&�G�*Җ��Y3cI4m�B�)_7cZ��=�a�֓Њؤt1��BRO0f�1Gc���V�[�H;W�t���8�{Qe@����L\�I������$틊�e���Ԯ]\=b%sw7.~�j�JPHZ��{ᨫ��;�@m�t�k]�4�#��mlU�h�'��r>
��\���,P��"*I��#%(2�������?j�V�p�H�81Pe@�
I�������#�!�M�&;P;ݭ�T�q�5��;^q���"�.E�X����9g9-��E�
�Q�[ƞ����q�s6�d���.��@7�h����1p�����$��n�{���nYڅH;W�t��S	��΍�cl�&&=��Y��pY^M:�GR/I;��5hP\ae��T����rB�Oa.~�فA��t�I����.X�4�����8'|�d_ywlMޢ�/~�o��.iklDL2�U�jVc%)(,�m�T;�?�xJ�`���#�"�
H�v�&Ӧ�ѝ�-�.K{�i��J�i���RK����j�����<�㲫da�!$���7��<>9�O��n���unR�z4{��:�@�ĀV�_U�����=_������ߚ���G�z���d�%+'?[���,3���h(���ɒ�`:�ሩ���ý�#$���j�{���Ҟ�[Vf%�s2n����׼����������z"O�H��i�p�.�9���w���/jjSGK�;�S݆%o��r�浫���hl�:I�����㗗��V$�n�5{����c�E�]ǫ��V�u��x�#��p�TH5�����5m��{�w��24�I��q��TT��d���-a��)c�p����e .N����$bF�!<�|�R2�}x�gS�#l}����<�����[�_#�ex��n�s�i�剪�?�Clo kM�m4�c�G�p!*Z��3������jishfGL�T������f��h�������ݨP(aR��3а!�7�4��Q�"����G��O��pg/��nh� �'1�6��p�Ra���evͨ)Zl���_?;c��;���j��X��	�xzP0�u""�>X�ɰ�S[�,3���z�����" Q[���[����^'�9�b47v��+?��+Ш��.Oի�#��俙t�����=P�v���e{�axh運6��`w��������6��q2�iU��~�
���(���I~󗭆���|Z��v���]�3_�UE��U��X(M��v��Vxf}��ʩ" Q�)w�Zg#�<�ǉG�>GB��_�����W@@�Z�DW�f�H?��E��>��|�2UD���#�FK3,�������xغ��ƈ.Q�M�M�O��pJ�_[bA�ws�E@%�P�V�\�O�gT�fu.N����0�,o�ق�<�_L�r��i��R��~�B�j3�2O��Ĵp�'���xR��д@��_����̫0s���>CHʴW���KN����{��F��<�M��غ��L1.]��d�+��e��nA�_�F�W抐���-#;��߈���B����锄3ȜZˬ�����iw7�qo��UL�S�??�eL���F��q8R�P6$�8$)���(�&޿q���*�#}���иF��i8���{z ?�=��]�it2T���o������L��Q����:��#;��������ոZ7�S<Ի���QՈ3��#�!VHtah��*�q~��{�.�����B�}ݴ��28Z=_�[||�5�+W��*��=�a����i�m7i���cB��mH�anĺk�dؾ��>��մ�����]�ϓ�G�O������:�4�~�utS��țZG�Zy�3��#�1V��a�i�?�}���{2�"�e+\�@��2�#�	rr��E���p���G�����PKȹ�D4�^z�I�Fո����5{�~���,?�Kܡ�-ZG���gO�5:��[LR�|��7Ջy�������:s5�I��Ϭ��� ��:A>���x�("&YLS*(?o$�Tv1M����:�NTE��Ϳ.(�^y�״Ɋ��d����1t��R1\1�sC�5�G�@��­�˿hz*�-�j���?1w�I�|�>Ԫ���<o�	�3w��V/h�Q����Η�_�I_��2�p�4�j��D�0f��R����Q��JXZsě���;խk�������㩗��B-wQv�N��RȯX�����
4���њZ��r�Xi礯���{�YI����SW��O�����AZ["�z/x��u�w.
zҿm��/Ӭe�E�i�#�aV	HU|<1�K#����ɿmQX�1��a
���sa�G!��6�<Y\M2���y�a��;{E���؇��P�c�<iPL�a#D5�6���7�M+��"�"�&�J�d�|�d_tkVL�h��[�������R�I��6�e��i�UғZ����E���ʫGE��T��://�Z50�5b�Ν3{�]��$<��9^u�Qm?��㻊�۽�跧�	���6to^5䵐}�L?��w���rl
���څ�V���\�V�<��9[���6�^jtϷ���:�p�t����!�����=�'a�]���Sp���T|�mJ? Sڧ*8�2��嵤��ݣ��-<��l?>}�w��quvĐN�����`@fN����7Ύr~��r�,���yHJ˂ެ=�m'���a�����vgE'/�a�/�t�����F˺�R����=�Z�e��N�{@�Ӻ��y}�7Bvn����-��f�ժ�봫jUÕv&�d����\�x�,��i������xet'�z����qݛp@��(�.��>�U�9i��o������74��F���)�:�ʤ){&M��M��S�-���F�#:˝�H�����Y�#�#����hb�1�����*~�gn��f��U!�vQȭS��M�Q<�O߼���!��M���U��΃�J}M�jS/HV�.�:7�f��KS5�����i��WQ��x������ ���B�Y�9~��^�R�w���Ol#��tC����9U�Y9�#788;��rC8�?��hz�)o3��*{��w�:FG?`($)�W�-.l���V�����U5k��~p)*īɧ1ٯ��?��M'�$�H����.����:��(�=���Ҵ��t���ѳ˱�x|�*��c����5��^�4�~ݡK�T5��pw��}��M�)��T���_>z����f��G�4�ž\Ҩ���$cm?���^K:%.l�V��w'�&�af��Ci�һ!�8y�\)�X��<�t,������1�p����/s�D�)?l/�z^���=)WTZ�L�r��߁g���}�����y6�#[��AU\Zw$�]����s[��=���rH�Mh�G/�(z�y���l���Z�GTEJI
��i�������E�%;�H�.N�צ���Q�@_�6����<ث��0}��F0�KlR:ޞ����݋��aL��hf\zV.��:�����T���0����~ދQ7D��i��<0���rH��TB����۬|ߣ	i���,t��zu0rq)���̩v#ӯ�C�f�vt����$*I�Z�h\3���3w;���>9�1�b���}״"-+?.��_��4U~�
������9����($ٚ:A>�c�h�8ɽd����	���E���@�s���t�oҤ�ە��]�1!UA/8�w�l�3S1ZW��"���OS<�n�3xb@�RӧUm���-^��&����X���'����V�ٓ��Fj�ͬ%��Q�xc�Vq�P�z4�}����3ZȻ�H8~�x�Ι�U���V��w�J��g�\#*HLc81Pnɔ	J�OG��%&��û�̻Q@�*`:F��h}��N��JM�eg���"�����p�"�o�?_��o��o������v�N]���s�q�VtǨ.�1�s�;���D�N\{I8�������3�ɵ9�_sXTԙ�p8b6�\RHpe1���pT±�Ϧ(����+�V�*U*�4����Z���i�1ǫ��O<<W�RP3����7\�r@��u��0{��0���s�7/�#�ԕxزě��v�!qT�tEh���ڴ:z��%Z����*�����@LC�jĊ�Z�ߧ�2�>e���]�iLy�#GǿFys8b�Q.�WK������c��󊞧Cv"���dWW�re0@!�6�5��41����D�m9���K���.H]����0Ң��D뺁��D�AWg�~<F���IN����Ah��u���R�:U���������g"���Ul?qa׹��^��n�;cм���

�|�\��2)�pT��YY���Ҫ��5��d��M���*����&�)h���S.��E_��р���".��7���茕���W4��q�`���v[bj����q�UiV�
Z�S�:Ň5>О:a�#<:������Clg$����rմ�bp�l4d�����4�
����Y< ݺ�3f��0E��S������d�P���!�)�����ƕl}#M���CK78 ��FjF.�($�FԲ�:e(^�n�n>V��i���[hZc@%O��!ֱ~��]�{�x���Wj�*��F�!:�'�"�p�$��ZB��*�75OU_/�zoj����*F���������(�$
GΎƿ�w����yF�_S���k�l����ͪ"����|[#���̈́w��4�Z��l+���d����|w,\�忥�|�>qQO�������tД<c�-؎�G���~\TT�ׯŏ)����6�JW;����@��o�+�9���#f�,�Li�;}%^쇠��t3�N�Ho��&U$Ϣ|�Ɍ�Z��f?���W�ܐv�>�n���W��X�h�ؓ�W㗗���7;^�Y��Q5�Y
@���8���5���ݱk��t�,�~LCt��^�AVN>�~U��H����M=��҅�5���*;ɼ�}}�G?3���\�"~����HEi�9� а��xe��ق5.��9[�ѣ�,r��{7��.�1��=�~z�~1��(}bHLC
�S9zj�jD�$��׋�;��]��ע�.&�0^��}�̵C�q��9��6Û3���e�fE$��<�ۛ��pFv.^��v��K}\��@,���?�="FR�2:�"�Ծ�h������0fm�m�w�f��SK��1)�:ƈER��UMjw٩pS�J�3x�4-�0�"���ͮkV��6;���рdB��Fw�]�-�G�u�k>��-ARZӢ�^�Q]Y��4��OW�8o-�p���,�L����P%wb�
��1F$Z��W���^�1���ӑ�<�S���*,Mh��m�4����vx��v��f���1��x}����b+K�pD7�J�4��cw�l@
1��V�z.P���)Bk�(,�Ĕ�S{e�*zjڗ�6Ivq*��HUX�S��}��;s��mh�%��K�?~X��o;��6L�,=��\��!�m.�4��cw�X@��:�0И]�#=O�L37���*n�c�����g $7a�^f=-���篣K��>�i� Hf���F�BU�~�:
_�8�i�� cju�����e�s�,(���Ñ�p8b�,�h잛	o��O\Q�<��fn:G����֢��K��ͷɹav@"�fg, 5��Vv�EE"$Ups���{Z�ޭY<��r�Y*cj��c��x�V}ڠ��Q\r:�Fp8b�DH!�����~���o/�/h�Q�fŊ@|ٿ';g�aa��}�����iZ���($=1kr��1�{�=m��{ƣ��n㑲�Řl�>����b͜%Q(��"GZ�ሱRY, QK�1�1I����ܛ�F;����;T�`V@2�����h�{4��j�����MH���Z�{K�$Z���b���?oc�ҭYM��������Q9���J���cFY, ��dʅai�νY�R`�d�[�ۉ���T͌w4o�+q)FCk�h���f��c����\��=9�5:5�&Z�x�+o�i"m�hi�cS0�%�W��3�U[�.)��8$��^��ؿ�$3�!5�M�3�����V.�1!��9 )D!�՟6��[:$�M��3��_��ڃa`�Ҩ�������v<<c>����`���$\��Ė`���8�j��X@��o�n|x����9f,3+����º��*j75����9Y�+$y�:c�+�������F0f)SF��1���\{�\Ø���,n��Ge�h�]Fj`go��H@���"z�Q���ɯ��w���0v/��\ew8.��nj�Mf:
Ia����=�Kl*kI��kB^��M�z�ǵ3y�����l��,+��Ǥ/� '���LG���ER5?�r�ö����^�f~�f~P���,1�u�����EDL2�NjҶJԪ⍥o�ºCa"��8p�Իu�sCڕ��}��0��u�hUe��1�X- �����9B�̼c�����̓�^��p� YUtN]���c�-���h^�����{�XY����_��峞�#
HLC81f6$�k%����5s2�ױ�88�5���0��ȴ7�%u)ڔ
�A�ڋ��k���D�Y����X/2�G�6���)�}+���cD�����Y�x�uX����p8bL�� o��	W8�����r�c�$;��,\u6�A{�������`��$��J�w�Ġ����9�*Hmw��㵟6�HpvO�nΘ<�#��.N��tj?�a
^�r��1�,�N��a�J�lf��K�|3G�r@b���Hj�[8�
rp�h�E��-���3R2�_��JGS�&L_�����{�ٱ|~��׺�7��/V��e����MZ|eT(*{��Ϯ��"�،U���4��cRX& �0�.3Gٛn@~�y����Jef�.Ȅ��F�ҝdH����c8v)�_*�2Pe�F5?ܻ9�\ys6Cv.%[տm]L{�;��SP&Zo4㏽�h�nƠ5���j-v����O�5efo��l{f����h���&h�
+G/Š�˿��^�������T��{��ݚ#�q��f����$����}оAp�?7M�}z�jQ=b��1�,r��_�x@�P��\Q\`�:G�fV=�$�����6m^j,���-ħ����i+*Z��y��f�3��Ԩ��N�[Z��+�x��e�J�ή�LG�Ig��-gG�URA���uH�f~��qI�

��E����5������^��_����Ol�y�O���}��Pҋ���:$�*�Omt��y.��kߴ��ca���L$�"Ĥ��>1���L���;f;O]E�K?c��~�צn�??��'����'�0�˱<]L���%����T��$�d`җk�����$G�Y�E�������dn���L�h��Bit1���h�ɚof�6�q=���z���:C_��L������{q!J��۬|x{����x����*�J�Q(�p���l�,�G�Y�E�)�4(i����adf@r.R�?�)79 ���m����5�yy��
�ڟcXhq���;N���SՇ����XL�+�}��%��.؉�V�)uZ��1��PɄ�����,\Ab�0�J�e?����`f���S~�䑝�0kj[?H�=�k\Ģg��`����Sc�hx�V�����q-É�X0��p�X��А�ؙ{׋� '��c3M��[������b��s����ذ���8ؾ�8hd3������`�W��c�7����Q�je��5��r����#㵌�c��")7���br�2��	b��9��	�e�){999�A�_����YFDL2�� �j���a�fٖV��U���9,�q���µ�,�Cک�tk���ա6����7��\��q8b�\Y$ Q�qwq*�1nJ���'�NYu�����1?��Z����Ob�|�Dh��Ii��	ǁ���^�����iU[�+�6D���s�
0s�~|�b��=�0G��;��������3(��%"�(3�4��	Y\AR?Z��Ч�E@zB�����o,�O�'Z�v���޳�G��+E˺�mT����Cê�������x��u���q��
�$�+�S���(��fv���1S�B2��Pqsv2���HZAC����C���a���b�߷���$ڈ���ݧo���\�*ڸ��!u�@Ԡ*<ݬ3ҽ,�Ҳ������� �#Ƭ�2�\�/f7E��;���LQ`�#�k�\Mh�3�-�Y�6���Ğ��c}�Y����x~h{����c���5��=�Д����Ԯ~�CT%�
����2���q�Q��c�y�G�Y�e� ��bg��mnOb��3��Hi���)-v\AҤ�ix��=���B����UM��o+�;*1��'!<&	a���>2�&���������_C��+�~U_h��[��>X�S3����:U��$S����9��KYW#q@b��7�J��0 �r���Q5��˿`d�Fx}lgխO2����8�7�y��i�iDL
.E��^.Qx2�z���e�� ���}��?!�!
E4�O/hs��~�,�|LG81�
	H7M��T��M�s�ppAPA�.Ǽ�4{ekL|*�x�;}�}�Y��w�{6Ŕ����9Z���(B	�BkcҲrE��͌l�^Zf�S�J5���;�������_ oW������Wwx��ww�����_�k�d:��K�b��0��pĘjX$ ]K0^���R��=���������T�̀�,�����[C�F~�x�����ۈu?=�;M	�
n�`������bש�`:T�����81V
�$���L��	����5'ÅlB�?�.~9 ��d�W�LpPvq���Q��O�u�o��PUp����u�q�����Z�6(���`d�=Q�HYK8czg����a�1���U�"=`���0�s�m0��d��xG��W��h�1�iY(�I������������.EU�A5m`�m?qE����t��c�d��eR�](�df*�G�2#���vtG���/����_��x`�G����|R=[�¤Amį�6��Y�����/�G���e*Hɖ� �9��2�"��"3Ӭ}�"�=�)�LY���e����1�Oh�]��L_h@ů�N���p%.�p8bL�,�n��V��Xii`�D����݋X�@�	$���v]�J��6��_�bx熘л9��Ӷ�Q7�㺣X��`�%�S=ˌ����ɽ�K���S1I����θi焊Ee�ԓ6�5� r��.�����1��Δ�'L�h�Â���AU��z7ŘnMxB��Јs�p�i�>	fc81�	�v�Z��~�3$���D��VF�,3����0v���Ui�([LO�c.^S��BU��~�&�!`T�F�߶.�:�>���`���E���pĘfX, ��o4 5���
F�v13 ��p@bw�=�(<�Q��8d�^T�e�@��	����e��⠍U��'��unR�vv`�Ac�����?�h��0�&������#�4�r�h�s�kWQ�{�a�L�?1���{HM5���:{#G��{4��X;*M6���J�����[O����ѹ��X������G�E ZcF4��1G�i�E[�iQ'@�sv�w���6@�����Ӡ�?��^���O�Ӛr��ld���$>%߮>$
�ݛ�D�A#ë�*[3�n�	t��FQ6��ٝ͜81�Im�3�V�Jb�x�`�l{Gq��I�!�"(hLG(|�0o��n7e�G-j�|n�cJ�E;���{o�5ѫemtjT�G�����q8t!�N\ƺC���=q8bL�,���e����.}�qӚ�&���{�RR$vM��3o��a�돚q@b��rl2~Z�,��!����Cêh� ����4v�V$�f�0t�b�q�R�hye�T��4�$r�pQg, 5��, ����R�����NE��-�%`Za溴k��wT6bٔ�lN]�c�B-�t���80Q@
5�u��~��b������� ��aŁ("&��	�#�4Ϣ���.�q�Rӱ���wpR�}��^w7upt���!�؅����`�b�� " JH+�!q�u��������ۚ����ϼ���άw�3�w�������%A*��03?�B�2�_�u�#��`axݟ^��b�@}Ti��0jq1-7K�^�h\+T�R�!h -u#�P7*����l>��#�Rq�l�ă	�C��JX�잲�b��i.�꧰����n�rlE�Ͻ����vUnӣE����u�H��NNfAb������ֶ�Д0o�Cg�-��c��-(�f��5�� -�� ��a�b։���x�ۘ��d�#)#W�{�IΔ�l�M��,�K��FVX��$H�~�����I�g�x��(*H��CQI)<����M�"m;r����*R-$*�\Xxz�qbRR,{��[��l�*f�-V��2�P�oZ�8�{��"��A����@�����.p����ګ�vu��é�r��aP�^Y���_�o�bT��a
E��b�����]tki�O�H���0;"5�Q�c� �!}�t���Mm��f�s`{�ft(l��q8X���P�B��6E�ޚ���cXf���� �q�9�0K*�aֆ�uon����3H�06
��8$*���T)ɚ~H��av���3��`�����?�#����a��#�qX��]M
�U���.�:d�qV�D#?��:NT4H�b<��\P庂�^��o-U���	�0cc9JTQ�"X�FE�����s�i��Ҩ��ul`� �i=�OM��M0��4H�Y$��#b��q��
*�ܨf����cA�/�aF9�ʑe������^� ;�Z�_���:��J�T�����E�#J��Z$H�"9����޻<�q�ú�/�;52��(��/�?b��X��GW�C+sͣ@�B��}�"Hk��3IT��*�����mG->儜s�A�R�4������q.\�����׷���:50�͊'�D�0c�)G.��!Gc��"H�����Y�I飺5�J�('d�^N�g�Μ��8��ѡ���@�%���:|�����0���^�0c�.GQ<a�jDA"(�Θ j_��H�ʷ�8������,��Q`Qp�Ry�o�1���$��_]!I�0�gS���a�.��0S�T���1Lu�� ��y����h�ȮM��;->N��;f��aR��v@�W�����rͨ��Jb43���o�>-�n�v�i��0�T#,GL5�������Ǌ+��w�ɶoL�4	7�t��/"���j�������Ѳnd���yS���*��:OKJ~K'C�;�Łq0
��=�ٷ�\��z4���mt�ջN�a��FX��j�o���ѣſG�777|�嗲����7߼����;&N�����q�~���jAjX#���`B���It��l��x ��*�M����T��		��|���pk�fF�I�)�����a��&X�`�����<x�`��W�^��<v�X<��(��?���� ���޸��=ܪ��֞�0e�:���QPܙsʲY$��)�U+��� $'�����_\Bq�V�� ��Ÿd-�xE��1�0��r�������L!wrq�^�>>>�޽;V�ZFeAʗ}�m;�q=���N9S�oFn�e�"�"����Ĝ���T(ԮN0v߰�01ݵ�i�(� �-�Oߧ��m���k��a��X�'������{�O�>,HWPU���W�5*H�^�P[�X�ͪc��cs૳�DG킃I���1ZWj��n�K���^�iI(�L�����m�>���R�0è��D�Y���s$HL9����E~�U�#���ٲ(,��D�����Z��8qh�B�M���b�B����k\�۵}��%I������8�B��x��� �a�a9b��cǎ�ܹs�Y����Z�j���`i�d���Q��Q?ߺ�w���x��~����;�:��0&���X�
�:yh���A���O[������$]���$ 8�dI�<���m�8Ò��7Jf�a,��qRh�{���V��-Zg�Z��Ч���h��G��[-HE��7Z�2i
���c'PHݱc@Y�Żأ���.�g:I�h&	U��޻"�|a.��0�2,G�ѲeK�]�V��ժU��sfǂTM���] �Λ�NZ����^cE��ğ��X����������;�B#�,U��{]\6��X���2#�����&o���s�a��D��2ԭYm�F���4l;r�s�x��!�Sm�5/���nW#'�'Ft�Z���C�a����7�;rh��6�蓩FΞ���7�K8�hM��$��z�3^�cŎŅ�a�Q;�� _O���H�os��� �w��f�iРjԨ���[īM�N'f��M��V���1ݛb��CV/��$铔�-�	�mUH���	���\�P�X�9��y�X�^cH�&��d�����aF.�OX���V����k��[���V�a��f�fϞg�ZK����6�����,��� �ZA"��ŢO�%��;k�N�?���@3I�ܭk��LRR���{=� �_̄$�I�\>�80�>�5�:�=�ʎc����_7*�^Hǻ�T��U�H���������GK�Ʈ/�a��}��k[O��ݚ��(R5���H���E��9Z�@�B����vi��;��v4�Ը1K��@�O��z7���n��yfڌ������F��\�Sm��vx ��Fi����;<�*��t:��!+�g�3���Й�J�3�A�V����Q�x�<7�ALnjS���Ş�V�x�I�u���׽�!q��_���*W2�e�+�@}��k�mDu���%�FRy�b�����믿гgO0������"7�����Y�7&�²��Ġ�2]�q_xg���V����C��g����T#))�حd�6 �F[������8I�A�딼�^?&��D�vq�d�~H���9��ێ��aI�������]�JI�.xtx{L��j�㹱]*�����X��ؙy��b�46r��߇���0Le�]�L�E
���4��Vs�g�
n��ӭ��*,dI�NH��b���J_���P�:��x�V�f��[�Jдv^��/�Z֑e���zH�b������߯ރ���0vI��p�G��>�H�o}P��T�nd�ݿ5n��\�{���]�Sg�(�n���uI�ć�Mи(���YaI�F�nK�HRt�GC�h�	�������a��@�G	I�������^�p�Jw��":�o���h�'�X�-�΁qh�H����� �އ���盛�M\�[��H+�������ڈ�Q�b���&�&4�4{�^qr0�ǏD�ǿ��O�w@���_�cݎH� 5��jA�'��30�-۴�Kq��-ЫC��}�yg�}=1��UKޥ;���~�H�c�_�>�P8��b����(������]�Z�F�<� �a��&�xg��ܹ1B��N<���G�ŋk)и`|D7����e%��
7�LR����B���c��:��%�\�	�Y�i�ǘ��LI*N'�7{Dԅ/�����;���}.�B��6,G��1�����,����p��X>�3�`3���]�W܀Oht��u����iE%�+����;an�F�6�	YT���"#����:zȱr��
�݃�Lh' ��Z?���=�n<�Bjf,����w��W�U0�}}|��0Ѽ�������FlP�*�.�;���\>���]�v�S���)�޽�:، ���������@��߽�/�z�,�]���BZ፴���O�Ő�׮-�4��,��Ǐ�����W���|7 �ڴ$X#Iq�"���L�����"��r���{e\K~Q	68��."5+)�y(,�<��xx?/���^-c`<tt@�8L����b�a��#.��X�]w݅���
-[�Ċ+0u�T0�`S�D<��Z�z��	�C;6�͝a�֣��ӀF�\�g3�oH+�������9���b�������\�\<1"�Γ�(��6=��c|���&m�b�~,_����F�ۺW�Mjv>ޘ�ii�9����v�-�RUPI�����{�0c26"Gr]��lpn�?�}��	��='.�����vF��p�}��D�9x'�9��2&e�eb��z%�� 5j�Y��啗�1�6C뎛�{���`�$EB��h�$M{j���ݮ��/�X mv�h���^��/�w�6�O�=ӗZ�?l���b!A�H��En��������9$��0c6 Gr]��-ļ���������H�0�alN���ތQݚ-��%�>?���E%��n���E��s
�A�ii@����/#Ь�ŋ��d,�Fr42�'���p��I�H��1���6�đ�{3\���2��)�F�j�`D����9��	�.F^��H�aݾ���m�O��u����ĳc�`�W��8$�~��jǛ��-�.=��Y��*�@7|�[��l>�o���IA��S64�*��h [��a�ţ��T�/)BT֪ŹI��\��'e�5"r��B��yW��$I:I�`�$ՌƗ��m��O�M?\��S.I4� K�d_CwKJ�p��d��
R��1��X������y{��R���,0�ݠZ��j��2 �U�I��*�@a��Lb��ߋ�֗^.�Wy�@9��(�M
A���+r��A�7��K�5�$)[�G��ɶO1B�M3��qݺ\�Z� �5�tI�]�j�1<����("��N]�C�9�</�I�T����E�ݍhr2�+���������\�ݪ=�7�����BL�����ESn��U����K�ׁaF�A�������<�~�^��s?�s
nw)=u"*�N\L�0�a��D<��*�������r�#���F��^K�+o�$�&Q9p*�@�I�� 8$F$�RW*�E/FG��i73�"�$GI�tI�$�3y�IyG��Y+�q�a���堌�a�$Ս
Ց�����	3ơ3)�⏝xbDG��wi��X�d���H�����a⠶V]�\�oV�ƚ�'M:7����5��oW��0�aӂ��W��>X��o���3��H�'��p���'o�~Y2�����Ç�E�����lfP���g�*s������=��b�]>�($I�ە]}����q����r�ۑ$��R`�$uiZ�ຝ�/�\J6�`��q�����\(":��b�ϱ`����(4��놻Ftm,�f�Zw������*B��!7�XQ����6a�?��a�iA"v�{�/�*���A�HԬ�w~��=��[y|���:��$W	��'�(Q���`ǭ�Y\\.FT�T����0������^$I���$�\�Z7���_�Ǥ�f��7f��8U�_� �I�Ϻ!V�8���/�'#�4һ�]�h$�a�C%9��ջ0�W��Y~�B9�[�h��-��ه��c���A2Wen@�բf͚�������4|�~�HUs322p��%i�$�I�����xO�>�cѶ~��m�����㡏���=������0'qj�*t�"Q�������� �!���_D�����ѷ.�k�b�Le�]�%)Ϋ?|^��&�l��?"9ͼ��rI�I�R�vb��:	jR� �t�0c6*�Ս�o�����+Ev��/��.�,GL�j��ȑ#1p�@t��	�&VH����_�����cɒ%HHH ���2��@�v�޻�>�F�ӽ)R��������������7�]Q�fYΜΞBC��S��Y%��HIRSe�J��p�1�ѯ�����ƒ��#����Ղ���}K��+���:��|JH6z�F5C�+�ށ�$��lV@�0D�h�O0�TB��B�sTta��EH�(A˖-��o`Ȑ!b��\���a��2c��\����
v��	�z�B��3�Y�hì������C�E9⏖�-��Hw����>x7e'���X\tˈ��I�����TRB�(ʥ(C���Hr�Ą����
�	���o�ߊ�`�~�GO_��-��B��t����1T=����j�ڰF>~d�֏?Ӷ���m��ZcU��M����ť���yqQ�	6UH4X��2��8$�Q��D�:p�-ہ?���4�b�Ic���z�'O�H��A�x45`� |���x��PX�r_���L�Qo�I7w0i�W��!�gRM9�Э'��c�W�%w5�r�xP�7Z���+Ѭ=z{W�����K��L��W��!B��\M��1_/w,~u��2��H��ŝ/|�����h
%ёS�$y{�����,�4����>��a���w8v޲YQ:�eI��Z�)���9��zx��D-������㋻�Q�M`�Ѭv8:7��c�RU+��8��8o�ҥ�ٳ�"�'Qz���/f�R�7c_�D�9w�4X��N�`
3���|E�)�k�48�4y;�+�s�T�fg*fhH�||�[h���S~i��R.IP^^���nC5�6�{ş4��A-P���񮇛+JBѬ�iM KJ/�g���s�C�LEHR���������^��)�����Տ�N�* ���J�
��;e�&��H� y�����C�P�Ƶ�����&���删�ä����X��$�Y�[�ed9puuŲe�н��ʹ�G�m�6\�x���ǢZ��;"66V�6�˴b�
q��ý���$�Gz�����&\�<wn~}>68#������1��T�!<�un�j� q�(�p-�4K�$Q�oz�6-�3-���������f��ц*������x���RP���M�uD���B�8xZ���)����J��7â�cp]���uƠ����AEnA1��|j���T�����9��C��5�;r��|:*�,��k�ҍ�vqb�&�T����Ĭ+�X
�铣��||��"4���+�ޠA<��C���{+wh׮�M��I�&�ٱ;A"�J���aݻw"��ۤ��}nn��+6<+��)�h�Nps��[S�٤��(�]�8'h�]�Ӄ��+����2�BEf-٤���T�]p�p���bQd�F��#���^b��*��(T���XLHFצ����ٲ��D�[{53�^ΪaL5��]���9z�U�w`4�mx��q��x��>�rkw���h{�L�Uo�Vx ⢂q�|*.��q|�����OVz����3f�9b�~�?.���g�᧟~Rt->� �y�1#��إ Rs0��������t7���#&��6w����}\��D�=j��C��y>J�Lrbvycrh<x)v�pX��-����N�%+�2���� H/���"��D�Ij�:UPUO�3Up`����������,�єbBߖz�D	�q��C��j���3�?��'��bp�6ڱ���4�au�M-Ų��y~G�R3���>f<�#�67�Ϝu���7kDY�q4hP��-�֭��P:s�}Q^�֭[ѢE��ϻ��c�С���/��ح � ��<����~�fqg�N|J1=�)f�������sJ�%sik8�������>1�oR�<� _O,�$���M�Й���o(��6M���*{Q/��$!@�!~z��I;�U��O|C��Ɏ�W�>�:���4�����pW�V�v�E�M�}���ip��#�D c�؈]�3h	\'Dg��D��\:5�!�Č\��ffK�����C�|���{t� )#��o�PNЍPȝrTA^^^x������C��,Hv��mG1��PL����|�`D��[{_�.x&,_6��ps�Y�kcT�$�xᝠf��/�e��lP)��HӪ�I��m�ۿ��u��:�bU$�	�D/#}4�WW���:tF��L�C�*7:���k�]O�9Z으b���SF��QCPƎ�A9���S����ap�"��KӚf:2�ώ邧Fv�I4�D�K�Ծ���Y�����Jϭ[�N��P�����&�v/H��?��$̑$:AQ_�MR��n~�7�3>�D�9I��p��12�n�"�>h�B��Q�_�ƭ4�PA�t�����ǂ_��$I��ۖ��G0�sS��I�W��4p�}�LÆ�	`j�`H�(�s�1���8yI�>hԻ�FVYj��;o�,��l\���BH�o-k���1=��y�
*lss�Fb��/�)-�x�E�_;�1�z��'.z>�%%�-J���uq��2����D�$щ���Th����R^����ƭQ=Ф(�dĐ��P���}p��K���ѯ.��|4)<l���Uޙ���!����*q�L�r����ኌ=��+5󤦞J�Ȱ�+��9���l.�h,�|�o����0Ƅ�a���"G���ʧ{`p[<=���<ӗg��&����э�L�3_��s�¸��pπ�"��\��yFB:o�A|+�R����Ȇ�%3���~DTPa͚5��U�V��KI����#�0�DT�̙#IC:4��7oǘ��Rq�G �슸�l<�ucs��4����#�h�$F%���o�"l����-�/Gh�咔�M�2��݇��	�����qX������op���qL�|�N��
���WO�c�;`�_�j�I�2aF�>ϭ�EbD��۳���e�����J{Ŏ��Zr����+v��fW'J�40���C7�����ڊ�4����[9䥗^av�/�wtʔ)&��p(A"H�J���㺚�
���]��_q��:}4N��cRX{���Ob\��,̓3��;Z��zX�cz�!�x~l<3�t�&H����i��I��I�����\l�w�[�Oq\7�Ԧ�u�Q��ԏ	F�u0�s#�pl���"$��y���<k�;D�p�c{�ͻz�ʣTD��o#�vwCT�/�����J;�_�k?n c�8����g�By�w�k��}[�Pds��Z��P�ֲ�2i8�ߍc�4�|L�8YY�U�����̙3EźY�|9��$b�/[�Z!ޙ����Pr��w'�;�j&�^p������R��ܚ}
�r���9�t��?�����zHӚ�&a�>�5yx��&�A3F4sd�U�ՔK���_���Ǡ Q^-rA!N_<>C;60i{����p�#��-h^'��LڞB�h��۠���n�`w8�]姾5o�]��;5�}۠]�h0���:u
����yt-#G�D۶m��ob�ܹ(,,4k�T�{Ĉx��WѸq�J�-[�C���qHA"�2LI�e�k*n�x��~��*�|�\�^2T�z�g�X�m��I1�(	�˲�k�t��O���S�<���K�f���Sëll��c�S1���"��lH�B���_�����_��{,����L�#��R���]�1�����/���o6Y��f��z���d�'��k�^E�,��ۛ8���i����/FF��+�=������:u���o����ӱq�Fl۶M4v54������h��ǣG��_799�>�($��d���G���B�37ϸ��]�}��6yZW��
?�'ã(��rл4}�2Ѭ,��#��M���;
�%1��j^x�P��c�ۛ���G��֩����
I�9ܮ��?,݌Go�	Jc�1�]��C�?��'��4$e_��%�2��l���L�nd��$L�l%^�>�w�i�{����:#Ð�P�ؕ+W�-� B��ə�2dΞ=����>Ig�3E2~���u
���W~X�Oہj!8E�$m+�`��?�Bm���I��s�R���0�@��Mu��~�`�����{��V���ώ@˺�0���/V�SN����+�de��/��}�{�Cốy��碒��\2�@�B���%����nT�"ǡ����Z������Ȉ��ѵ��'�+>[�}Z������5X��qn�`Bǎ1o�<��v�¸q�p��	0�8� {O&b��s0�[6�4�z�Jw�}����eJ!I�.-���r�)w��"�
bʊ�B��&�|�.+D��s�#ɔ�L�y�Z\p��o�w��	�"� pT�W�%<0�^�~^��:Q[E-���?�$��$�X�Р��l�Y�G���,�zT��0��۔����kv�º��q{�"߂J�b��DSM.�m���>�k��-4�D3J��n� _O0̵$$$�k׮x�����/��ȕ�yO�:���~HΌm�l�tb&N�+$����������GK�ƴ�[T�3�	����@��@��7��+�.Ң�E:)�h���9ʤ��,�/{z�r@��U�s��
[ C�����G�:�f��f�h�h�B�*$�f�䒤f��mC:�Fz#�*�/�~?�ݏ�}[��#��z�H�g�����v�XZՋa�T�����&�r���`B2��K����p��&X�L"!)SD����&����A˺��ǀJ{��"�h����BϞ=i^�Iц�x�b��[��Y�����P��7�����2����p�t⢼�;ԝ�4&I�(�D�Ds��Bs���.*�.'�@�f�l�)zu|QZ���A�F�w�4rJ�"�:�SD��e�W��:Q�x~�������F���+1��mb�KM<���Q����ɸ��ƹ��{Z���,>+t�<,��^��5��t��7}��3��\��#�),.��u�BU�V�y;��1�QTT���hԨ�X��Cppp�<u:�fff�ҥK8v�>,�c�Ʃ�����L�Oޒ��n�f��k���Y(
%�#��P�rI�.6��Vn��AG_� �;�Wc{6��{"4���g��p��E8rV�>XI�&-I�{Z�f˞�\�s��ꡑѥ1ָ��Jw�W�����~O�0�9е�f�ia��#����Ҳ2�k+�wr�'s��G������
>�u�:+f�,�"C����y/�[�3���(��6=IqI���g/ٸ$Q�
���ļ��k�p��f������B"$�G��BSZ
�4X���"���H4�)����?��Z;��1���k�!�P'2P|~(��c2�UX�d�B�*���r��l`%qZA"�9v�'���-]�\(��;z`�M-1}�6��� �F䰐$Ѡ��y%�f��Y$�[JjV>&}�+wVo�!I$�E�K��}�yR:�
aN4c&G�d�5y򖎈
���)�!}���8c{4�g���3ܺ5�����Q�0f�#y�����٫����0��ԂDЬ�},ÊN�&�>�W<�����Gu�9�'��'I��VP}^��vx ����jn�~��}.�d�-�$�,����jF�\b:Vo9 $�^��/��e��!Ϡ��䩔zE�<�V����M[$*�1�ä�K̒h?9�#�~)'��Hv��c�(�gߖ�K���_�7�0���T��[�`ۑ��n�0Q��h�>��<�>�u��R
5%I�_�gU��D��g�t���ͬ�U |�ǿ�͊]6W2�\��%I2�GH�/~z�!�iR��sGN]Đ�f ;��>H� bt�}�o�>�7&�Ϗ����`ԍ���y�����]����x�۳r1����/EIL�WV���_�ƛ?mDD�����7�0Ut��sD)�G����q�L.K{#���<��LU.JT�X	��$y���=�$I�p��2M AbD����hj����J�#�,W����Á�h
��l�����Ѹn4��/�~����� F#}n.KR��XW!�M�(��+�0��>�\�z���v��8�Տ	ƈ΍�(m�E!��>F��sq(!�O\������d��f���q.���NJJ�*t*����pM�1�I���1���d���ό��߉y -ۼ2�Ơ��.X��+/Iڼ��$$��.���B1��*t��b���ढ
����$T-I=��ϛ��Ȩ 	���\�jzVHR�����=�lg �(K��7v~r�ȋ�\�	]eT���r/��	m�$2FT��X���+"$����+v��5��[E�ۃJs���o��)S�X����p���"?��Ն`A2 Ug�8�7�Z�<����W�� R:�>��XV�:��&Z�%I��d�7�Q��ݛ�[���M�y��${B(I���� _���D�Q]�/�:W
�4�k��:G�r{�0�����t�ܰ?A���ǵK�Z"����d;ǕU�I�Q�P�|x �Տ�u�t�{���xvtQ���e;D���_|ļy��~���7~��7������X�v-�z�-l޼��� aӁ3���xhH<��IT���~m뉅B�n=&��A��d5W$�¦P��$�f�p;j>j-�=�[c�������b��$L�b�x�W�$�R�)��8�P���l��%0Lu@ax�;5�=RbV����^{ݝ{:�>��((��0��r����F��!���������X�����`B2�Z���;�8q;v�0�u�?���#�����_��{L4�e�aA2j.����X��޻��K�c-t߷�X��悍�� �5M8��nPZ�49�$I��L��th Jj__��eo�t���0(Ic�(5����.��wn�s)Yx��`�I�h�=}p�����I�0�x�v<��
y�N����K�,A||<.^�h���ԩ�����u��ŠA�P\���P��mS���Wn�.Mkɲ_*�@%�i9y1��ŖC���Y$g�90�j�$�L���J���(�I2A��֏Fצ5ѵY-thOy���\���w㣥#+ϱ�I��@����G�U������cAR'�� nh�U����a"���0DGGI�ѣ

LK#��x@�:�Y��Op����aA����/bث?K�Z�Y�\�Dԋ�]�Z�����&��$K�4�0�ԷG�$�|�J�� I"�����[�E��]$)�ب|���rU!F���C����J�^�$�ޑcV�F���2!���02�r���vf���>��-
-�������1a~�5�Fᴉ}�~)ڄa*�$
����[M�~���"��$h���p���E3I�-ªU��� Y	��W�
Qz�����TP?&D,w_���\����yi��~��I7��.�HR�zѨ_;Ƣ~lH�5N<%㳉��R|�z�(���bt-咤�ڗ�a�kf�\��ˍk�Јr8�Q����{�.)3�V���mGq�iC�f�Mm�at�&hWua�hSa�#�R�,�8�ƍñc���k���=�-͛7��ŋQ���i#S�NeA�,�(�q�(���خhQW���T����k_�|NAQ�4I˿�8�	:5;�y�Ȼxy9y��1=��������ye�@��04����"�06R��6b������	�h�˒����r���ٵ�E=�Ԯ�ǘ��ʑ��<0@����ҍ�����] �n|�|�X���[w�F�X��wW|��0�~v6򋔍al�C�����k_?|��Wq��Q����&�����ׯ���'�YA�֭Ųg�83,H2B%�ii�0w��R�PRz&����<��Fʎ� O���<i�/Dv^<�ݮJ=�����NM(7뇵�1w�~d8y�<�$]7ʋKJ�}�IyF�n���r7��-��0�A�t^���j�4kFti,�<h.jT�c����9zhH;4�bp=��m�"l=|��c�>�<����O��hp;jJ���0m>�evFRSSŌі-[��}�����s�Ήu�r��)|���x��{�ĉ����]�����=��ξ-ѸV(l�!Z��б%h�h�֣�����.G)tG�?��*�)9�#�խCL�6�^Cq�S�_�9�H��;�?�? ���?��a���Y%���fkop=U�������ČQV����nĹ�l�d����]���oT4 �<,��_�<=[�1y��ǾƩKp$�Ҙ1c��ￋR�Pe��K��s��8~����[�`A%A��;{��[:�ۺ��}��?6�7&�������K�z�bVid�ƲWps4��M�k���y�	�����؁L~MBR&&���
	���Y�t� ��*q��
8�cz4Ex����/~���rt-��<*�WT�Շ���N��`����E���uχ��`�ʕB�M����HX��)��J�=�(��f�Ǡ�8Q��O�X�(��I��]'�|�	�R��,�d�>�{���	4m����?�}��(�F�˞�D�čl;b^��&Y���(���q{o�w�)B�$FI�Y�E̔
m��,H��_|���8L�<���ccc�b�
Q�;;;��~JJ*糹��|$����7%~vl\CT��׶.ְ�0<5�ӿ�'`��SX��.�s�s).�,�@n$���Y�:1�x��[�#��ɯ�-���|��\Ʊ���/����6���h�Y�i���'����ߺR�W��a9B��W�9�o�ۤ�{�p��g��b�Q#�_T����0��3�<�����t-�Z�!xT�;?��P̨���ବ,8;,H��e�Haiy��"^�_�8�m+������tZ��\���;�:��K�[����Kf���E�Gn틧�/7�^C=>��ی/����qL��JrsG�hT#T4Ϧ��K��U��Y�y��yl8�D�*�Q�S��	(�Ck�rݱsi����L���5*���褋�wމ����u}9�nݺ�F�C�EQ���7��0'��QaA�!(1�/i���F5C�	����o��� ����}$;��?Ҳ�B2J8s@N���s����E%��x���Ӻqm|���hgzձ�[�����B�m'	3�C�q�/�)����˓_��+�׋��������6N��UZ�F\GC����G
R�z<�� ���1b6n܈-�oh|�M7a�5j���F�Q�SO=U�yڗ�Âd��y*V@��5��s��ވ'Yj-�#Q+"��Pݤg��RJN�IƎC���>�Pi;MPt��`�J��yn6&��k��Tb��Ǳ�\6��_oL�&��a�n�$�e㥙�����Q���(1�ak�)(Ʒ+���fЩ9��N���22�rtk.����Ɏc�src��0��4[�nE�Z��[G3HT�n������o���Θ1C��]Kzz:֮]g�G6v�����X�%4��!~����i�?G�"��S$CS�$z�p3�O��WX������\\L���dZ2�>�<gzGoMF
��$+t���~��Io_�I�,����wm�w'�Ct�iX�Ɵ�l+^�t1�s�+�iʤ��^�.D�$W>�0�Ae�i�V	�,�$Ku"x0�*ʑN�2�#".�pj®&ǫ8yb���߿?6mڄ���g�)��Μ9�Fdd$��>t�޽�~>��C:w�I�G5@jV�X��J2i{���hĬ=R�HYi	tɗ�cY�r	%,I*A�D���랎�z�Sc0�gk�wu�l�����;QiI�F���P�$F~�W��K��oێ�'��]�3FPY�t�y���0 ��(1ü|;k�\O�J��q�<e�8AAAb�Gg �Jv��Y�Fl{-u���T�vڴi`X��:��%0�T��Y��$��/0
��S>�tE�+^y�f����{/.)�Gs����+ſ�+�>7$I�����y�87��+r����59�1�j�#��G�����ǹŨ4���*{�vZJl��"�<XT�3Į]�зo_�ɜ~Fiii?~�޲���Wb�]�$I*S�īMOFK��H�T�f>xx :��g����O���'��h.6:w��ȘH<���W�9%c.Ԝs|��pSKQʘQ �#��L��/*Q����7�~��8Jv�
��Q7��\��Ín�{�nt��Q�5k����4�4d��<yL9,H�uh\�%I�v�<�DA�$�D �G������N�4��ɉ�_���K0{�f��S�F�|��ՙ������v��O8y)c
ݚ��E��ׇ��)eF�`9����0s}3�>��7�lR�� ��32Br��,}^a�$%%a���&m{��)����^��?����y����/1u�T���:,HL%H�t�$!-QIJBY0K��tnR3��1�0��7���3�Ju���}C+��E���q�*�`�j?������>[GϦ���v�����x�֞�E������}�b7�*�\*�Qˑ�J�'��P蝒��g����ܜ[6*���z�M�>]<R��ŋ1g�����w�b���*�~�mQ��iӦ���Eff&:�-[��-�Ͱ 1�puSG�t�$˝N���oL��{���Ĕ�H�����j���ٵm�Ϸ�3|ag��-c1�őWƩ?�.�����v���i%^7�Kcx�[~��-��b��8q1L9R>2�й\���b�%ړ2r%A�,����%��������QSFlT����~Z��P�X*�@c,H�a*$��1t
K�$bT��%�rFti����#r8L��H��u#��r)��-OJ��<_��RR��וQ���u�TM��7'��(	�/&�g�k�z����{�d�QQY�1��rD3Gv,G5m���?�ٲn��KP�}D��f�����7%ذ1�S5��$��cI�Jd�~?�mS���NHƓo����W.��F����K�CФ��|�57֔���b,�xH�5�fLDm9�Ӱ�k���^-��]�:.J5AzjT'�� Gϥ��<kj,GL� 1�qS[���;��AI�n��v���i��K��/[Eo��YYP�p�F��Tƒ�
���y*���o�%�=�(I�^������Y�Y��/\wK�Ƙ�h���AL���h��[����#�,H�i\��KbЫ$���+9I<�����&�ps�z�B������g��[���h��eIr
����>-1�gS��[�:��D�w��`�i�`37�rd1����2���ڍk��S�f�ܙKd�/f=s���t��fRa9bL��1I��D	�De%�Ԓ$Q�q�b��[ŊEu*$IT,�JG��{����Q8Zá3)�������5�YEZv�KԥiM��ߧ���~@A��� �A�vqxdX|�7�Zc
����#�DX�� a)�h&��$]�u`Ir��4�J�+�$G����b9�A�ҭGE����X	ˑ,�[�� Q����3�Y}��ԇ�������k�k����X �c,H��I
��<JJ��%�)�$]p8t��ʙ9v>?�هy +Ϻ0O�
,G��h��:�'������y��x�UVg�3#Ч�y��o��)���e�a0&�rĘ	c��J��
7��V���utФ'�,INFq�e�����-�|8FFX�d�>���o����6��ĩK��%Ą��-GP���1���XN�$�]R�0"��j�h�$G�$�f���Ʊ9����k�b��6�tX���U�qg�����!���bA��<�84��"(jS^ꢚ줸��Ȯ�����?�)�dAb����j�%��I�B#Eo&�1Ц'K�͒䈔^.Ê'Dх��(ˑb���ᑏ�c�������������E�O^JGfn�؇��?eG�5W�Ou�Yi,Gv��?;�~�L�'#��JRKq��){ ��ct�O_�S<T0�L�dIr,Υd�ǵ����������r�8�O\¤�W��G�m�J�-�#��9���zU�{�ǿ�0�r� 1�P!I"'I�È� K�`��� ���*7y��Q#"���i��&�%ɾ!^���Ͳv�)�������������(*6V@b���k����k��|J6�wj��`_���*��/ƾӉ�?��a�`Ab�$)8B�&�"Ie!Qи�GXQ�|P��@��bp�ͻ�cܠ���߲�Y��x�Ol=S��m�"0*�r�:tCj�������h��������{��ȉ����0����KF^�=�%)M��hP/&�L�%IY$a!q1$I�g�@�.��s��Ԍ\|0���t�$ۥ���o�\�[=X���3�Yx��5`���%#?B��Ō���]�TF�\���($I��	R�c�[�}HgDG�Bb:���I�YJHR`���bl����оaL��w��^U��aFxT�(���j��I�Rݎ%IY���&J2D3IrAyObȒdS���,|y4|=�k�Le�)ԈQ�#�a��%�*I�F�$Ir�z��(L�	u����t��`&(��6�7m٨��k ��
��D|4gvN��P,I��?�. �ѯqO�ֈ�ƿ��͊�H���F��r�0��u���%
W�eLb�ڳ�p�z��� 1�"�uAa�T��/�tɩ.�[���G]�zD�ojS���Ş�
�\�A�z�7���H���>!�kGb@�������v�:��$�T�{��͊�?��5����檷�rUP�]�*۸ZuX����kV'\ܴ�	������1}Fs
���_���LJH��)"����o������V㹈�Q%ܳ$���c�V*	���"�,M����/��hғ����W�����n�Z�!IT7�����/&A��-���տ�c8,G6O�ֱף��/wˆT$GT�n��cX����}���$FԖ�2�B�q�}��p�G�r|��' IR�z1z�S��\P7t1DdIrX޿��Ur�p��44���m�Ѳ���[�}'�7�셯��Ɨ�DN�:b���Q�$]��Bs���(��|�-�Gt�f>d^gvk����������|�$�L��>8��ܾ>�+��,~��x��~ݽ�"���������0��ubF���C� 1�b���lH�+�dqC���Caw�iGD��^>�Ē�PP�s�#��~L0L�Z��+2��>5����㟭�%�� (�Y5FX������Ph�R�=4�.A焒�Ȑ$�t:�|��TZ�ee:Y�u6%K4ᬭ��Ӧa9�YZ�F��4ã&#�6#Ǿ�)Y�pZ$9�f(�6�
:wO0S-�˫�)-Ii��$�C��!Y����m�Ȱx��ǩ�L�el<d�>I���r5�8���=e9�Y�^rT�9���Xy�'d��騐#y��T	ɑ��3NSm�.I�LV�G�%I}�o�����tg������e,�b]�ĺ}�1��9֩!b����aQڡ��%�m!G�,G6�,�y���(��kw��p.%��b��Z\�Z��T#���D�b!��CL��m��2O�
wԖ��p8�Ʌ�$�Z!I�I��|%)��$�B"X�!I�����Q��{��m��7k���]���J^�\e��̑k��"�#��v
�*�V@��?X��W�C~Q�Y���q��u����֬V�۶o#
8�o�F8,GL5�T?޾"�^qI*-�"I4��a<j"��uZ�4�S����.�K�FY�F���HT�`9�i��ÃC�U��=��r�f[�D�.�-T�qƃ����z|x��y�� ��利fX��@EI�H�T&f�S�(F���~W�xs��E$��C%Ii"4:e�ڼ���v,I�b���;_J̆���y��U��-�x�l�J���_1�J�t$g��s�za��9pXX���j�� I��i�ҕ=Ni1�B�h&��N�E%�X��jǫ���V>0KUG��n�.�%Im�[�0,G6OÚ!�ۦ���ۏ�ǣ�.�M�*��������o�.r���0��a��p8X����)t���mԐ$Mz�trtLI�)\�%��С�$i�s�#Kc���6ZGyF��\�X��i���%X;m���ٻ��r<Ab9bl$�� I��mv���є,I� IRYh���PI�I���)X��3��op�GK�ƅ�E�Ñ�����o<7�����Z��J��>�,G������&>��9I*I��i�d�,��B��y��DM~�xdIbl�#��m�h��/�PP\�oV�V�}|��QZ?зr�Rʍ�ժ�ȃ�{X����]T�$��,I
��Zރ%U%I*�A�M��&����ޡ��\�mƗ�Ȯ�Ҵ��u�ߙ�[�����J�m?�	}[�]ߪ^���c�� 1��$I�x_�T)4%E,Ij�R!IIҀ�T�Ci
� j�Ē�(�Ե]�h0z`9�;�3���=��&$d��El��#ƆaAbl���xTE��%I
fIR���۩!I�:���0��rd�4�i���)���dߩ$��B�K�yX�����%I'IR����ۏ$�^��k�������h��P�S��
O�@N�('��e(����SX��`9�["�|�>O�'/*\a��2r���]���y�1����:� ���6/[��TH���$�09����������j�!���ຬ<���]Eu;U$�,��b�0J�rd��y{�}>��E%ʞ�n�r����0W;���(G�h�P��U�1aAb�����*HҤ�t���s
��
�����|v~���q-�32�&&2k�W$)-�R���3�Y�a9�k�Z���-,��P$w"��9^VT�#�1���$Q�����J�).�iI:���:�z�5�����)�:6�ap��0�$1c��$%I�d�	Ό��rd�е��j��X+,���<u���Bu��Xc��is@IҥK'u�q8����Mk�]׳e��n��ګ����O\2o�W%)I��(����%IFҲ��٪oק�^�o�#����PH����;%iQ��9*!�NB�X�;���[H�t�����P�tr/�AI:p:��Qݚ����E��RP����z�� cþ�wz�L�
��F�f,I�rY��s)ʆ��4,G��V.�@�wԠ�����
���t��k���r��),H�}R��䄒�n�i�I�/�vx ���
߮ܣȱ)���=��v����\�ғD_%��$1V�r�pйK� ���p�\�*�����7�~�i�%�m�#ƎaAb�%I��]�m��N����Cgѽym��_���X/��<,�󧌪2����{�;IR0IR�*��IKD��W-dl�#��tb&��E�]צ^�j�4(�>B���:�+,���ga��1v�H�$
7�)zMQ�4h�I���~����鎅S�`��?��%y��6���^i�8q�L
o9b����rI�v
W�����q.s�`�DX��='/ad��z�umV�6T�=��єۺ\�v�)+[��bX���qt����Ր$]f*��f��#xtx{���"��S���oֈm-���n��Gueg����롓��H���$�LK�~(��r0*=_�^N�M�r���8z���aʬu&�1���n�1!���p 6	�� � 1�Z����/�F6 IS�_��^��`��@_O|��P<6���u�v��)f��f�z�ѹ1��l�`?/���j�.l؟ Y��$5����$��+-KҍPXgt�_��S���4�9<�N\D��Y�0P����x{�&E�M7���I�!�B�ݧ`s�1�p�$��Y��$��UT���_����]�ܮyl���ƛw�ƅ�����������y��!*��k����������E���(�$+4�#�ɪ I4c%��%�:��s��������	��I�0�F���Š�W�_���)��߶�}��]�䈎�t�6ɔD�Y�ճE�hQ[�Ԫ�~����q0X��D�Q�A�p�+��nIzw�4����q&mO�w����yk!�J.C)(�$�%=I��)��cI��s�BlT�u��n<�i�7[�oJF�����TE��j��ȩ�n���D�볞�7��s��L���}��@��ky������f��̭�r�тaԀ�q\h&�LW^XAAlA����ӗ���7�,IrA3Xw��Yy�JQ!I4�Ē�>�9���"��nT�M��������I�Y��rd+���U;O��zz��,Ϣ�Ǣ��?��w�����l�L=A�r޺�7��;��H�.I��y�+��$ơ���ST�$����()-�����xpp;ŏGR���]�(���	QH!-�����IJ眤�s2Q,r��-ca��9-���/�Ԧ��^sD��>~d����E���6[�*�Ը&���H�R�2�▘�쵅1����+ Ă�8<jI�a_�j�$*ڰa_޾���˯R��W����ET����TR!I�?#?..6*�,GN͎~�l���6Հ��Vܠ2k���(?c_%�!G*U�+������ܰ 1NI�.=Y4{U�$4����� �,��}��:L�4�'�����%�@I��d�����ϖ��E��HXa�>�Ja���0B2���kv����ɩgzfzz:ujno�PU]�Vu���=��]5}����;�C=�
Gw�#�/����>n|��X������on��v����F�!i2����r;!��bѐ���F��pDQ�V���ׅ�.[w�?�En��A����}���V>{��28�鼖q8�ͣx��� $�N�,}�wH������ǵ�քWܰ=�����ͫ.z�т���]����W1����Z*��d�f���g�tdk��?�����ǡ�� �V8"153~�w�2|�7_W�{�t��;5X��?���������F����S�ß�F����f��&! �\�,$-����G�6�k6��+��B�����9_|��#�'NO�C��K#�K�ِt��R�w}<$��j,��u�/��RU��ý�����;>1M8�i��:~��~�g^~��	-ɞ������}yQϽo�dxŻ>�v���\`�:.�{������ՄpD�h>ś���bgz*��T*�Л�>�j���Xu���K���f�IH�)��R�!����\���8�8p���B�7��z�L��GO��b����S�G��2��рpD}	H4�����7���?Q���|w_ }��t�p�M�\����Ŏ���Z!i��(C<\;>�J��(��:�hZgCҁbHJ�<��q�&WI�����ǂ����RH�Z����	Gpn�MJ@���o����?��t������RH�?rg��CCR8r@�w)��܄#���DS��r�������KH����p�\�zH��IBR�ͽ�-uI��܄#��ws���!)::�nHʟ8v�0Y!)��4�����8��;�k���B8�s�@@�����I���|gO }�}C��釤��!)�I*��64��m���?}�?
�3��k��t���C"ː�-}��q6$�?�*-�ÝK��	I*�pTE�3��#����7st������䉐t����}�bH�/v�Cgw }������\R��1.�H��Hx��I����$x��������CR~���=IBR&bH��2��釤�Bu;!�1Gpn�<���?�rG�0#$-+����vH��ϝ�n�X�
Iu%��	GpN�O��=IY����n��+��bH�/v`�⛞RH�z�y  =#IDAT�_����E8�s��$��|>���;R�($ec��/�
7$���%77���8��Ȑp�&�	Hp1IH���r3ө�TI��\����w�-�IH:���NHʄp�&�E	HP�bH�/��K���������BRFbH��R�O���:�y!)3���pe��\�!i���9[�!��g"焤�Gpn��M@�J,��#Bn6�ӹcH�/��y!)1$ř����N1$兤tGpn�TD@�J�B����O=$�!)I���>;��UH�����@Gpn�(�����Z����Ly���E;�5[+����Rg�CȢCR����L�\�S��\�_�Y
�,B,�>1~v�W�/�#vt����&O����G�:L���d����r�,�qA�K��^��+ P�������ձ�H  Te��=�w�XN$  ��	�Sg,'  @B@  HH   		   !   $$  ���  ��   T�m�Bxp�he_4;ѐ��i*={�P-~�333r'*lU�����#,ks�!�M�g%����|��%��hxӓ!w�x�/�֟zYx�M;43=(��w<�x�@�_;�G���\H�|��7?�&���@F�&C~�`��ߩ����;,K�3!wd�?#�|KK�^r{'4�ɉ�?v(K�O��9���Y*��.G�!i>�`鹋ALH�P[{�+^�|���cGC��,��T�p�o	��2
G%-~&@@��-������5��$�m��T�%�"$����	˂p�a8�o�X�Kx��C�BHڟjG�)3IBR6�!� �rH:1zv&i��$��-�p4?�: �O1$-,�J5$͝IsC�Na��|&B�h�o�~H�/����ް$	Gpn�ԍ��Q.Y�UNHʇ�Б����Z|��C!7ZB|̅��E:��,>I��Y1�"[�f���|�v�UbK�O{F/���G4���=y6�Z���L�5L�;��|!L��	���6���p�$ A�-����m���6ZN���Й?SGӋ���@Ʋ̣YlவL���O��=G%Ŷ���a|�=����3=aj��f/+��	H� J!ipMȏݹ�0X��p��-�/ �Ғ�����&֣��4:����\�~�X8����A��au���9* ��t�L�H��pd�/�3�u�#�0	�w�p�0qoh�? �qfiu����t�?=�˘Q���$����TX��08s0 @�V�}-���5��\�y?O8��HP}3G¦�wCR
/ ����3a{Ǟpd�/�~f��|dl��a��  �6�::�a���0��M��2d$??���zf� HKg�T��cW1$���A�*$ A�R�KƿV̪P@�b�m�{�ÝC�x *! A�Z�&¥㷅���  Y�z���X�e�H�� �G@��f�N�Ѽp@}l<s_�ϵ��m�pq�$??���v�� ��M���\kk]�� %[��]s�����#��}So���	H���g
}�G 4��㷇{��f�87	j�sf,��|8,5---���;�X�"ttt�>����B�Pz�?�������G����x8u�T333Χ��+�����}���U>�/}����mkrr�ԶN�8N�> k�]�����½0��xo�������\���Gl��Q�Sa��]ᡮ�pn�P��L�b�R�������\�B�`����㿞��G�gΜ	�֪U�B�Sy!����Ǔ�^}���ь!<��cǜ#Fz�=n͚5axx�4Ht1���O����G�	(�F�7s$O�	G����$�����C��dhd�\���q���H~�������K�؉������@sY�`�p��@]�8j�V|���֡C�J3MP1��v?�{d-�{�J��x/������9�h]���xae�ɷ�$��3'��齡Q��������#��;�GP���[�gy�#�#�Q�:��C��͛K?v8���WZ�Ո�E�֭+k�Z��a!���{��	���fÆ3��G:��S	HP#�&��*vb����A�GP�o�^�ĠG���������ʕ+SFO��׮][
��)(Q��^c������u��]z饥��F<�>��'Cx��500u t6`I��yݶm[i�Q��1(�����_*���gqb'3�`�t��Ҩ��i׮]a����'ދb@IsƨܿG�'ƶ�q��^֝y0��- ��	HPk�j]���؋m��R=����c�=V=ei���.�����El�[�n����h�M��_�m�3�tO�A��k��k��=�gFé�` ��`����s�3#7���z��O��NJ�lGNm�_Z�LM"�Lw#����>�`��"�"q�&�jDO���'��|$<( ��$X�X*�Q��+��"�FՈ�k��&�s�=ιY"�l�RZ&��b����.+���"4�8���쮷xO�ꪫJ�Ĭ�J��sa:���	�  �"��M�Γhq�ӎ;J�å"��!����W:X�����Y�X�c����b{�G�'._��(���\\�CR<p6K�����-�`Qf�|u\:r�嗇�(��;w���X�x�R��u�����8�p�}�����@s���{b#�7*Wtq���{���`�XlH@��$X���RoqT?��/e�;3qs},Nc��(�מ����Žq&���Vf�	��x?�gu�Ŋ���f��zVn�J��s�;C$ �"��f7�w.�h)w�,n����ɬC���Z�9Z��hA���+�p������-�{b�^�r����L^/�E$�ZO��H���湜�NM��-�;,�eu�+�� nO���-�eu�0��'O�L���$(��J�H�.G���ˁ�u�˔���'ivv�t��B���T��\�{���w�yg���HP���$��x�^=,���X��!����K#�dg͚5��r�aÆR�0K9����K�Z]�����w�qG��F
��ab<��*ht˷�)k����F�G�;Z�by����JNd����T�\r�%��f���P{��f�'��1~���4����$�R�|��8��r���,b��$�a�鋳v�m�ƅ��7.S�˖T�[�V�^]z4���ƽH�w��������U�����5��͛7�f�iӦ�!�Y��l�l]lc�$V��k׮]��'�Ō3*�&~�1$�>�NI�ӧ�T!�q����\�fg4���C����^���u�hݺu� n?��+-6ˌ���9.��w�������e�  A52^�7�/��h�G��50�_{mmmM93�dqD>�������ח��5�X�<^�ݻw�����&4;	��^���� �f)�P��-!?�����\�+v"�������*�ŽH�V���b8X���ĥv?�p��ť�7n�.ř�Z�$��:N Ūbi/#����C�C��p���-v��/�;~�D;�=F���q8"�ɤ���łͺ���֮]�=��% ./���f�pO�ˏki��
  A#��ׁ��T����3��V�^W�u�b����u[���t8rh_ؿ��p�d�+!������Y�f)�]�x@n<{+�sfX�d{{{g�{b�&���@�HР��b;���m�٠�\�\\6�]=�a��u���������k��cǏ�ݏ>����kĥv����T����X��k����B�]ƶ�eK1��$�9�޾�hnn��1.ጣٓ�����r�XJ_Y����d�ܸ%��w�^;�:~li)<~�<�Vg��n���d��-^�C��C5$ A����7�R���(��PH�21>Vz�N�Ξ��[����?\z?v$<����t�Ng�31$)�P���5\��I���.~l}�����NZ�I<}�T�c4�r$�
��J��J�����b[:�����18� ���xb��EEcŊ��}�#	9��2��0>9y&LL���ށ0�j�t�ˏ�q��X��w���Tfӟ,^�xm̬C�HЀb�3v�*��B\z�o���Y�����o��܋�����7b�Z����u�K�c��}�ޚ<g\Rr���p�r�Ո����������Bggwy�_lS�v2��v1`����W��G��Meϛ�fcZL��3�g����_���=����4�Y��s�7l+��XؿoWj�{̬Cm	HЀ*)�3E##�J˗�3�O����y��i_Q��7]V�����0yfqK�b�>.+y������qv�q�=v.�_�m���h)�w�����P���C�kJ�X d�c���ղpG������"5�8`Ti��x_�m�����ĸ<���f;:���v���5��l�����}���fj<jfjK@�g�*)��EFF6פTs,�}l�`1$�+�j�R\�r����������指��ٳ�,R���Q%�b]�z]i4�Z�]�8v$LN�����tV/,���g�분��8c ��G��*�Q�*޿b�����Ʌ3�ǋm�t�\:j0h���6m�<�]�9<��=��w����b���t�b	H�`��r���Q�M�=Ǧ�~=v�p��s�NAy˨*Gc���ុ��^\�$�]S��NV�ZU���٢5k�C����~�9<|`w^Z[���|�޾�b�~qػ�������q�-.�SѮ��`H�b�,���ᚔ���у���/���f	r[[G�l��a������S'kWZ>�[�O@���+Y�tv�(�Jdc��BaU[��X����p�ݷ�Ç�V������Ė'��r;�q�hժ����q6i���Z��f3IQ|�����;��w��s!Lƽn�Ol�����ޚ��'�K�ⒽZά�`�5���;5�O'�CmH�@���ˮ\74����.-q���уax���^���
SSg���U}��N�Nl9*߫V�+U�J���LiT~`xm͟;��Y/
w����ňsm��*�'�����#�"g������v������Ғ���Z���`����	H�@��r�7�X�.m3����铡���������}�T ��J:�1Ţi�3<g&�k���������{~1$�N�8V���C8{zz�ɓ���D�ʽ'FqƳ��<]I�4��n������<x���/{	G@���+G\c���c����DpǕ7�;n�jUU�:;;���@8v���p3���9<\����8q�Hh��
i��vuյ�w���E��x������r�qi]GGgH[4�?�J�X�.�l�}�z����B�$hq��\�3���'�O�*0�%V��v�ե��Ո#���ř���Kg�ь�~�3'K��!V0�y�M��}s� �j�����^|�*���+�;�ʩb�N# E��\&'O���wW�'
HP=	@\bQnu��f��U��������k6�C��㣇+��8�ˣ;���b�*w_Fwwv�;�?�Z@�b����<���V9��=��Ŏz<����Z�Q����m1����Iu�h��W��3g��c���k��#��'B�$h ����Q�r�U��B��W�\�;ߺ�K]����u��VIi���ʹL�V,�����(��k�=w~�����W�=1�x��~�ejr"���Q]���۾Z|���y��1^�Ç�Y��$h �,%I{��u�Y��G�m)�6_)��έ���؁,��V��Қ�?[11�����0�~kط��s����+V���l
��X�3��5=��a��`��W\_*4Rm��<T@��HPgq�/���+��(�35�o�^U@���-�3g�q]�*�h�����g��q��{�Zjg(��2�/.!��f��Y��M����?V�����U���kh�TG@�:������r��,L:�j$9Tْ�cЉ}�J��ꔏ��,��[�]�����V��N�֕������۳i�e���}U?����@e$����2�t&�i�ڍ�(^K��'��QI�1W����eצW����~(����W\bg�]6*�'֧�f�f���u��]�����HTN@�:�dy]�\UZ�_��x�G\�3�ў�F��T�3ϛ�f)v6�t������5#���Gﯪ"]���f5K˅�u;�mmm�g^9R����$v�=��h&�֬�>r_���,�����]��5���F�vX�zCU{��=1^ӱ�� ��]���G�d`peU�b�����(�p�f�����ʵ�/���3�ynq��b�}F@��HPG�3Ϲ��W��0Κ�ڵ+4�xJ��-�`�JR��0�.������:;���ӧ*���}�� �O@�:�& ����zhi)T�!���T�;���j;�Rz⬧A��^�.<�뾊�.�$�k[�&hV�IWWWUk�u(i[/m�+�1���fH��]\�ઊۗ|z���vV=���رc(��uRm��|S����.�"5��1[@����t�]� ����T�.^[	�' A�Tہ�KϚE[[GU_���.Ͳ��V�5����Q��FK���-aE\Z�^��L�����Tۉ���E����V�,+O[[{��
������j��v�o�A�j�{T�y�*�@��jGKs�&
H-��f�7Z\��|ܼ^���;�3�g6W�F�7l� ��x}�cjj* ' A,f�#�D3H��o�q��.K��Vp�������[L�l�A�xhl������h .N@�:XLg`~~.pqq�Y5��^�jN�j��x編��D�}-�{�v����u���f���NP����ZŶK���T�4��˿��L�}1)$(��u��*}ͺO���FE��Z�y��R�,��<i1�	;흃�	HP:��k�Y:�;�:���jcq?����d-�[�����tb��@�j�ss͵gK�ʆ�f�ăOWXv�:m�' A����y'}���arr24�l,f�O�9��R���ci(\�^d�YN}o��Z�<\����㞘	�# A�t�ӌ��f'�!��N���1�7�?P蘿1���4cg@@�F��f͸������N
������ε㞘�a���ٌ��f���j`:��(H5��fǵ���CƼAe��FK����9�a3;�-��]	2�*;�5i�3vB�⹆�qO��H�1��������fǵ��H�1oP�i�k�Ӷ2�z�Դ(� e��e�rh|~N�F#  uc&h4�l������bdõ��H�1oP�i�k=�m��Ȏk���eK` M�|׆����P	2�*;�54>?�@�� c:�q�I�٣��s�K�<d�Tvfgg�����P	2�*;�4���Zf�=�# A��jd�ٮu\�;��L���T�6tڳ333��� cFK�3ۄa4v�;::隞�Ԇk��YtP	2�*;���߳��>3H�c�(;��<dLg ;͸�D�=gΜ	�ƌe_�q��<dL@�N3vtܳ1��Y3qV�޹lh�P	� vb-�JW��݌�It��1m�LM�v���H�{�O@�:����R699��%v�0SW[��
H��f�|���ӧ���@ =1�6����@���}�%^����@z�Y(��u`�?}��(q\^�D"q����ڊ�F�K@��	HPͺ�+Kͺ�$����@:t4k�5M�K�l���eP�k�i)]�N�
��i3H��n�|�Aɳ)9]�B�Ƨ�H|��6g?[ZZ��0��G@�:�x)����M�O��f:jH�6���Nb@R�.����3U'O��^�R:�@e$�oX�9~�xhf�mŃL[[[��q8p3'N��V�
�^��@�$�oX��.�����@m�=J������P	�$���{e:::�G�-1�Ңm�'��ko������;֮]�#�g��p]����T[�,TN@�:�o\RmY�xV�����ħ/.a\�zu�v�����b@����\.PFK�`�]m5{�,���=�FP9	�ha��Ҷ�ߵG�	q	��T;����t��X����3�x�Z��
���Ύ=* �H��<�ȑ#a۶mf(k f�A�Fl�7n,�P����b�~ӦM����jvv�ԩw ���ٸ���	H�# Au$������&Z�H���ٿ�L��$ -^Hd#�-�[�x�����Xf�xf��-^��[�Zf�qy���l��- -�{"TO@����D'�zF��-���U����Չ��rE���ׯT�=�' A���tb�799i�>|X�Z�C���QZz\�x�����	H� tb�w��A�/ ��Xġ�����H|}�v+ UG�����A����-[BKKK�|1�\���\��[�.P����xO�K��+���T����zr��tO �*���u��W��/n掣�\X�l
H���+�sO�\�Y��E��R�)	C���L�pqqOB,����v_.���+��W�^�v������؁�g�؋T��yU~�|����*�o߾@}�{�b���yp�x���Sh{���ʴ{�n�*�PN���#pa���
XcسgO������x�U]��#h�b�Ӌ���m��L���}������Mc���'^\�F���(l_;��%$h(FL/�Hiubсx �Y��G�)5�ċsO��)l�? ň酙=��Y��3{�x�/���Va�ځ�p~��p��W��H���p922:;;Ou��q�G*�;v�I���*\�n�� 4�X�)�k]�re�	�=Z�Gy$�ܹ3��8�&hL�beܣ900xB�&�yBmF�z����w���H ʣ�>���B>����R�)�����abb"иv��U���xV<`<v �U����+7}�힟
@C���Ĳ�6l���Ƶ�Ԇ ����i˔��ӧO�Χ��F8{VW�C}.�ٕ��vn�����$v��(�WӁ����~�x6R�{��Jm���l�'����f�k�1�B�fW�)x�����q���x��p�WsY�����#�����.�����I�����Ҳ�f/���kQk�ֶ ͮ���޿qe�#�>�% �qP9q�Di)źu�B3�g��������\sMS.����)}�,-��u\~ܬ�������ih)�hv�ϣ��ˮ�����W�����w$�H�/�l➃�z(��x�c�K/�44�8����=t������}�ifhm�=�^���U@���Z�_��R�s�=a���9$./���{K��HW,���m�vEh&��KS�?�����kn
�"��=1~�i�����������k���o����-=�s�d�����v�+�B3�#��.g'�ix��,gΜ	��G��9�񼣴g<�z$x�0�/��?��<gr��3d������,��l��c)�I�PA����e	��^q���޴���G�m�������  ��L�-���	�잱��-?���{�G��'��S��  �ŉB��syF@�ٗ]������������ ��DKO���,K`�;Q���蜥���c���{?����N��Ӗ����l5��9�[^����������?vY �k�u����w�e L省�ys�������>�8���Ua6���<U� X~���	@�x�~����}��/���O~���y/����� ��c����ƕ����k���>�w~���ŗ���������9l�$ �di	��� ��o�/���;�}���'~�=��8�3-=a�e(�� �����ٽ�'^�Ϻd�7������𕷼���w����pN�Vl	}�$ �����0����n�|��������_4 E�yӋ����{�w�S �!V�+��!	��c��K4��������?�O�oe��S���W��������$�9<�bG���� ��}���d~E�f��V8���|�+F�z�<�����;F���~�ů|�����',V���.�����֝y0 @#���@�� ���z�]�}����Hњ�����o|���c��l�t�}K�:��N hT���*@3����~�΍�?�( E�{v�?}�����~���mx�]]׆��������m�N�4���/��/�a�ߜ��+HQ\�����M���O~��������ˮ	F�?>����p�W> �����~���t�?�r�cY�zV��}�7^��/�ƅ>����=I��}o|�O}�ӟ����ze�&��?p�E>������g?��  �`ժU���á��7@�Y;س����?pɺ��.��U����p�S�zݫ��ɛ���O}��x�/��/�����/}) @=uuu�~���M�yW�����W�v���p9��������{��c������������ ����o�N�
��zk �zhkk����FFF4������_��U���$ E�w��/���7_����3����^�����}��}o��fg$��8s����?\~����ʾ��?��]���*�ښ�h�`�����7��|힟|�����;�. �=�yO���?>��� �B�Ї>6n������������y����:^���4 -x����W�t�g��_~�]��-�@��_��iӦ���� �t�W�w�����,^qö�����_޼����<O*)�lo=�?��w��+����_�������Y�&��?���n��;�z�  ����~��~.�����,����_x�^�.��ϗZ@Z�f�{�������^�����oyǟ��;����lG�&�:�ɟ�I���?����, @-�ر#�گ�ZذaC�f���o��;^���\�mͷk����1(���?�X��3_��u����o��޽/Ф���7���E��@���� T���#���o�~��,w[����^��y��(���4^#��������Ͼ��?���GNn�n�����}�=qz�?@��I��>��χO|�a��� ��ӽ�U�
ox����p���K�~�yWl��?z���~�%k����e��l�p���س?���{�ȕ߼o���xx����}d�}�����̽��//=n����O~2�u�] �epp0���Pi����,'�-����e��j���o�l�7]���Y�=���n����#�k�o'OO��������m����gf������Vh��{{�7�o}x�?}[x����{��/�η����G+A@X�fd�O�����������=B|��G�G��@>��k/�L���t�m������=+����!����D|h*��+�����a�޽�|������{�7�����/��?۶e�]HU�$hv�֭{0>^�������n���{�}?��7����{��db~~���{�ߡ�����~M.FK�c����'/ 5" k``����79������b@
�d�Ν_okkUe	;r�'�) Ԋ�  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��     @B@  HH   		   !   $$  ���  ��   аr!� �	H���r���$ZZZ� @�$Xb�i64�|K�t  Ȑ�KL�%7�Dk��x  Ȑ�KLK>�4����[�HS��.W�y�[Z�'�:	��B�p"4������(�����|�y���|��A�z�`�ii�5M@���?@��Ғ����$Z��eB$Xb�e�Phmok� E�|���[�Z
���$��[� uАz� E�|n<����|.4M@jk� АV��M���t};��
�S�I��h{4 �������ά���R4�����%/�k�=H���� u�pV�}��%�4���G_o�-��A�2# g��&@��-�S�}�7X"���6 ����2<������	����i���"�a�2!3�P�o^��R�z���D��-	��\.7���W�~WW�]R�ӵ�;C�����mX���@f$Xb
�֓Y�f1�����-��myw�n���3�y�|���e���*~�,�~�|>����p�g-;�l	H�Ĵ�2H---��ƕ;��TKK>��'�\�^9�W��G+���*�l����f����lB}�=ڶy�Ȕ�KLGG{��`��R}��#+�hp�����3H�Balff�/����f/�l�?f������ǲ~͖��L^g������dO@�%������_�cEWj����u�%���j�!����������^��ڞ��hd��G{{:�XVV��F֯�ޱ"��hkݽmˈ�5P,1�B��ʕ�_=|�ȋ�z����T�����믾����D�!lܸ�3Y���識NG�×n_�����ٹbw�������x�\>Z�:R�+.���C}H�]~��?�* �٣|
{����uWm�ҵ�e��u�ioo?899�:�׊�ή������;���%�,K;v\����vǇ�x�����z���Sˎ�~$X�6n\�?��=:z��t_)z��j��CC}u�[ߐ���J1���暝�������kuv�CR�@6mX���b ,[�\��O������OlI�ur�|��L�%Bgg��f;��$X�n���_����.�N_�oi��mb�տw��u�hX۷o�����?;yUZ�;�ݽ�!m۶��c��5�,k1�_w�����[�"����Hu������믺��f;��$X���o}����On�������w�ށ�=_�?|z�e���U��4�x�K_�����p����ʚ?>�V���Li˦����ǦM�����k��T`�QgwzG�C�	H��m߾�Ǐ�]u�}�����Rh�kk�|��}dۖu���ZȼD9Չ�_��������/���׬dW��=0�&�,�3�_��[;������k�z�cǯ޿��+k���m���c�����vn}M>��@�	H���põo-
�w�}�;j�|�|m_�[���U���}뺷�X��``�Y�r�旽�/������$���КTK$Z�Ǯ�b��{�w�����K^�����>��C�~�����𚐖���ζ-#�
@��`���+�����з���ߟ����9b ��
�ݽ����]3��7�[�8\����������n��ѣǞ]��C|)x���7s�(]�c�O����4��D�9Ϲ��]]]���w,f4�{�k����b��j��7�V�G@�eb۶-�q�����~���{���TJe^T�LL�-�wm�WYQ,�ύ����C�j��ӅB���������+^���)��7�y�=�>y�ԥ�~m,��;:��ϧ��F�oY��u#�)�v.@�UW���m�6��;��}?���T�������r�Z�/Z�f�^�m������H�����~��o��cϞ}?r���8zt�Ƹqynn����{���ݹk���_޺u�ikk=^��Γ�&�95>q����+���6�����+9�ϟ������;��=�uw��3��mٲ��q���5{����Ç�<wtt�3g�_�R(�jmm-�::�Zi�E�GV���-#�Y|�� O�ٹb�s�{���x�u�Xl�������w���Ǐ��ɟWhm+�����о�3�r�T�>}�]�pɶ����<46	��8��~~1��.�i#>\��@��q��ٷ��/<��௜���Q�׏K�FFV��MV������ Q(�X�.>�����N��݇~����?���ǳ�6�k_��hx 57�v���q���g�?p�9��ə��>_�%wjh��kW}|�p��PC1���������G���c�?q��y����o�Z5��c�mk+��! ������z�o�����zzb��c'^Z�x���Ԫ�ٕ��ӫ�����խ�±��¡���Cm��#���C+��w'�ׯHY��ٸ~���czfv�ر�����b��tpj2�zzU����b[mo�_l��mg����~ɲOX��M2_�lq    IEND�B`�PK
     @^�[�z��gW  gW  /   images/c64d4bdb-8b24-4d1f-9af2-aab9cfab9f47.png�PNG

   IHDR   d     �� 	   gAMA  ���a   	pHYs  �  ��+  W	IDATx��}�]E�������M��B�� ��P�_A�O�C��ϊ,XPAz	B��Ki���M6������;���;sgnye����?/�޽sϜ9gN�937
Ny�}�^?�ٕ��#���tú4�Nel� �"�_�@	�B��)�D��*�ף`�w�X%B��e7�;�f�lH�{xa�b��Ϛ�O���N�m����ԊZv���t�JC�P~��� ��}��}5eUlO�e���Q��!4b�����So�31K�x]�}�	�@�o������i ������%������#-#$��nozuݑa[�P9��)���xh�脃*�[������
���sl�O��Қ�5nPN(j�xs�@��!�S�3�+�	�L��VW�,��ms:Jh�b[4֓zhsπ�𓺣���M�TSeY����28o+���v�[�L�7�QXVdp(��G���W#6�-g`��ȁI�_D@q�ߥl�0d�O�9o��(��(,{́�rO���16��+F>F"b�S/��,�z����N�3 (s^0�����4�L<`�iٳIv9��(^�P��msB�㬋���jNlHg2u�8��ax�Z��cgl�ߞG�.B\a�������I�2yK1$� �` Bʹ&����o����3r�ʓ��3B- j;��\�r�}HkGo�ա�T�Q�:��� �y��ŋx�J/�<(Jqa 툝��b���	���T:Q"L����1�.?��&��&�R�ȇ�c�|�5Fr�9�v�ԣ��T�*\��� �2��] =�^|L�=�c���%jV������qK�@7i��R�;�XR*(UF΋((d��;��V�޶ѐ�d����TS8Ø:�j�(:�K<tU�@P�ǰ�Q�i�3�B5��p��6�̓�i�Ȗ�T�́Č���xTR!��8n���eEYH�d#q�GD'��"q�0��؃��� *�� 2�x7Fw�W�m^����x�Z�Tc���{E��r�Q��.���Q���5HB~�wбj��b���i�ބ����$K'|���y���Q�Z�}���o ��xE]��ђj����#�@0�pJrb�ttk�i߂3��	����'��? �jm��'Am��r\iU3a��GAD���i!����U ��#u4g���tY��������cV���8Qˬ@�1��l]TI��.28�Z�n�6��sN+z�OE�G�G#�c�D�|�[֏w}zss4�3?8��P9ԇ��zAԔ���y��:��w��2�|^��$tR��Y��X�՝]Y$���o��@'T�@���4�)��RU�'*DD��mF�Ċu���k/,-�~����5���/�o�o��P*}J�k�d���X�5%@kKM�蝓٦���X�3�d�j�v�wG����\p/�}2��*�C�Æ3��l��(zSi�N�K��nj���t�w�a*�*�_W�pG) 	]�s��3���!�H&5u�"j�f!�	G]��d8�'8�Փ8ٮ�C�O�_L챯C��D�����Ġ��{��g��iA���u(<�)�9v�b�H�>T?�p�i��uꏻ�C����۞HS�R>�:[��r�g1��f�E
��A���^�8u��RUJ��z�����&~������Caޗ������@�h8���W��ď�#G�7R� ��)Q�RL��B�a*��ĞF�8�:W�z���9�8y����x�ħƔP��ax%�q���QS����y�.�����PL�S4��	{�%��D�kӵ�$l��� �.��C�B���-C�p=�m��$����4{}���J_7�q�i��'���2��cT#�r;������ QJ0��jD�R�bX]y�UX°�Q�6��3dG7D��y@\]��̬�Kc!v���I����/���,�f���ZH7T��O#�>���Ⱥ�`�2!�0&TCj&�3R|=��J:.�b0B�9<��S�$�|��4gN���1�r_H���h�l��NȄ��̐���$3άDH����'6�B���� �Ż �`�(�gQR"��A���M:��%����Y��tY�A��8Y��(��T���Q6K1W�B�AMͩ�6��
�;��y�z����=,����w�H�K`}*��:ԩC<�>����D
�F�~ee���ߑS�Py(f�����j�H5l���(/J��U��Z��)@I�Cr� �M~h�ʔ0צ�8�c���`H�7~�}z�Y�'�wPzp2=Zw�Ki��H�SZ��b�����~�,�g/�,	e��:љ�ҙ���4���IX��y�Mw�ޑ5%Va u���[h?����(�!��⹮��ğ[�h]��zטpR-��QDu�h�ruZ�F�pIYXK������\E�-PBF���mg�ϧ]�a�f��*B��z� ��4� �U�b�9���:�UI�vq�R��8M�F��9$�W���(5!�<E2���?<���1���\7R���bz�ސ�f֗:�"�HH(���&]�G����,2�@�	�:C�W�E�J�IZ��P���n��,�2����BW�A �,j��Y�
l[�c;����RG��`�n���*�H��/n9p�`z�h
���]=jK)�����`�P����qR��@���k���a0^�("KP�Z:��,R1�ZR�����&�ܦ��
�y���;��H�%q �`��0%3?����e9 ��vG
M ���Ԣҭ�U��Q�ː4�}02=*W����%;�)GT{��~��hP��g�lW0�Y���x\E��=���ns\fP���e ��3�f�\��CT���bxnԬ��:��4�%Y�w%b!�3D�mz�bN^�3���wט8��I�|b���J�����^���5�9�IoI{�����3\�fe�1���^�����R��6��Ut��X:4UlX�@-GI��{Q�J���{]�C�5�編DՆ��af�E܇��=Rg�N#%�N\#��j>H(�l� E��R�� e��z���D7�����8׎ȶ����$?,o�V��!h�"��g��Pn
_GR�a�yH�؅/��ψ-�����nAU1��p'�'�$8験un9��*�
=$W(]QQ������r��1�����!2�ҝ �L)*�ү;�����BZe�����a��PH2�@�S�IB./˯�&X�rG%��1<#�G�Ԅ����SL]�hPٲ`$�c�IG%9*G����DY Zw�Cט����$��&51q�q�c��Ɍ�!"�=@�v���l��iN��}z�!5� MM���;{!����,��Xi8��ֆ��
��/	�um �G�7]8��=�2�*y(9S�tc,��v�T��T��PSɹ|	Wz�J��qbu@t����ͪ��dt� ؚN�!|�,��:c�0zj��z&��E���D8LUO�!B\�ыn~��P�df	U㜻��?��s�cW���ވj�����^j��r�j4dc�T��}����'F�3$4�I44zh��l���A��Lf;#�c�峆TI��C=�,C�j	������15���?yO�PzZ��`QoC�M}_x	�E �6�m�̴���C�E���S�Y̔�ua)�;���[����wH'
�h�`����Ǵ���}����#��WI�uB&��v�`��	ً+�Y�gZZ7^/�P`Ɯ�{�P5�vr��"7��1ڂ���S�UV�%(�;���0X��~>Fz�g}����y��{3�.��-P)�![w�����t��y�&/_�O��>�VB}�V�T��"�I�ȯ8P�c ��\8������xoNN&J�DG�W���Э�1r�C3�#�!wt�Z�IsT��tz��B9h����Q,���MI�7_W��#�){�T_.ŀ3��䬲ǽq[т+�<��� 869%�^����	�������+�mk�2z�zTH\;��L�
h�iį�M� �1@���J��|�u��f���f���C����.�{|g�g�u�#��TwQ5ۙ^���8/ħ�ȁ#;&b,���ԉ�S�	�p��[�դWO�,p��c��i08��_�� ����a�����!:��"�l�ͱ4UY?�^�O�����2c+sa#�O��q�/	�V��SnH�@.q��&'b�d�,S^dT7@r�]���*���m�'N,f�P���Q��t�8�>��[�]WS�s��ޠ>E�?��]��p�͉�_ғR��z���ђ��ۑ�C��Q���4�.8*"(!����ǀM�;�m>u+��:���@y�u���Rm����^��iOڴ�.���T�����
���������8Z^�7���Ц�f?<�+>P�u�	�S�ܰC�a�G1:b,���ŗ��|h�05�z�����Ĕ�ȹ9q�!���3��Y��mߐ=�����3�Yff8�)u�f�4#C��:���m��Ld�	
����Z_�io�\�x��6��#��*fP)f��5���$�	���Ҭ�K���?�.�m��ϸ����3��u��1<�:��A�uek����(�T�� 5�0V�K��t�P�8�&�F+w�JBP)��hL2�d�U�Ĩ��>�m��J?3��1�9�	��8�Cģ[tz9�l��빹ϩ���mh�ȑ*��S�K�i�(.I�FH9�d�X���/�Z4JL�L�=x��8
:���f��"������_��qЅ7��Ҩ%֭�,WUJ��%�C	2W8'�b�?��d�K��r�o���3�[µZz�*��:�R��kg�c4�:�
�M���'��}�Z{ ���Z��9s~e��;VD� T qz/Jf����ޜm��|	wJ-d+x���h=��_dm�X��j�g�ɪ�!5k��m���%�]����lf%nR����܊F�ޓ`��	���ї���d1�YP�FɈ�����a"6��5G,��R��I�q'<�� ��!<�8�yuL�w�9�va�}t. ��KD���C�|������<=���!��T�g��3UGt\Nz7��	8+z�'9H��;.� 25/H8��S5�Yg��w��܀*Uy��/���2������%����1��5��е�Amo����5�?k���䩯C�=7��P�S-i�a��\�+\g�(wX�c�d�ޕW'x�e\�`Ɏ�%8������	U?s�S������;>�\',���2H#�qTbг�o��'ڿ�pC���� ^�g�^�G��{������8�vX�󨳐����Z0K�H:�r��2�&;4^ӑD;��6�P�x��J2r�A[к�YuQ����<6M��s	7��P�H����h����O/Rƨ���z�0�D���N��+t�uY�k&]�K�-���%{���\���F���+�D2j�z���i��Q�a:�Y�K�����ȫ5��Rz�%\=K=��ۚ���JW�B� ��W�����ǝx{�6G��e��b�O�S$��Z��㴱\��U�)�(~����qe��(��!rE�X�S.����Ϗ;�����&uc�Gtfx��t.�A g�S�6����bܧ�_���B�iY��<�G//^z�Ѝ1�)&CX㙆J�cxr�)lgā;xt��S6�G�}#�]�&�n+ �80���;H@�ܡ@�nfr���'^���:X�#�����R�5���y�Q��p�-ξ���~a���e�FR�t��zB�=����;ax�ƹ�:L]�ʻ�]�tn
�G�=�:p,��K���N�z�I�j�I?"�jٹU�������E�/Y����1�� ��`�YS��:·�!qfʒ�[bnJ�xi�q���#�m��_6$��ڋW��ݥ�R��L�݇�5+�5lk���>�=���Y�	R#��j�8
��>̭TBJ���}��\&����7�\��l�Q%0$K
Yn@<-��:#�8Y7x^r�,�O]�� �f��}��� mEM����6I���|���*h*��S��+���ޠ��������,J
�6t1����T>@��ԙAi�`��ם�w�ڵ��)�!���)@Nj�G�|j�a��0 ,G(�!�j� ד�OI`��$8p��FO?z�z��6P#ܘb����zq�ޕ:��qZ
���Rr�,�]��iV����8&�!�rP��2�1��Y,ED<��/�2P5A��`D�pe]����rOr�axǢ<�U�"T9����{�_B&]-�mj�����:PuwD[{ܥN[$G����8�>(8-< �0�Ġ8Ne�ӝ]�r@�I� �������"Z�����	D6�:S�Đ� `����vP�j�{+�=�qG�߭�U[�/L#&s�� ���֖�:gZHw�--#�4����p���f�h���{��Gf��k1�
yM��*!g.�!�I�*;���:r�)"�"p�[�����F�t�"U~�g�Pk����׽+����h��)Y"u����Q���T�f�S+��|i��g��+}�~'R�K���z�6!���g��~��xZ��?ǻ I��M�W��*��l0u=%��I���9*�^���?v�b���IASGGD]a)��_rr)K�/F��4�D�O�"D����k���w�H��$4Ofh!Xh�mCԈ��mӀ(	����׶�uT^�y� �%h� @K�!�p�"q��D��d�X$��C��������W�u6	�p!�Y�1;��Zp�R`U-��:�9\z0'�`�����%���7��G� �Hh�/��nՈ��S)&RU��d����Ï��/q2$ݩd��U�"�C��w�I~�XH_
&����_���hC̭\��pHq�)7�Q�P��b�0{�����{���>T^����1� S.)밥���x�(_.)�)z����xD��Kz��#�;�DY��,&.�eE@+���ZE����x��?�ƣ@���0������"�;寂�Ǉ�
���p�Kn�63̵Gd29\��5�J��7�@�x~h$>jM��d�57F@�J����G^�^6hmqAv�������례�W�GD�F�g|�ы�1p�j׈�r��Ԅ�G	L%���8�'�qɆf�=���l��Ug�<�!B����0�!@ia��/sq�$����u
 i<�\�W�$��'O�r5���U?`	����Z�T��AT� ���=�R�o��u�d+��!y����͔�地 7)ۨ
���{,p��3n��
��*j��Ou��R,����e�u!/+�;�}*��w�7�R5r�N(lV�F�º�� �(�H�j�ٖd����A\�����Fi��@��$$*޷0xڑ���Q���0Dl9�+!��DP�vb�LiDw�/_6�K
��s���\;���, �`%��}p���A�W���L4|D5����pb#}+�������R��B���u"~��E[]	�-� i1� �
�u��;�겠��H\&S%��! �)�k��s���e@��� �KK���Ii�>�F|�Kԉ�A�η3����qSI�R'8���3��ܓi>9L�{B��e����o[4���掐��\~��I�`3"�o�Q#aw�k��&5��vE����x`H�!��#<Z��l�g��i�V:)��`�#;��$���YSO֋����e&V�D��q3tR�����LLF���G=9%�$����KX9���?�~��*="߃�LY�} ����oz��Z�"�Hh����1���Yµy���v�,6f;��lU�,qHq���i�,�w?$�{ي�*!����;�������^Td�/=R�p�ԏ�3�}A��nU?L;႕]s$��5�?]����1���V�Ԗ3�%�yE���7�]S�kb{��8c��<�^�d�͗���6I�o������w�~�n6�y}nl�cjPdW��(��tm�>����q�����L����n�!aOgۦ\��/��wwII�Iz��	��y�����Ѩً2��������ͅ�0����F}��f��	��_�kR˱2�HK6H���V����W8�c����O�5bJ��|����x��3߿�a�@�q%P�9��z����f;�V�$�!:�>����s*@�9�eL�������Eޢ�@&�@���譹�A��:Ï�0a7��g�(O��1��m�3�l�y��v��V:�)���n�M.q���!�(����K&K��pt$Z^�O��P��b������&�b(�"Ψ��t�#���5���3-�)U��T����}z����9k��!p�!qM=3�Q��|=�A#����B�AgC�0 �����!�?���@6R5F�'[�p�nS�^6�n 5�+��52���ZxQ�y<@�%�����0����Ŋ���{�Խ.4�ĩuM�Q0$=N��p+�v븖+�b\����a��`:�ի*����5�A#\]&�5^�2ugӇ8U�T�t��U��� ���E�h[��|�eU�+	�j�xU�N������qL�ɰ��Z�$��0䃎e���pB�C4#K��H�4���z�~�^�t�a�9 (&:(wLy{�������$���(��fi6�r-7�8��;�����W�捣�$5xu��IY�CxE�`R�!�����f�s������Î��@�&��i�hw3�<C;��&�}�Ho�f'g�Q��ڗGO.�_�B�0$�k�%St5��Y���!���4/�qU2��O��Èh��)��+�ɐ�!����T��aF��:�?{�Od��2cK�5��7�@��TV�nk � 5#�U�-����T��(�R�ة��ф��C����km�� �NGg�����|+� *��g��N�i'�#D2�Q�T�Gځ#aR9�2o��;����%��4,�-�2��.��m��p"���h\����s!Fz�T͈x��L��㪵� 7U(�[����]1��3;����[㘾������M)����wh����i6r"�Y_��.�7ӹ�@�k9F�;� G���Җ9O$&`M�lC��PO�Ӥ�xy��)	P��@4"��k�rDr��c���oY�l���~q�Y�.���b��H�7R�p��$8�#��Y���D��]&����rZY�����5��	I(���Jd ���!��T+�@�{�2x���GV$�э)�Tn��8��fOVtF~>Vx).�f3�TWl�	�S��ߗwF��?��ӟ%����)�p�GN�/�n1�o�d��B� ��z �=��A"�j���uj��j8�2�� }g��~ֳ(gH4Na�������f�D'��H$�1fX��� ?�3���b���)^i�B���!��N�A��u�bx�K�q~���&�`FM����;��k����1>Xť6L'	w��/�T�	�GSi�+�����͌�k[�/	�n*iR\lHI�ʲ�S^�4��l-�*FNF����$e�e��r���f�%vQv��ng� ����� %���aCz�!����`�@l;M,��!�&�Q�S���8,wC�x�O$�w;�L�l ���H"yf$�Y�9����f��I�{R,�]I���،78k�(��2AH�4�~��HU�óϾ�]'�hvM=�Pf��su%p�QMPٵRld#�mV�4�Y�`ٶn�G�b��ZIUk���/UZ��-6w��9�� AY�����o���=�9zv#��쁁DR؈(1*+���.9��Z�?������vo\u)|�̣���v�K�c��de���J����&�=�����Nţ��������_�Ę6EA��,_<uo�[��D8V�L��=|20�~��
�v6� �\w�p��:X�g<m�p�	3��#��ky:���r39W)�!���'8:�z}� �:�f���à-�?���B��PU�o\|�[	]��>�a�"&_8�`h����k�x,
��y�\z87o<�d�'��L�-����P��{,�:��Le���S�S���]m��8C��G�h�/_p|����@�Z�fH�Y�#����L��d&�"�du/;q6<��vu��w6�ئZH���!��>v�lX��<���g��9c~�@�	���=b2����^��1��`dn]E1����E9�����>��9��*y3�<�q���,Ă��:t����k�CL$�E��'0�KU���GϝXS�z[���Ɉ[uY�y�$^7��5jY�#��F� ���S�`b]�����B�����ےC(�a�gq���m���1!^.�E1�gLs�w�@&(�-f�����bx8 &ԖBcU)���
�p� �q skY��=	�#J�<��6s���ϼ�T�H�*BCϐy�x��*��r;an �Ʀ^N°��cPH�Ie�Ӊ�A>S����8����XC|D،��g��t"�H@9gv�{b��z���f̜�W�P�kڌ�PS[�񌌐��%��J/jgנ3jD�f͙+�]�t���9�������<pNgp(�<���423s���&s}���b�F�hkg?w����m@��ю8L�6Z��a�����H���&s"��0�H��E'Bj|fí���tvBEe%�?AI����.�u��J���xau|��Y"��!9c����� T�Բ��X�V����ol����h�_\�
�L�����&O�
�uu�����P^Q!$�٭��;`Ӯ^q�����͌Y-�(S*�ޯ���N� �2���;ab�MK8�(���٢��`W5��-��-{`,s�~,c¸	��epC�6���*���oɛ!1F�7�/�g6��.<ݧ�����w?Hl$�=K�����@/��c#�׷��7���U�Q���+*���JpsqN�ϾǙ��"M{���[����	(a͞[|�H����W7�A�����K���Z��	I�3~gc������읇�%�X��<�.T��ู�x���-���q�S��K���C<������p˽o·/;���b"Ϙ�`��t82U�m������ʪ�y��Z�7q���h)�H|�yג��tMkvx���d��I�����8~��A������A�!}�CDG�W����T8��I��F$�)ؼ��}<�n3�_��	���-�p���e���n5z>د�����	w����ܞӿGb����ކ��	k�����M���5�6XrE�b����O��U�:��Eӹ$����j��O���e�'R����3�(p����7�*I����vؙ`�Ryy��d
��>�.����1���d:�k`�aq.�`�<Ĥ���7�������j�?�����>.��$k`����D	m�.���7���&9����˲�I6�u8q"�zs�;���Vy%� �� ��;���u�9טZ b����;�{V�Ћ�ָ� cֵv��{�� ��gQ+WA�#��*��*�Qyv0�n��}aA3\�%EPT�|��'����L	##$�c�\��tH��O��%q�WK,�f$),��Z[P߻���'�ep4x"��j�	Q����"��߿��Y����+��=�!���a��W��/(�$�07��R{5�,l���A\R-)��-��$k+�ڌ�������k�;�{��%�YJ8CG{�N��C�ioeg�a_��&a��N�NLK���@�>@
-�^oX]�@��������j��a3JYI<VQ�/��E1w�Q�D�u���?�Qfk/�i���22��ݟ�;be�_NLGb:���2�o�����}��b+��Uz+�3	���+<�J�!)��|��!��h!��e��u�N��I���8�j~+���WF�i���|�a�|��)0sz���5�%P�B"����ؼs�k������DTT=�ۼ��K#��=��a��7'W���p�/�s�jj� {��i>�z��I�������'ô�Y�C��������Wê�mjy$N)��)��M����WA �i�? dP,���2؞�`<��W�SB�;�(�0t�3�s:
�=`���}g'���[;��;�������G��X�'��������?_~~����|�N(���#��e�qӯ���Yc+��d�3R���m��էM��:j��N�V�`R1��
��ѓ��c��k��|y-<���b�j�Jڐ�i4PR`���28j�D��p�3�����͙�c�I0�AiA*�j\0�
n>k��)�c��7X��XF���2Ȉu�!S�Ϟ�+��_>�����a����@| ��������~x�5���k`����I�%L��|ɱ��I�'�lk���#YP�S�	����8���9��!����N���6Íw<ooh���gRQ��B]�&�,��X|�"��X�u7\������ރ�t8��I��-��e��X�m��3%���F���Af��p�����5��>���姡op�3BL󴇒PVR
c�U�sF���@{�����P��$�#�C������9��f��{��a8���ֶ�3���3$�;�U��]�g$�|дF�5SSH�?<��x�����(�	�=.9�d8a�<hWe̘�ܰ��!�غ�{W���6���C��}/������Y��Λ΅n�;_2��diLYZ�r�ײ{�&ǩ��HE���N��w�R�Z��S�0`$�0�=\7��u���x�����<��DB#?ul5|�����.�b�j}U)�,�3�{W�y�-�郯��V�dN[� \�?��'�}9���ˎ�;�"�#G��m۶��w�T�Pl����tڜ�\ƟS�a$�^zYH��.8
��;��|���#�����#g�/�?������b��ŋ��S�ڟ<�Y��҆L���0	|�[�§�9�������;��B�3����b<�s`ڴi��3��5�\w�u���[��������b����.b{�_��ޏ�<[��9pח���?|�xx����u/�������[��'���?� ��w������r�E�]}�@#��dΜ9���k׮����y��a>�a���T�D��N:���rx��U�8����-����b��{f���Ͽr��#U�3��?����6��+�$%�~����76@7��1��?�<<��000��黌�����/C�r��H��B�*J�xІ�T_8z��(����X��Id8�9_�d��p�cʆ�N���ULJ��O8 �_�� �H\dps&"�"%�����n���Z.���o��Ȃ�
��iF8�V/����������f�N\��@��H���� �Z���s�#�+����3�fk�+K�ҵU��e9�JAO�w�y�L&����x�p�i����ޫp�CGņVЍ=z^�����ж���=�4�ߏ�vȈ���w�)��LJ�!�yw�.�u�^ܜ�1�
�%n�L\��#����^��z+�����ŋ��/�!#lBpd-�>�e�v5!��:`�&=ca4��̀��m)7�<ǘ��e[9Cp2r�JT[������^�ux��`���ӓ���s{ӥ��Ų��S������#>U.�9��
�logn�ȌD�ˌq��;�O��"�r����7�̥��C��c��C=���y��$#gC�ؐ���Y����(T���U�{�/�NW�UЋ_W��H�lm�1եMͣ�]Ĝ��N9>���a���M�R��.��B����7�|Ӹ�N��Yt`S|:���*(hTQE��= (/�ѢX�8�g !������{L0��	Kd�g��駟�;���~hhh�;v���9��%���3$?U��r�ݽ1T^���G/�����+v���6v�[�
�/Qgz�DD`�N��I�ܹ��2s�H��|ҙ���x��*����z�9���x0Į�	��"�\2L�(z���=}0���"q�Kw�;н=��Ep�M�C2�.P��|+��n�FN��Hb�.c�����a�!3� ��U�r_7�oom�7�^K����g��o�h��[�v1Wwޤ1�Č��k�8#�qc�J�W[vu�\[�H��}wO�)=��ϕ���ĉa(���{II��^V���8��^�������5U�bs��i'�D1�,-�p�YG���7��O��
��@��mJ��N:x
2m,ܳd�@���r��q�#�����V���+t>z{,�UE,��ެ�Sg?#�s3������2'�0F���gBê���4<�b'l��A��'͐O�����>���t��W?̓
���g�wp(t�;��{�|�u�M<�XR��IΣ���k�8F����Jn�Pˣ�ǵ{�?pV�����-n�����8u���`"v����΂��Y���?��}�m���h,l��~:ڠ���g,Z�ՂO����w�W��O|�
���si
�)0J�%Z��8��� J���N�y�-����l=��v�㯭W�y�pX0����I�ֶ�a�%�����	+�]ϷeؕBf�7��ɩ�'�cJ�Yg�/��i���0y(��4��ކJ{Hd�������Ȍ�5�c���?� ������3����_����A��C�w��nxf�&>㊳�o�o�Af���?���ƕ'�H�o���S4�O�_q�|~�"�q)) �^�bq�䇟:�E��A>Gסz;��i|���4г'���L2n��3�+`�;���T@u-��� �In<�0	��	3v���;_��g�gj����1��+��9.��}!k�/�"C���A������J�̟�郯���{[���%���M�X0(���yp��	������Z5��oA��ҼV��Θ Ε�������l�N�]�.��5����۟ZG�~�G�h�� 3f���c8e�|4� 45�| �l�Kw��2�c�G�Qp����?�(\y�A�{�ʼ{�Pu��������W.=�����B��A��S?�{t�5�[�����c�lH�mz�_��8�B+3����7a�'����^�G}hi�8ΐ�����g.E��æs����Y���*4� s������r�e��g��#���xܜ����#�q���c̢�������^���
��x <�|�i�;\���C#�i<_����XH�N[W?|���ߞ[�U�<X��7�*�ЕL5����?	��=|7��'b%�nT�Q�$,JJ���'�<��~mjn��L���p���H�4u* �>�g5�_6	�{e|���p	���JeȂ�Z���1�y���> ?��i����Vn�#��#��??���n8�H���3�<XPAt�����1@C-W!�V���5̃C	��oC��MrИ���чυs�X��VpL9��	⸜�1��ڸ���-�z���u�������S���V��&A��w᣽�z8~u-����\������#o�xW��r�p�?�����T������?~�4�����3�n���\j�;D⿹���-,���.�d�h7Е��kO�׾����n�ߐk�@�'�J��#���\w�xf��}&�����.C�|�1�>V6�c�]0c��1c�PC�H�^��UL|�+��f��8 �}w+���)
����鳷?	,���|�b��WO��*����7��pT���:,�9.	�щ�A,>��+O�˸X������G�`�ax̠�l�25ť���Sn��{�El}�L���;]��F�(�b�f{�0��$� ?3��j�8�Ө����6h�	ظ���ֆ�r�����!��`T'W3	������ן�p>�$��}/ö]3ʒ9�8a+2\6k<��U'�Y,��~�����G�����pf��i�?��=aJ��^����mO��3��|��y�]4���8�(��;j����f��NAF�l����6W�DFՃyT5�yA��}�~��2�P�y��%O��� ��b<;��c$��=}��_?23F�ja���!�GaR]i�sYe�S��i�#��Y�8_$?�Hh��?��K�~Go��1s���/�v�y�q-�6��i�34�8r���p��SY�!��c�h�Л�ܺg�6CgFPA�q:$��<g�[�3���;s&���a��2p._�?�24ď�b��K�9P��w�D{{}+Op�h���p���9~��JB����#f=c�ӟxc��y}m���b��c	I���$ �;�j�2��#�n�F��^�Wð
��h���vR3OG��($�&��a��XgL��s�v��
����$�=0q�L%�2�����Vm��������Df@^��$�=�{`ٲ��K ��w/���S�d���?�
�i�s�V�[`[�&�nno���h�1��1乪9�Κ9���ٛ(8��1:�m�-9<��ID	�K�����E\�@q��?
�]w੬o��"�p�}y7?�b�]r���1E�����cf�W�솿VN����f�.c��񅹾8��o�%pWI7\���Nf�m~���u�8�*h[��ЕM33��4�xǷK��d�T�PYDp�9O�_q<������R���|^x�شi�����A#�����������W��x�-��5.��
3���KK������a�6f��(�7���A���	PWU����<���O���ȫkv�`2%f)�nN8h2��v>���b���tx���������3h�p�r,`���<��z�Ez�	&�W\'�x"L�<V�0c���Ʉ�-o`����ן{$|墣���>�p<��,��Y0c��B���%#�aȌ�[�����4�g��'�/��
lo�a�����SYƧ/p�sc�-<������O�_�Q@��_�~�ό�=l4���1��*���E<�gޣ#�{q����H��Dċ�}����n�	֯_�,>���N'Ŏ/��8�e��r>r�^�."ܹs)4�Y��0�ٔ�21="���G�:1oifnM<[1	�n8�$m�çO�Nf���G ΢ګN=~���|Sή�~���g��&���~60�o��)�Ӆ�q�Zl8�}f\yޱp��g�̽��{^��|�;a+�"�)��l�28���yN/2ӂ��s{�'=Ġ ��w�񙳙�~��©N�[:�ùm��BC���r�
�"1�]��Q��p8��|6�?��)p��Yp�'~��D��-�7·�H���?�gc��`!�5&H��gY'�W�{��y ��'hO
:N�c�q��;V��~Ĭ{��G���wЉ�
sp0An�ܹ<���+��.�c�=Z�7$�G�˳+x�p����R��#o�E�Gâ�p~�F8����D��d,[�c��q�ϒ	�����r���a��1p���͉�0;���%/-���~9�|�H��o�V�C�$8���ˏ�S�xh �w���?5���2o����z�qN�[%p
���t���7n���:
�8����uk���:Uǝ�'�y^?�?��ͅ���<�.��i%�mP:$�dE-��V��:7���~�|j3;Nc��O�.-;� �t+lٱ��������x�n��o)�2���n��~� N��/+/asm	��h��T�/���(�a�@�(���7o��������� �y���=�0|��ϼ�	�����������q������-мi+�	(//��s�Ñ�&��3��<+�C�t<*s�cnb0TY>{;
���_�|2s<��TY ��������)}�ʀk��S#�>�uGm�8m��~�dx��|���a�t�Í��쳭c �����z*߰s�Yg�u�]/�����+�>���@.��򜰬V/��v˟��폼�37�.;� �<����������m���^�7�5�5��U���B^\��~���T�&����<��ƂV�F ?��G���s<������w�Y�]����Y���!S�a��o>{\p��ݓ�|��w�|�"8�ƻ�?`kɒ%����ok����=Ӈ������/�)w梜�����xq܏kLG㔆�A^�.H��<�;Q� ZQ���ֺ��5����(|����!���L���ޜ�����pv��pB�����KG82�G#^��E�z�APLY*ƺ��;�k���(���p��O<Ⴡy�r�"��U8k��`��Alk�0UC!������ـ��^�x́�0�
������T8t���;{���:?o�X����8ۋS�,]��;��f�97�*U�G΀�Y|q��s�1?-He�Ӏ�{I������!XZ[[yL�-����H7��w�Z�Xk�8o��7p�$l�K����͝|=���J��M���.�vw ��ŀ��F��i=O������-�Q���\����sS�����wx ��ˎ�0�c�"��I0����u�0{�Xx�l�c}
��>K��;���v$�Z�����){��-qћ:���|���#�5�-��Ǐ���x��$�4T���.��P��л�����;��c*ç�1��w6�S!�=z\��GU �
���E�>��M�?��t!��� �[�[η#�22�C���)!���|�/��KW3q�̞���z�E%|�ٳ;�9o{�஥E�x�/}��@f�: �b&�!<L<�Y<�Eu'(&�_����Uu�����h%�X1��l��a�FnÎ�T_I�T_�ի8�����:�-�u�%p��q.�ԏ�����ݼ~�-' ��ï�������yE�p���1�3ɘ�������Z%�|d(!����A������@e��ӻSj�)���!]��d��R�I�q�r���N�{�z!G�C|m��V5�L���$,�)��-��q'ԲXX\K��1f�.P6@���3����;�/���؛j��d�x6�x�X�e�sus7��ܦ��pQ�������Q���2�t8�ÈMS�����I�b�*�\ѵ�;�LA�JR*�P�ʧ�q4�2I���Or"`�AF���T��-GAÍ^��%��J$J�Som����(�:Ό�׮�ᒁ��;�\Z;��?d�$�5�V�3�ΦO����#O�)��`[c�b�"jQgm����Yd��n�օ��M�%�S���~
<N�/��n �݂���U�;W��� �}���:�ꁪ���gORC��洪��[�w�y�gς8I+�2*���_�|�˸o�b�P$`4��"�Rtg��m��xp}�����8]/|�9�8[/p�G���9x���P�$c�Wnv.b�H
�ڶh�w`!�KV�B���K�P���xq^@�&uh�����p���hQi��ϧ�7���j���.8�0���a�m%|bs����0���mrq$
��Ǚ���/��
����uPJ��]�S<Y�h"1R	Q�2R� YG.:Μ
�ç���1����=��T9L�5�:q��^��dEGFG�� L`��*����UPZ��<�9���N,yN���8�;;��ut��ڟ!�����Y�y�H���[(��/҄�+��T9`����Pj���!��UU�|�pYY�4�#���̧r��Ō�J�����F8xRB~p���5��H��}�8��� �F�hr����jT����.�Hw�]�D3f̚=��Aۨj γ1���`͚5�l�\�D88�={�l��i�J��rg���y��J����y��<aO]@x�ҷe�.tuC;���(���Y'���x� ��D̘1�E�1(bƹ���IH��:x��ȠQ����'��s���{�S�!	��{��%2tܸq0~�x_f�%-͜�I�&񵌖�f�Y,�9��S޷�g��8�jjꠎ�E,���,��g��{�����@���5v	�����A�T����e���q�J&=u�u�{��ɹV��P=555�g����<����ضZ[����w����#����!�|uv]]-TTT3fs�����^V�ou^ ˗-�'��gz�A8U,(+--�DK������5q�[��~p2$���$|]xm��Ę!�@�IF�Q�^h[v2� ��Q>�}cHEE�X����I�ݼh�KSP�UVt�T� �,���I�����I3���j������d���� 8�)�M&L��mͼ^{G'�fy�T���9�8:��;��S�B�E� 	3���A�㙹apd��[�^2��G�,澗�z�5z��͆H�����X�:��ނ�>'�^be�#	r���YJSEŋ`FSi�O)��\#��jS2��LG��,;ϭ��@IGw�|�(g]i���MxX�{#u�$�<j�}aPV� ��w��T�\�
��s��g�%�f�p���~woo���`a�k}}}N���.�Eh�x�.N����7�1��V������n`٧��C�8x3N_������w�������t2?���Lj�^qI)�f�F,�'���wH./����f�3g~p"�c�LC"�(8�	q��mW޻}Qz;�@�6�.��g���������_2��Z�S�}�h5`;�=�H�ݶ�w���§��0;�������r8�wCww�|��0�gg�~�b��D���Ͱ�h�mڎ�b��B���QR*ъ��[S=��3��K	z��P�i��ͷ��R���X}M�5g��Np�L���X �!Ȟ��'��:���N����y�0u�&��3���8~y"�בb�D;q���p����?����`_ǎ��/���DM��T�E�eu���D�����~�d}U����C72�u"N����d:CLk�_��<��Ox���	��Ĳ(S]4��wVq�/���aX4߀mQv޾����g�l�������8�����Z����c���b��4V�r[[wo��/�����D���;xÍZ]�aW1?�s�K҂!�T��u�1�Q�^z	ݸeK��qܣL�,�>���G.��w�x���!�d2dv__o��q��3l�x����������<rGCCCI>���Ι��F�c��g0,/����W�ylӸ����ݑ�8�ڂ3��I�0��@��t���������θ� ��>��T��N<h2<���41}H��
������2�$�����N�M�!�g�=p���jՒ=
�,8�S��� 8L�l��O����G��w���p��o۶50i�w�uv��v����'�aXKGϰ���8���a��5���O��߹����"0�-Y�Q����d�+P"RxB��r$|�O��|��G�����v��Ȥӑ����?�r{Z���q��ų�F2�t�}w'̚6F��_~R}�g�������!�X�ϐ}��g�>V�3d+��������~��ce?C����!�X�ϐ}��g�>V�3d+��������~��ce?C����!�X�ϐ}��g�>V�3d+��������~��ce?C����!�X�ϐ}����c;����##W�7��ˈ�3�m+nr$v&Q����M.�y4�(o���;Z#b�Gp�����	��eY䝐�<���@��˲6�c���*�{u"+�@i��,�n���.�C�<Ě��ͪq�t F�#�M�Dr���5+<�Ʋ���2����`�������C���e��l,�dw23�Z$�n<�X��w���[wv�h���!H���2<���`�bUTT���-+�Gƌ�ƍ�����)uļP8	F���"F��	zDeu��ǘ�XQ<z}_�� ?�7��M��;�������:�L}��uDIi�DvkG4�����_����F��_�9-�{� �    IEND�B`�PK
     @^�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     @^�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     @^�[�<��s  �s                   cirkitFile.jsonPK 
     @^�[                        �s  jsons/PK 
     @^�[�.��  �               t  jsons/user_defined.jsonPK 
     @^�[                        ?�  images/PK 
     @^�[�R�W�  W�  /             d�  images/e30496d1-6e1c-40fa-a66f-2add70ecdc94.pngPK 
     @^�[$7h�!  �!  /             6 images/a7fde0f7-2836-4f0c-aad0-66dcccec46ff.pngPK 
     @^�[Y�u�= �= /             FX images/1615224e-fb94-4bec-8b91-0567bb6a6470.pngPK 
     @^�[�z��gW  gW  /             K� images/c64d4bdb-8b24-4d1f-9af2-aab9cfab9f47.pngPK 
     @^�[�c��f  �f  /             �� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     @^�[��EM  M  /             -U images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK    
 
   �h   